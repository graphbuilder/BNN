module test_layer1(
clk, 
rstn
);
input clk;
input rstn;

wire P1000;
wire P1010;
wire P1020;
wire P1030;
wire P1040;
wire P1050;
wire P1060;
wire P1070;
wire P1080;
wire P1090;
wire P10A0;
wire P10B0;
wire P10C0;
wire P10D0;
wire P10E0;
wire P10F0;
wire P1100;
wire P1110;
wire P1120;
wire P1130;
wire P1140;
wire P1150;
wire P1160;
wire P1170;
wire P1180;
wire P1190;
wire P11A0;
wire P11B0;
wire P11C0;
wire P11D0;
wire P11E0;
wire P11F0;
wire P1200;
wire P1210;
wire P1220;
wire P1230;
wire P1240;
wire P1250;
wire P1260;
wire P1270;
wire P1280;
wire P1290;
wire P12A0;
wire P12B0;
wire P12C0;
wire P12D0;
wire P12E0;
wire P12F0;
wire P1300;
wire P1310;
wire P1320;
wire P1330;
wire P1340;
wire P1350;
wire P1360;
wire P1370;
wire P1380;
wire P1390;
wire P13A0;
wire P13B0;
wire P13C0;
wire P13D0;
wire P13E0;
wire P13F0;
wire P1400;
wire P1410;
wire P1420;
wire P1430;
wire P1440;
wire P1450;
wire P1460;
wire P1470;
wire P1480;
wire P1490;
wire P14A0;
wire P14B0;
wire P14C0;
wire P14D0;
wire P14E0;
wire P14F0;
wire P1500;
wire P1510;
wire P1520;
wire P1530;
wire P1540;
wire P1550;
wire P1560;
wire P1570;
wire P1580;
wire P1590;
wire P15A0;
wire P15B0;
wire P15C0;
wire P15D0;
wire P15E0;
wire P15F0;
wire P1600;
wire P1610;
wire P1620;
wire P1630;
wire P1640;
wire P1650;
wire P1660;
wire P1670;
wire P1680;
wire P1690;
wire P16A0;
wire P16B0;
wire P16C0;
wire P16D0;
wire P16E0;
wire P16F0;
wire P1700;
wire P1710;
wire P1720;
wire P1730;
wire P1740;
wire P1750;
wire P1760;
wire P1770;
wire P1780;
wire P1790;
wire P17A0;
wire P17B0;
wire P17C0;
wire P17D0;
wire P17E0;
wire P17F0;
wire P1800;
wire P1810;
wire P1820;
wire P1830;
wire P1840;
wire P1850;
wire P1860;
wire P1870;
wire P1880;
wire P1890;
wire P18A0;
wire P18B0;
wire P18C0;
wire P18D0;
wire P18E0;
wire P18F0;
wire P1900;
wire P1910;
wire P1920;
wire P1930;
wire P1940;
wire P1950;
wire P1960;
wire P1970;
wire P1980;
wire P1990;
wire P19A0;
wire P19B0;
wire P19C0;
wire P19D0;
wire P19E0;
wire P19F0;
wire P1A00;
wire P1A10;
wire P1A20;
wire P1A30;
wire P1A40;
wire P1A50;
wire P1A60;
wire P1A70;
wire P1A80;
wire P1A90;
wire P1AA0;
wire P1AB0;
wire P1AC0;
wire P1AD0;
wire P1AE0;
wire P1AF0;
wire P1B00;
wire P1B10;
wire P1B20;
wire P1B30;
wire P1B40;
wire P1B50;
wire P1B60;
wire P1B70;
wire P1B80;
wire P1B90;
wire P1BA0;
wire P1BB0;
wire P1BC0;
wire P1BD0;
wire P1BE0;
wire P1BF0;
wire P1C00;
wire P1C10;
wire P1C20;
wire P1C30;
wire P1C40;
wire P1C50;
wire P1C60;
wire P1C70;
wire P1C80;
wire P1C90;
wire P1CA0;
wire P1CB0;
wire P1CC0;
wire P1CD0;
wire P1CE0;
wire P1CF0;
wire P1D00;
wire P1D10;
wire P1D20;
wire P1D30;
wire P1D40;
wire P1D50;
wire P1D60;
wire P1D70;
wire P1D80;
wire P1D90;
wire P1DA0;
wire P1DB0;
wire P1DC0;
wire P1DD0;
wire P1DE0;
wire P1DF0;
wire P1E00;
wire P1E10;
wire P1E20;
wire P1E30;
wire P1E40;
wire P1E50;
wire P1E60;
wire P1E70;
wire P1E80;
wire P1E90;
wire P1EA0;
wire P1EB0;
wire P1EC0;
wire P1ED0;
wire P1EE0;
wire P1EF0;
wire P1F00;
wire P1F10;
wire P1F20;
wire P1F30;
wire P1F40;
wire P1F50;
wire P1F60;
wire P1F70;
wire P1F80;
wire P1F90;
wire P1FA0;
wire P1FB0;
wire P1FC0;
wire P1FD0;
wire P1FE0;
wire P1FF0;
wire P1001;
wire P1011;
wire P1021;
wire P1031;
wire P1041;
wire P1051;
wire P1061;
wire P1071;
wire P1081;
wire P1091;
wire P10A1;
wire P10B1;
wire P10C1;
wire P10D1;
wire P10E1;
wire P10F1;
wire P1101;
wire P1111;
wire P1121;
wire P1131;
wire P1141;
wire P1151;
wire P1161;
wire P1171;
wire P1181;
wire P1191;
wire P11A1;
wire P11B1;
wire P11C1;
wire P11D1;
wire P11E1;
wire P11F1;
wire P1201;
wire P1211;
wire P1221;
wire P1231;
wire P1241;
wire P1251;
wire P1261;
wire P1271;
wire P1281;
wire P1291;
wire P12A1;
wire P12B1;
wire P12C1;
wire P12D1;
wire P12E1;
wire P12F1;
wire P1301;
wire P1311;
wire P1321;
wire P1331;
wire P1341;
wire P1351;
wire P1361;
wire P1371;
wire P1381;
wire P1391;
wire P13A1;
wire P13B1;
wire P13C1;
wire P13D1;
wire P13E1;
wire P13F1;
wire P1401;
wire P1411;
wire P1421;
wire P1431;
wire P1441;
wire P1451;
wire P1461;
wire P1471;
wire P1481;
wire P1491;
wire P14A1;
wire P14B1;
wire P14C1;
wire P14D1;
wire P14E1;
wire P14F1;
wire P1501;
wire P1511;
wire P1521;
wire P1531;
wire P1541;
wire P1551;
wire P1561;
wire P1571;
wire P1581;
wire P1591;
wire P15A1;
wire P15B1;
wire P15C1;
wire P15D1;
wire P15E1;
wire P15F1;
wire P1601;
wire P1611;
wire P1621;
wire P1631;
wire P1641;
wire P1651;
wire P1661;
wire P1671;
wire P1681;
wire P1691;
wire P16A1;
wire P16B1;
wire P16C1;
wire P16D1;
wire P16E1;
wire P16F1;
wire P1701;
wire P1711;
wire P1721;
wire P1731;
wire P1741;
wire P1751;
wire P1761;
wire P1771;
wire P1781;
wire P1791;
wire P17A1;
wire P17B1;
wire P17C1;
wire P17D1;
wire P17E1;
wire P17F1;
wire P1801;
wire P1811;
wire P1821;
wire P1831;
wire P1841;
wire P1851;
wire P1861;
wire P1871;
wire P1881;
wire P1891;
wire P18A1;
wire P18B1;
wire P18C1;
wire P18D1;
wire P18E1;
wire P18F1;
wire P1901;
wire P1911;
wire P1921;
wire P1931;
wire P1941;
wire P1951;
wire P1961;
wire P1971;
wire P1981;
wire P1991;
wire P19A1;
wire P19B1;
wire P19C1;
wire P19D1;
wire P19E1;
wire P19F1;
wire P1A01;
wire P1A11;
wire P1A21;
wire P1A31;
wire P1A41;
wire P1A51;
wire P1A61;
wire P1A71;
wire P1A81;
wire P1A91;
wire P1AA1;
wire P1AB1;
wire P1AC1;
wire P1AD1;
wire P1AE1;
wire P1AF1;
wire P1B01;
wire P1B11;
wire P1B21;
wire P1B31;
wire P1B41;
wire P1B51;
wire P1B61;
wire P1B71;
wire P1B81;
wire P1B91;
wire P1BA1;
wire P1BB1;
wire P1BC1;
wire P1BD1;
wire P1BE1;
wire P1BF1;
wire P1C01;
wire P1C11;
wire P1C21;
wire P1C31;
wire P1C41;
wire P1C51;
wire P1C61;
wire P1C71;
wire P1C81;
wire P1C91;
wire P1CA1;
wire P1CB1;
wire P1CC1;
wire P1CD1;
wire P1CE1;
wire P1CF1;
wire P1D01;
wire P1D11;
wire P1D21;
wire P1D31;
wire P1D41;
wire P1D51;
wire P1D61;
wire P1D71;
wire P1D81;
wire P1D91;
wire P1DA1;
wire P1DB1;
wire P1DC1;
wire P1DD1;
wire P1DE1;
wire P1DF1;
wire P1E01;
wire P1E11;
wire P1E21;
wire P1E31;
wire P1E41;
wire P1E51;
wire P1E61;
wire P1E71;
wire P1E81;
wire P1E91;
wire P1EA1;
wire P1EB1;
wire P1EC1;
wire P1ED1;
wire P1EE1;
wire P1EF1;
wire P1F01;
wire P1F11;
wire P1F21;
wire P1F31;
wire P1F41;
wire P1F51;
wire P1F61;
wire P1F71;
wire P1F81;
wire P1F91;
wire P1FA1;
wire P1FB1;
wire P1FC1;
wire P1FD1;
wire P1FE1;
wire P1FF1;
wire P1002;
wire P1012;
wire P1022;
wire P1032;
wire P1042;
wire P1052;
wire P1062;
wire P1072;
wire P1082;
wire P1092;
wire P10A2;
wire P10B2;
wire P10C2;
wire P10D2;
wire P10E2;
wire P10F2;
wire P1102;
wire P1112;
wire P1122;
wire P1132;
wire P1142;
wire P1152;
wire P1162;
wire P1172;
wire P1182;
wire P1192;
wire P11A2;
wire P11B2;
wire P11C2;
wire P11D2;
wire P11E2;
wire P11F2;
wire P1202;
wire P1212;
wire P1222;
wire P1232;
wire P1242;
wire P1252;
wire P1262;
wire P1272;
wire P1282;
wire P1292;
wire P12A2;
wire P12B2;
wire P12C2;
wire P12D2;
wire P12E2;
wire P12F2;
wire P1302;
wire P1312;
wire P1322;
wire P1332;
wire P1342;
wire P1352;
wire P1362;
wire P1372;
wire P1382;
wire P1392;
wire P13A2;
wire P13B2;
wire P13C2;
wire P13D2;
wire P13E2;
wire P13F2;
wire P1402;
wire P1412;
wire P1422;
wire P1432;
wire P1442;
wire P1452;
wire P1462;
wire P1472;
wire P1482;
wire P1492;
wire P14A2;
wire P14B2;
wire P14C2;
wire P14D2;
wire P14E2;
wire P14F2;
wire P1502;
wire P1512;
wire P1522;
wire P1532;
wire P1542;
wire P1552;
wire P1562;
wire P1572;
wire P1582;
wire P1592;
wire P15A2;
wire P15B2;
wire P15C2;
wire P15D2;
wire P15E2;
wire P15F2;
wire P1602;
wire P1612;
wire P1622;
wire P1632;
wire P1642;
wire P1652;
wire P1662;
wire P1672;
wire P1682;
wire P1692;
wire P16A2;
wire P16B2;
wire P16C2;
wire P16D2;
wire P16E2;
wire P16F2;
wire P1702;
wire P1712;
wire P1722;
wire P1732;
wire P1742;
wire P1752;
wire P1762;
wire P1772;
wire P1782;
wire P1792;
wire P17A2;
wire P17B2;
wire P17C2;
wire P17D2;
wire P17E2;
wire P17F2;
wire P1802;
wire P1812;
wire P1822;
wire P1832;
wire P1842;
wire P1852;
wire P1862;
wire P1872;
wire P1882;
wire P1892;
wire P18A2;
wire P18B2;
wire P18C2;
wire P18D2;
wire P18E2;
wire P18F2;
wire P1902;
wire P1912;
wire P1922;
wire P1932;
wire P1942;
wire P1952;
wire P1962;
wire P1972;
wire P1982;
wire P1992;
wire P19A2;
wire P19B2;
wire P19C2;
wire P19D2;
wire P19E2;
wire P19F2;
wire P1A02;
wire P1A12;
wire P1A22;
wire P1A32;
wire P1A42;
wire P1A52;
wire P1A62;
wire P1A72;
wire P1A82;
wire P1A92;
wire P1AA2;
wire P1AB2;
wire P1AC2;
wire P1AD2;
wire P1AE2;
wire P1AF2;
wire P1B02;
wire P1B12;
wire P1B22;
wire P1B32;
wire P1B42;
wire P1B52;
wire P1B62;
wire P1B72;
wire P1B82;
wire P1B92;
wire P1BA2;
wire P1BB2;
wire P1BC2;
wire P1BD2;
wire P1BE2;
wire P1BF2;
wire P1C02;
wire P1C12;
wire P1C22;
wire P1C32;
wire P1C42;
wire P1C52;
wire P1C62;
wire P1C72;
wire P1C82;
wire P1C92;
wire P1CA2;
wire P1CB2;
wire P1CC2;
wire P1CD2;
wire P1CE2;
wire P1CF2;
wire P1D02;
wire P1D12;
wire P1D22;
wire P1D32;
wire P1D42;
wire P1D52;
wire P1D62;
wire P1D72;
wire P1D82;
wire P1D92;
wire P1DA2;
wire P1DB2;
wire P1DC2;
wire P1DD2;
wire P1DE2;
wire P1DF2;
wire P1E02;
wire P1E12;
wire P1E22;
wire P1E32;
wire P1E42;
wire P1E52;
wire P1E62;
wire P1E72;
wire P1E82;
wire P1E92;
wire P1EA2;
wire P1EB2;
wire P1EC2;
wire P1ED2;
wire P1EE2;
wire P1EF2;
wire P1F02;
wire P1F12;
wire P1F22;
wire P1F32;
wire P1F42;
wire P1F52;
wire P1F62;
wire P1F72;
wire P1F82;
wire P1F92;
wire P1FA2;
wire P1FB2;
wire P1FC2;
wire P1FD2;
wire P1FE2;
wire P1FF2;
wire P1003;
wire P1013;
wire P1023;
wire P1033;
wire P1043;
wire P1053;
wire P1063;
wire P1073;
wire P1083;
wire P1093;
wire P10A3;
wire P10B3;
wire P10C3;
wire P10D3;
wire P10E3;
wire P10F3;
wire P1103;
wire P1113;
wire P1123;
wire P1133;
wire P1143;
wire P1153;
wire P1163;
wire P1173;
wire P1183;
wire P1193;
wire P11A3;
wire P11B3;
wire P11C3;
wire P11D3;
wire P11E3;
wire P11F3;
wire P1203;
wire P1213;
wire P1223;
wire P1233;
wire P1243;
wire P1253;
wire P1263;
wire P1273;
wire P1283;
wire P1293;
wire P12A3;
wire P12B3;
wire P12C3;
wire P12D3;
wire P12E3;
wire P12F3;
wire P1303;
wire P1313;
wire P1323;
wire P1333;
wire P1343;
wire P1353;
wire P1363;
wire P1373;
wire P1383;
wire P1393;
wire P13A3;
wire P13B3;
wire P13C3;
wire P13D3;
wire P13E3;
wire P13F3;
wire P1403;
wire P1413;
wire P1423;
wire P1433;
wire P1443;
wire P1453;
wire P1463;
wire P1473;
wire P1483;
wire P1493;
wire P14A3;
wire P14B3;
wire P14C3;
wire P14D3;
wire P14E3;
wire P14F3;
wire P1503;
wire P1513;
wire P1523;
wire P1533;
wire P1543;
wire P1553;
wire P1563;
wire P1573;
wire P1583;
wire P1593;
wire P15A3;
wire P15B3;
wire P15C3;
wire P15D3;
wire P15E3;
wire P15F3;
wire P1603;
wire P1613;
wire P1623;
wire P1633;
wire P1643;
wire P1653;
wire P1663;
wire P1673;
wire P1683;
wire P1693;
wire P16A3;
wire P16B3;
wire P16C3;
wire P16D3;
wire P16E3;
wire P16F3;
wire P1703;
wire P1713;
wire P1723;
wire P1733;
wire P1743;
wire P1753;
wire P1763;
wire P1773;
wire P1783;
wire P1793;
wire P17A3;
wire P17B3;
wire P17C3;
wire P17D3;
wire P17E3;
wire P17F3;
wire P1803;
wire P1813;
wire P1823;
wire P1833;
wire P1843;
wire P1853;
wire P1863;
wire P1873;
wire P1883;
wire P1893;
wire P18A3;
wire P18B3;
wire P18C3;
wire P18D3;
wire P18E3;
wire P18F3;
wire P1903;
wire P1913;
wire P1923;
wire P1933;
wire P1943;
wire P1953;
wire P1963;
wire P1973;
wire P1983;
wire P1993;
wire P19A3;
wire P19B3;
wire P19C3;
wire P19D3;
wire P19E3;
wire P19F3;
wire P1A03;
wire P1A13;
wire P1A23;
wire P1A33;
wire P1A43;
wire P1A53;
wire P1A63;
wire P1A73;
wire P1A83;
wire P1A93;
wire P1AA3;
wire P1AB3;
wire P1AC3;
wire P1AD3;
wire P1AE3;
wire P1AF3;
wire P1B03;
wire P1B13;
wire P1B23;
wire P1B33;
wire P1B43;
wire P1B53;
wire P1B63;
wire P1B73;
wire P1B83;
wire P1B93;
wire P1BA3;
wire P1BB3;
wire P1BC3;
wire P1BD3;
wire P1BE3;
wire P1BF3;
wire P1C03;
wire P1C13;
wire P1C23;
wire P1C33;
wire P1C43;
wire P1C53;
wire P1C63;
wire P1C73;
wire P1C83;
wire P1C93;
wire P1CA3;
wire P1CB3;
wire P1CC3;
wire P1CD3;
wire P1CE3;
wire P1CF3;
wire P1D03;
wire P1D13;
wire P1D23;
wire P1D33;
wire P1D43;
wire P1D53;
wire P1D63;
wire P1D73;
wire P1D83;
wire P1D93;
wire P1DA3;
wire P1DB3;
wire P1DC3;
wire P1DD3;
wire P1DE3;
wire P1DF3;
wire P1E03;
wire P1E13;
wire P1E23;
wire P1E33;
wire P1E43;
wire P1E53;
wire P1E63;
wire P1E73;
wire P1E83;
wire P1E93;
wire P1EA3;
wire P1EB3;
wire P1EC3;
wire P1ED3;
wire P1EE3;
wire P1EF3;
wire P1F03;
wire P1F13;
wire P1F23;
wire P1F33;
wire P1F43;
wire P1F53;
wire P1F63;
wire P1F73;
wire P1F83;
wire P1F93;
wire P1FA3;
wire P1FB3;
wire P1FC3;
wire P1FD3;
wire P1FE3;
wire P1FF3;
wire P2000;
wire P2010;
wire P2020;
wire P2030;
wire P2040;
wire P2050;
wire P2060;
wire P2100;
wire P2110;
wire P2120;
wire P2130;
wire P2140;
wire P2150;
wire P2160;
wire P2200;
wire P2210;
wire P2220;
wire P2230;
wire P2240;
wire P2250;
wire P2260;
wire P2300;
wire P2310;
wire P2320;
wire P2330;
wire P2340;
wire P2350;
wire P2360;
wire P2400;
wire P2410;
wire P2420;
wire P2430;
wire P2440;
wire P2450;
wire P2460;
wire P2500;
wire P2510;
wire P2520;
wire P2530;
wire P2540;
wire P2550;
wire P2560;
wire P2600;
wire P2610;
wire P2620;
wire P2630;
wire P2640;
wire P2650;
wire P2660;
wire P2001;
wire P2011;
wire P2021;
wire P2031;
wire P2041;
wire P2051;
wire P2061;
wire P2101;
wire P2111;
wire P2121;
wire P2131;
wire P2141;
wire P2151;
wire P2161;
wire P2201;
wire P2211;
wire P2221;
wire P2231;
wire P2241;
wire P2251;
wire P2261;
wire P2301;
wire P2311;
wire P2321;
wire P2331;
wire P2341;
wire P2351;
wire P2361;
wire P2401;
wire P2411;
wire P2421;
wire P2431;
wire P2441;
wire P2451;
wire P2461;
wire P2501;
wire P2511;
wire P2521;
wire P2531;
wire P2541;
wire P2551;
wire P2561;
wire P2601;
wire P2611;
wire P2621;
wire P2631;
wire P2641;
wire P2651;
wire P2661;
wire P2002;
wire P2012;
wire P2022;
wire P2032;
wire P2042;
wire P2052;
wire P2062;
wire P2102;
wire P2112;
wire P2122;
wire P2132;
wire P2142;
wire P2152;
wire P2162;
wire P2202;
wire P2212;
wire P2222;
wire P2232;
wire P2242;
wire P2252;
wire P2262;
wire P2302;
wire P2312;
wire P2322;
wire P2332;
wire P2342;
wire P2352;
wire P2362;
wire P2402;
wire P2412;
wire P2422;
wire P2432;
wire P2442;
wire P2452;
wire P2462;
wire P2502;
wire P2512;
wire P2522;
wire P2532;
wire P2542;
wire P2552;
wire P2562;
wire P2602;
wire P2612;
wire P2622;
wire P2632;
wire P2642;
wire P2652;
wire P2662;
wire P2003;
wire P2013;
wire P2023;
wire P2033;
wire P2043;
wire P2053;
wire P2063;
wire P2103;
wire P2113;
wire P2123;
wire P2133;
wire P2143;
wire P2153;
wire P2163;
wire P2203;
wire P2213;
wire P2223;
wire P2233;
wire P2243;
wire P2253;
wire P2263;
wire P2303;
wire P2313;
wire P2323;
wire P2333;
wire P2343;
wire P2353;
wire P2363;
wire P2403;
wire P2413;
wire P2423;
wire P2433;
wire P2443;
wire P2453;
wire P2463;
wire P2503;
wire P2513;
wire P2523;
wire P2533;
wire P2543;
wire P2553;
wire P2563;
wire P2603;
wire P2613;
wire P2623;
wire P2633;
wire P2643;
wire P2653;
wire P2663;
wire P2004;
wire P2014;
wire P2024;
wire P2034;
wire P2044;
wire P2054;
wire P2064;
wire P2104;
wire P2114;
wire P2124;
wire P2134;
wire P2144;
wire P2154;
wire P2164;
wire P2204;
wire P2214;
wire P2224;
wire P2234;
wire P2244;
wire P2254;
wire P2264;
wire P2304;
wire P2314;
wire P2324;
wire P2334;
wire P2344;
wire P2354;
wire P2364;
wire P2404;
wire P2414;
wire P2424;
wire P2434;
wire P2444;
wire P2454;
wire P2464;
wire P2504;
wire P2514;
wire P2524;
wire P2534;
wire P2544;
wire P2554;
wire P2564;
wire P2604;
wire P2614;
wire P2624;
wire P2634;
wire P2644;
wire P2654;
wire P2664;
wire P2005;
wire P2015;
wire P2025;
wire P2035;
wire P2045;
wire P2055;
wire P2065;
wire P2105;
wire P2115;
wire P2125;
wire P2135;
wire P2145;
wire P2155;
wire P2165;
wire P2205;
wire P2215;
wire P2225;
wire P2235;
wire P2245;
wire P2255;
wire P2265;
wire P2305;
wire P2315;
wire P2325;
wire P2335;
wire P2345;
wire P2355;
wire P2365;
wire P2405;
wire P2415;
wire P2425;
wire P2435;
wire P2445;
wire P2455;
wire P2465;
wire P2505;
wire P2515;
wire P2525;
wire P2535;
wire P2545;
wire P2555;
wire P2565;
wire P2605;
wire P2615;
wire P2625;
wire P2635;
wire P2645;
wire P2655;
wire P2665;
wire P2006;
wire P2016;
wire P2026;
wire P2036;
wire P2046;
wire P2056;
wire P2066;
wire P2106;
wire P2116;
wire P2126;
wire P2136;
wire P2146;
wire P2156;
wire P2166;
wire P2206;
wire P2216;
wire P2226;
wire P2236;
wire P2246;
wire P2256;
wire P2266;
wire P2306;
wire P2316;
wire P2326;
wire P2336;
wire P2346;
wire P2356;
wire P2366;
wire P2406;
wire P2416;
wire P2426;
wire P2436;
wire P2446;
wire P2456;
wire P2466;
wire P2506;
wire P2516;
wire P2526;
wire P2536;
wire P2546;
wire P2556;
wire P2566;
wire P2606;
wire P2616;
wire P2626;
wire P2636;
wire P2646;
wire P2656;
wire P2666;
wire P2007;
wire P2017;
wire P2027;
wire P2037;
wire P2047;
wire P2057;
wire P2067;
wire P2107;
wire P2117;
wire P2127;
wire P2137;
wire P2147;
wire P2157;
wire P2167;
wire P2207;
wire P2217;
wire P2227;
wire P2237;
wire P2247;
wire P2257;
wire P2267;
wire P2307;
wire P2317;
wire P2327;
wire P2337;
wire P2347;
wire P2357;
wire P2367;
wire P2407;
wire P2417;
wire P2427;
wire P2437;
wire P2447;
wire P2457;
wire P2467;
wire P2507;
wire P2517;
wire P2527;
wire P2537;
wire P2547;
wire P2557;
wire P2567;
wire P2607;
wire P2617;
wire P2627;
wire P2637;
wire P2647;
wire P2657;
wire P2667;
wire W10000,W10010,W10020,W10100,W10110,W10120,W10200,W10210,W10220;
wire W10001,W10011,W10021,W10101,W10111,W10121,W10201,W10211,W10221;
wire W10002,W10012,W10022,W10102,W10112,W10122,W10202,W10212,W10222;
wire W10003,W10013,W10023,W10103,W10113,W10123,W10203,W10213,W10223;
wire W11000,W11010,W11020,W11100,W11110,W11120,W11200,W11210,W11220;
wire W11001,W11011,W11021,W11101,W11111,W11121,W11201,W11211,W11221;
wire W11002,W11012,W11022,W11102,W11112,W11122,W11202,W11212,W11222;
wire W11003,W11013,W11023,W11103,W11113,W11123,W11203,W11213,W11223;
wire W12000,W12010,W12020,W12100,W12110,W12120,W12200,W12210,W12220;
wire W12001,W12011,W12021,W12101,W12111,W12121,W12201,W12211,W12221;
wire W12002,W12012,W12022,W12102,W12112,W12122,W12202,W12212,W12222;
wire W12003,W12013,W12023,W12103,W12113,W12123,W12203,W12213,W12223;
wire W13000,W13010,W13020,W13100,W13110,W13120,W13200,W13210,W13220;
wire W13001,W13011,W13021,W13101,W13111,W13121,W13201,W13211,W13221;
wire W13002,W13012,W13022,W13102,W13112,W13122,W13202,W13212,W13222;
wire W13003,W13013,W13023,W13103,W13113,W13123,W13203,W13213,W13223;
wire W14000,W14010,W14020,W14100,W14110,W14120,W14200,W14210,W14220;
wire W14001,W14011,W14021,W14101,W14111,W14121,W14201,W14211,W14221;
wire W14002,W14012,W14022,W14102,W14112,W14122,W14202,W14212,W14222;
wire W14003,W14013,W14023,W14103,W14113,W14123,W14203,W14213,W14223;
wire W15000,W15010,W15020,W15100,W15110,W15120,W15200,W15210,W15220;
wire W15001,W15011,W15021,W15101,W15111,W15121,W15201,W15211,W15221;
wire W15002,W15012,W15022,W15102,W15112,W15122,W15202,W15212,W15222;
wire W15003,W15013,W15023,W15103,W15113,W15123,W15203,W15213,W15223;
wire W16000,W16010,W16020,W16100,W16110,W16120,W16200,W16210,W16220;
wire W16001,W16011,W16021,W16101,W16111,W16121,W16201,W16211,W16221;
wire W16002,W16012,W16022,W16102,W16112,W16122,W16202,W16212,W16222;
wire W16003,W16013,W16023,W16103,W16113,W16123,W16203,W16213,W16223;
wire W17000,W17010,W17020,W17100,W17110,W17120,W17200,W17210,W17220;
wire W17001,W17011,W17021,W17101,W17111,W17121,W17201,W17211,W17221;
wire W17002,W17012,W17022,W17102,W17112,W17122,W17202,W17212,W17222;
wire W17003,W17013,W17023,W17103,W17113,W17123,W17203,W17213,W17223;
wire signed [4:0] c10000,c11000,c12000,c13000;
wire signed [4:0] c10010,c11010,c12010,c13010;
wire signed [4:0] c10020,c11020,c12020,c13020;
wire signed [4:0] c10030,c11030,c12030,c13030;
wire signed [4:0] c10040,c11040,c12040,c13040;
wire signed [4:0] c10050,c11050,c12050,c13050;
wire signed [4:0] c10060,c11060,c12060,c13060;
wire signed [4:0] c10070,c11070,c12070,c13070;
wire signed [4:0] c10080,c11080,c12080,c13080;
wire signed [4:0] c10090,c11090,c12090,c13090;
wire signed [4:0] c100A0,c110A0,c120A0,c130A0;
wire signed [4:0] c100B0,c110B0,c120B0,c130B0;
wire signed [4:0] c100C0,c110C0,c120C0,c130C0;
wire signed [4:0] c100D0,c110D0,c120D0,c130D0;
wire signed [4:0] c10100,c11100,c12100,c13100;
wire signed [4:0] c10110,c11110,c12110,c13110;
wire signed [4:0] c10120,c11120,c12120,c13120;
wire signed [4:0] c10130,c11130,c12130,c13130;
wire signed [4:0] c10140,c11140,c12140,c13140;
wire signed [4:0] c10150,c11150,c12150,c13150;
wire signed [4:0] c10160,c11160,c12160,c13160;
wire signed [4:0] c10170,c11170,c12170,c13170;
wire signed [4:0] c10180,c11180,c12180,c13180;
wire signed [4:0] c10190,c11190,c12190,c13190;
wire signed [4:0] c101A0,c111A0,c121A0,c131A0;
wire signed [4:0] c101B0,c111B0,c121B0,c131B0;
wire signed [4:0] c101C0,c111C0,c121C0,c131C0;
wire signed [4:0] c101D0,c111D0,c121D0,c131D0;
wire signed [4:0] c10200,c11200,c12200,c13200;
wire signed [4:0] c10210,c11210,c12210,c13210;
wire signed [4:0] c10220,c11220,c12220,c13220;
wire signed [4:0] c10230,c11230,c12230,c13230;
wire signed [4:0] c10240,c11240,c12240,c13240;
wire signed [4:0] c10250,c11250,c12250,c13250;
wire signed [4:0] c10260,c11260,c12260,c13260;
wire signed [4:0] c10270,c11270,c12270,c13270;
wire signed [4:0] c10280,c11280,c12280,c13280;
wire signed [4:0] c10290,c11290,c12290,c13290;
wire signed [4:0] c102A0,c112A0,c122A0,c132A0;
wire signed [4:0] c102B0,c112B0,c122B0,c132B0;
wire signed [4:0] c102C0,c112C0,c122C0,c132C0;
wire signed [4:0] c102D0,c112D0,c122D0,c132D0;
wire signed [4:0] c10300,c11300,c12300,c13300;
wire signed [4:0] c10310,c11310,c12310,c13310;
wire signed [4:0] c10320,c11320,c12320,c13320;
wire signed [4:0] c10330,c11330,c12330,c13330;
wire signed [4:0] c10340,c11340,c12340,c13340;
wire signed [4:0] c10350,c11350,c12350,c13350;
wire signed [4:0] c10360,c11360,c12360,c13360;
wire signed [4:0] c10370,c11370,c12370,c13370;
wire signed [4:0] c10380,c11380,c12380,c13380;
wire signed [4:0] c10390,c11390,c12390,c13390;
wire signed [4:0] c103A0,c113A0,c123A0,c133A0;
wire signed [4:0] c103B0,c113B0,c123B0,c133B0;
wire signed [4:0] c103C0,c113C0,c123C0,c133C0;
wire signed [4:0] c103D0,c113D0,c123D0,c133D0;
wire signed [4:0] c10400,c11400,c12400,c13400;
wire signed [4:0] c10410,c11410,c12410,c13410;
wire signed [4:0] c10420,c11420,c12420,c13420;
wire signed [4:0] c10430,c11430,c12430,c13430;
wire signed [4:0] c10440,c11440,c12440,c13440;
wire signed [4:0] c10450,c11450,c12450,c13450;
wire signed [4:0] c10460,c11460,c12460,c13460;
wire signed [4:0] c10470,c11470,c12470,c13470;
wire signed [4:0] c10480,c11480,c12480,c13480;
wire signed [4:0] c10490,c11490,c12490,c13490;
wire signed [4:0] c104A0,c114A0,c124A0,c134A0;
wire signed [4:0] c104B0,c114B0,c124B0,c134B0;
wire signed [4:0] c104C0,c114C0,c124C0,c134C0;
wire signed [4:0] c104D0,c114D0,c124D0,c134D0;
wire signed [4:0] c10500,c11500,c12500,c13500;
wire signed [4:0] c10510,c11510,c12510,c13510;
wire signed [4:0] c10520,c11520,c12520,c13520;
wire signed [4:0] c10530,c11530,c12530,c13530;
wire signed [4:0] c10540,c11540,c12540,c13540;
wire signed [4:0] c10550,c11550,c12550,c13550;
wire signed [4:0] c10560,c11560,c12560,c13560;
wire signed [4:0] c10570,c11570,c12570,c13570;
wire signed [4:0] c10580,c11580,c12580,c13580;
wire signed [4:0] c10590,c11590,c12590,c13590;
wire signed [4:0] c105A0,c115A0,c125A0,c135A0;
wire signed [4:0] c105B0,c115B0,c125B0,c135B0;
wire signed [4:0] c105C0,c115C0,c125C0,c135C0;
wire signed [4:0] c105D0,c115D0,c125D0,c135D0;
wire signed [4:0] c10600,c11600,c12600,c13600;
wire signed [4:0] c10610,c11610,c12610,c13610;
wire signed [4:0] c10620,c11620,c12620,c13620;
wire signed [4:0] c10630,c11630,c12630,c13630;
wire signed [4:0] c10640,c11640,c12640,c13640;
wire signed [4:0] c10650,c11650,c12650,c13650;
wire signed [4:0] c10660,c11660,c12660,c13660;
wire signed [4:0] c10670,c11670,c12670,c13670;
wire signed [4:0] c10680,c11680,c12680,c13680;
wire signed [4:0] c10690,c11690,c12690,c13690;
wire signed [4:0] c106A0,c116A0,c126A0,c136A0;
wire signed [4:0] c106B0,c116B0,c126B0,c136B0;
wire signed [4:0] c106C0,c116C0,c126C0,c136C0;
wire signed [4:0] c106D0,c116D0,c126D0,c136D0;
wire signed [4:0] c10700,c11700,c12700,c13700;
wire signed [4:0] c10710,c11710,c12710,c13710;
wire signed [4:0] c10720,c11720,c12720,c13720;
wire signed [4:0] c10730,c11730,c12730,c13730;
wire signed [4:0] c10740,c11740,c12740,c13740;
wire signed [4:0] c10750,c11750,c12750,c13750;
wire signed [4:0] c10760,c11760,c12760,c13760;
wire signed [4:0] c10770,c11770,c12770,c13770;
wire signed [4:0] c10780,c11780,c12780,c13780;
wire signed [4:0] c10790,c11790,c12790,c13790;
wire signed [4:0] c107A0,c117A0,c127A0,c137A0;
wire signed [4:0] c107B0,c117B0,c127B0,c137B0;
wire signed [4:0] c107C0,c117C0,c127C0,c137C0;
wire signed [4:0] c107D0,c117D0,c127D0,c137D0;
wire signed [4:0] c10800,c11800,c12800,c13800;
wire signed [4:0] c10810,c11810,c12810,c13810;
wire signed [4:0] c10820,c11820,c12820,c13820;
wire signed [4:0] c10830,c11830,c12830,c13830;
wire signed [4:0] c10840,c11840,c12840,c13840;
wire signed [4:0] c10850,c11850,c12850,c13850;
wire signed [4:0] c10860,c11860,c12860,c13860;
wire signed [4:0] c10870,c11870,c12870,c13870;
wire signed [4:0] c10880,c11880,c12880,c13880;
wire signed [4:0] c10890,c11890,c12890,c13890;
wire signed [4:0] c108A0,c118A0,c128A0,c138A0;
wire signed [4:0] c108B0,c118B0,c128B0,c138B0;
wire signed [4:0] c108C0,c118C0,c128C0,c138C0;
wire signed [4:0] c108D0,c118D0,c128D0,c138D0;
wire signed [4:0] c10900,c11900,c12900,c13900;
wire signed [4:0] c10910,c11910,c12910,c13910;
wire signed [4:0] c10920,c11920,c12920,c13920;
wire signed [4:0] c10930,c11930,c12930,c13930;
wire signed [4:0] c10940,c11940,c12940,c13940;
wire signed [4:0] c10950,c11950,c12950,c13950;
wire signed [4:0] c10960,c11960,c12960,c13960;
wire signed [4:0] c10970,c11970,c12970,c13970;
wire signed [4:0] c10980,c11980,c12980,c13980;
wire signed [4:0] c10990,c11990,c12990,c13990;
wire signed [4:0] c109A0,c119A0,c129A0,c139A0;
wire signed [4:0] c109B0,c119B0,c129B0,c139B0;
wire signed [4:0] c109C0,c119C0,c129C0,c139C0;
wire signed [4:0] c109D0,c119D0,c129D0,c139D0;
wire signed [4:0] c10A00,c11A00,c12A00,c13A00;
wire signed [4:0] c10A10,c11A10,c12A10,c13A10;
wire signed [4:0] c10A20,c11A20,c12A20,c13A20;
wire signed [4:0] c10A30,c11A30,c12A30,c13A30;
wire signed [4:0] c10A40,c11A40,c12A40,c13A40;
wire signed [4:0] c10A50,c11A50,c12A50,c13A50;
wire signed [4:0] c10A60,c11A60,c12A60,c13A60;
wire signed [4:0] c10A70,c11A70,c12A70,c13A70;
wire signed [4:0] c10A80,c11A80,c12A80,c13A80;
wire signed [4:0] c10A90,c11A90,c12A90,c13A90;
wire signed [4:0] c10AA0,c11AA0,c12AA0,c13AA0;
wire signed [4:0] c10AB0,c11AB0,c12AB0,c13AB0;
wire signed [4:0] c10AC0,c11AC0,c12AC0,c13AC0;
wire signed [4:0] c10AD0,c11AD0,c12AD0,c13AD0;
wire signed [4:0] c10B00,c11B00,c12B00,c13B00;
wire signed [4:0] c10B10,c11B10,c12B10,c13B10;
wire signed [4:0] c10B20,c11B20,c12B20,c13B20;
wire signed [4:0] c10B30,c11B30,c12B30,c13B30;
wire signed [4:0] c10B40,c11B40,c12B40,c13B40;
wire signed [4:0] c10B50,c11B50,c12B50,c13B50;
wire signed [4:0] c10B60,c11B60,c12B60,c13B60;
wire signed [4:0] c10B70,c11B70,c12B70,c13B70;
wire signed [4:0] c10B80,c11B80,c12B80,c13B80;
wire signed [4:0] c10B90,c11B90,c12B90,c13B90;
wire signed [4:0] c10BA0,c11BA0,c12BA0,c13BA0;
wire signed [4:0] c10BB0,c11BB0,c12BB0,c13BB0;
wire signed [4:0] c10BC0,c11BC0,c12BC0,c13BC0;
wire signed [4:0] c10BD0,c11BD0,c12BD0,c13BD0;
wire signed [4:0] c10C00,c11C00,c12C00,c13C00;
wire signed [4:0] c10C10,c11C10,c12C10,c13C10;
wire signed [4:0] c10C20,c11C20,c12C20,c13C20;
wire signed [4:0] c10C30,c11C30,c12C30,c13C30;
wire signed [4:0] c10C40,c11C40,c12C40,c13C40;
wire signed [4:0] c10C50,c11C50,c12C50,c13C50;
wire signed [4:0] c10C60,c11C60,c12C60,c13C60;
wire signed [4:0] c10C70,c11C70,c12C70,c13C70;
wire signed [4:0] c10C80,c11C80,c12C80,c13C80;
wire signed [4:0] c10C90,c11C90,c12C90,c13C90;
wire signed [4:0] c10CA0,c11CA0,c12CA0,c13CA0;
wire signed [4:0] c10CB0,c11CB0,c12CB0,c13CB0;
wire signed [4:0] c10CC0,c11CC0,c12CC0,c13CC0;
wire signed [4:0] c10CD0,c11CD0,c12CD0,c13CD0;
wire signed [4:0] c10D00,c11D00,c12D00,c13D00;
wire signed [4:0] c10D10,c11D10,c12D10,c13D10;
wire signed [4:0] c10D20,c11D20,c12D20,c13D20;
wire signed [4:0] c10D30,c11D30,c12D30,c13D30;
wire signed [4:0] c10D40,c11D40,c12D40,c13D40;
wire signed [4:0] c10D50,c11D50,c12D50,c13D50;
wire signed [4:0] c10D60,c11D60,c12D60,c13D60;
wire signed [4:0] c10D70,c11D70,c12D70,c13D70;
wire signed [4:0] c10D80,c11D80,c12D80,c13D80;
wire signed [4:0] c10D90,c11D90,c12D90,c13D90;
wire signed [4:0] c10DA0,c11DA0,c12DA0,c13DA0;
wire signed [4:0] c10DB0,c11DB0,c12DB0,c13DB0;
wire signed [4:0] c10DC0,c11DC0,c12DC0,c13DC0;
wire signed [4:0] c10DD0,c11DD0,c12DD0,c13DD0;
wire signed [4:0] c10001,c11001,c12001,c13001;
wire signed [4:0] c10011,c11011,c12011,c13011;
wire signed [4:0] c10021,c11021,c12021,c13021;
wire signed [4:0] c10031,c11031,c12031,c13031;
wire signed [4:0] c10041,c11041,c12041,c13041;
wire signed [4:0] c10051,c11051,c12051,c13051;
wire signed [4:0] c10061,c11061,c12061,c13061;
wire signed [4:0] c10071,c11071,c12071,c13071;
wire signed [4:0] c10081,c11081,c12081,c13081;
wire signed [4:0] c10091,c11091,c12091,c13091;
wire signed [4:0] c100A1,c110A1,c120A1,c130A1;
wire signed [4:0] c100B1,c110B1,c120B1,c130B1;
wire signed [4:0] c100C1,c110C1,c120C1,c130C1;
wire signed [4:0] c100D1,c110D1,c120D1,c130D1;
wire signed [4:0] c10101,c11101,c12101,c13101;
wire signed [4:0] c10111,c11111,c12111,c13111;
wire signed [4:0] c10121,c11121,c12121,c13121;
wire signed [4:0] c10131,c11131,c12131,c13131;
wire signed [4:0] c10141,c11141,c12141,c13141;
wire signed [4:0] c10151,c11151,c12151,c13151;
wire signed [4:0] c10161,c11161,c12161,c13161;
wire signed [4:0] c10171,c11171,c12171,c13171;
wire signed [4:0] c10181,c11181,c12181,c13181;
wire signed [4:0] c10191,c11191,c12191,c13191;
wire signed [4:0] c101A1,c111A1,c121A1,c131A1;
wire signed [4:0] c101B1,c111B1,c121B1,c131B1;
wire signed [4:0] c101C1,c111C1,c121C1,c131C1;
wire signed [4:0] c101D1,c111D1,c121D1,c131D1;
wire signed [4:0] c10201,c11201,c12201,c13201;
wire signed [4:0] c10211,c11211,c12211,c13211;
wire signed [4:0] c10221,c11221,c12221,c13221;
wire signed [4:0] c10231,c11231,c12231,c13231;
wire signed [4:0] c10241,c11241,c12241,c13241;
wire signed [4:0] c10251,c11251,c12251,c13251;
wire signed [4:0] c10261,c11261,c12261,c13261;
wire signed [4:0] c10271,c11271,c12271,c13271;
wire signed [4:0] c10281,c11281,c12281,c13281;
wire signed [4:0] c10291,c11291,c12291,c13291;
wire signed [4:0] c102A1,c112A1,c122A1,c132A1;
wire signed [4:0] c102B1,c112B1,c122B1,c132B1;
wire signed [4:0] c102C1,c112C1,c122C1,c132C1;
wire signed [4:0] c102D1,c112D1,c122D1,c132D1;
wire signed [4:0] c10301,c11301,c12301,c13301;
wire signed [4:0] c10311,c11311,c12311,c13311;
wire signed [4:0] c10321,c11321,c12321,c13321;
wire signed [4:0] c10331,c11331,c12331,c13331;
wire signed [4:0] c10341,c11341,c12341,c13341;
wire signed [4:0] c10351,c11351,c12351,c13351;
wire signed [4:0] c10361,c11361,c12361,c13361;
wire signed [4:0] c10371,c11371,c12371,c13371;
wire signed [4:0] c10381,c11381,c12381,c13381;
wire signed [4:0] c10391,c11391,c12391,c13391;
wire signed [4:0] c103A1,c113A1,c123A1,c133A1;
wire signed [4:0] c103B1,c113B1,c123B1,c133B1;
wire signed [4:0] c103C1,c113C1,c123C1,c133C1;
wire signed [4:0] c103D1,c113D1,c123D1,c133D1;
wire signed [4:0] c10401,c11401,c12401,c13401;
wire signed [4:0] c10411,c11411,c12411,c13411;
wire signed [4:0] c10421,c11421,c12421,c13421;
wire signed [4:0] c10431,c11431,c12431,c13431;
wire signed [4:0] c10441,c11441,c12441,c13441;
wire signed [4:0] c10451,c11451,c12451,c13451;
wire signed [4:0] c10461,c11461,c12461,c13461;
wire signed [4:0] c10471,c11471,c12471,c13471;
wire signed [4:0] c10481,c11481,c12481,c13481;
wire signed [4:0] c10491,c11491,c12491,c13491;
wire signed [4:0] c104A1,c114A1,c124A1,c134A1;
wire signed [4:0] c104B1,c114B1,c124B1,c134B1;
wire signed [4:0] c104C1,c114C1,c124C1,c134C1;
wire signed [4:0] c104D1,c114D1,c124D1,c134D1;
wire signed [4:0] c10501,c11501,c12501,c13501;
wire signed [4:0] c10511,c11511,c12511,c13511;
wire signed [4:0] c10521,c11521,c12521,c13521;
wire signed [4:0] c10531,c11531,c12531,c13531;
wire signed [4:0] c10541,c11541,c12541,c13541;
wire signed [4:0] c10551,c11551,c12551,c13551;
wire signed [4:0] c10561,c11561,c12561,c13561;
wire signed [4:0] c10571,c11571,c12571,c13571;
wire signed [4:0] c10581,c11581,c12581,c13581;
wire signed [4:0] c10591,c11591,c12591,c13591;
wire signed [4:0] c105A1,c115A1,c125A1,c135A1;
wire signed [4:0] c105B1,c115B1,c125B1,c135B1;
wire signed [4:0] c105C1,c115C1,c125C1,c135C1;
wire signed [4:0] c105D1,c115D1,c125D1,c135D1;
wire signed [4:0] c10601,c11601,c12601,c13601;
wire signed [4:0] c10611,c11611,c12611,c13611;
wire signed [4:0] c10621,c11621,c12621,c13621;
wire signed [4:0] c10631,c11631,c12631,c13631;
wire signed [4:0] c10641,c11641,c12641,c13641;
wire signed [4:0] c10651,c11651,c12651,c13651;
wire signed [4:0] c10661,c11661,c12661,c13661;
wire signed [4:0] c10671,c11671,c12671,c13671;
wire signed [4:0] c10681,c11681,c12681,c13681;
wire signed [4:0] c10691,c11691,c12691,c13691;
wire signed [4:0] c106A1,c116A1,c126A1,c136A1;
wire signed [4:0] c106B1,c116B1,c126B1,c136B1;
wire signed [4:0] c106C1,c116C1,c126C1,c136C1;
wire signed [4:0] c106D1,c116D1,c126D1,c136D1;
wire signed [4:0] c10701,c11701,c12701,c13701;
wire signed [4:0] c10711,c11711,c12711,c13711;
wire signed [4:0] c10721,c11721,c12721,c13721;
wire signed [4:0] c10731,c11731,c12731,c13731;
wire signed [4:0] c10741,c11741,c12741,c13741;
wire signed [4:0] c10751,c11751,c12751,c13751;
wire signed [4:0] c10761,c11761,c12761,c13761;
wire signed [4:0] c10771,c11771,c12771,c13771;
wire signed [4:0] c10781,c11781,c12781,c13781;
wire signed [4:0] c10791,c11791,c12791,c13791;
wire signed [4:0] c107A1,c117A1,c127A1,c137A1;
wire signed [4:0] c107B1,c117B1,c127B1,c137B1;
wire signed [4:0] c107C1,c117C1,c127C1,c137C1;
wire signed [4:0] c107D1,c117D1,c127D1,c137D1;
wire signed [4:0] c10801,c11801,c12801,c13801;
wire signed [4:0] c10811,c11811,c12811,c13811;
wire signed [4:0] c10821,c11821,c12821,c13821;
wire signed [4:0] c10831,c11831,c12831,c13831;
wire signed [4:0] c10841,c11841,c12841,c13841;
wire signed [4:0] c10851,c11851,c12851,c13851;
wire signed [4:0] c10861,c11861,c12861,c13861;
wire signed [4:0] c10871,c11871,c12871,c13871;
wire signed [4:0] c10881,c11881,c12881,c13881;
wire signed [4:0] c10891,c11891,c12891,c13891;
wire signed [4:0] c108A1,c118A1,c128A1,c138A1;
wire signed [4:0] c108B1,c118B1,c128B1,c138B1;
wire signed [4:0] c108C1,c118C1,c128C1,c138C1;
wire signed [4:0] c108D1,c118D1,c128D1,c138D1;
wire signed [4:0] c10901,c11901,c12901,c13901;
wire signed [4:0] c10911,c11911,c12911,c13911;
wire signed [4:0] c10921,c11921,c12921,c13921;
wire signed [4:0] c10931,c11931,c12931,c13931;
wire signed [4:0] c10941,c11941,c12941,c13941;
wire signed [4:0] c10951,c11951,c12951,c13951;
wire signed [4:0] c10961,c11961,c12961,c13961;
wire signed [4:0] c10971,c11971,c12971,c13971;
wire signed [4:0] c10981,c11981,c12981,c13981;
wire signed [4:0] c10991,c11991,c12991,c13991;
wire signed [4:0] c109A1,c119A1,c129A1,c139A1;
wire signed [4:0] c109B1,c119B1,c129B1,c139B1;
wire signed [4:0] c109C1,c119C1,c129C1,c139C1;
wire signed [4:0] c109D1,c119D1,c129D1,c139D1;
wire signed [4:0] c10A01,c11A01,c12A01,c13A01;
wire signed [4:0] c10A11,c11A11,c12A11,c13A11;
wire signed [4:0] c10A21,c11A21,c12A21,c13A21;
wire signed [4:0] c10A31,c11A31,c12A31,c13A31;
wire signed [4:0] c10A41,c11A41,c12A41,c13A41;
wire signed [4:0] c10A51,c11A51,c12A51,c13A51;
wire signed [4:0] c10A61,c11A61,c12A61,c13A61;
wire signed [4:0] c10A71,c11A71,c12A71,c13A71;
wire signed [4:0] c10A81,c11A81,c12A81,c13A81;
wire signed [4:0] c10A91,c11A91,c12A91,c13A91;
wire signed [4:0] c10AA1,c11AA1,c12AA1,c13AA1;
wire signed [4:0] c10AB1,c11AB1,c12AB1,c13AB1;
wire signed [4:0] c10AC1,c11AC1,c12AC1,c13AC1;
wire signed [4:0] c10AD1,c11AD1,c12AD1,c13AD1;
wire signed [4:0] c10B01,c11B01,c12B01,c13B01;
wire signed [4:0] c10B11,c11B11,c12B11,c13B11;
wire signed [4:0] c10B21,c11B21,c12B21,c13B21;
wire signed [4:0] c10B31,c11B31,c12B31,c13B31;
wire signed [4:0] c10B41,c11B41,c12B41,c13B41;
wire signed [4:0] c10B51,c11B51,c12B51,c13B51;
wire signed [4:0] c10B61,c11B61,c12B61,c13B61;
wire signed [4:0] c10B71,c11B71,c12B71,c13B71;
wire signed [4:0] c10B81,c11B81,c12B81,c13B81;
wire signed [4:0] c10B91,c11B91,c12B91,c13B91;
wire signed [4:0] c10BA1,c11BA1,c12BA1,c13BA1;
wire signed [4:0] c10BB1,c11BB1,c12BB1,c13BB1;
wire signed [4:0] c10BC1,c11BC1,c12BC1,c13BC1;
wire signed [4:0] c10BD1,c11BD1,c12BD1,c13BD1;
wire signed [4:0] c10C01,c11C01,c12C01,c13C01;
wire signed [4:0] c10C11,c11C11,c12C11,c13C11;
wire signed [4:0] c10C21,c11C21,c12C21,c13C21;
wire signed [4:0] c10C31,c11C31,c12C31,c13C31;
wire signed [4:0] c10C41,c11C41,c12C41,c13C41;
wire signed [4:0] c10C51,c11C51,c12C51,c13C51;
wire signed [4:0] c10C61,c11C61,c12C61,c13C61;
wire signed [4:0] c10C71,c11C71,c12C71,c13C71;
wire signed [4:0] c10C81,c11C81,c12C81,c13C81;
wire signed [4:0] c10C91,c11C91,c12C91,c13C91;
wire signed [4:0] c10CA1,c11CA1,c12CA1,c13CA1;
wire signed [4:0] c10CB1,c11CB1,c12CB1,c13CB1;
wire signed [4:0] c10CC1,c11CC1,c12CC1,c13CC1;
wire signed [4:0] c10CD1,c11CD1,c12CD1,c13CD1;
wire signed [4:0] c10D01,c11D01,c12D01,c13D01;
wire signed [4:0] c10D11,c11D11,c12D11,c13D11;
wire signed [4:0] c10D21,c11D21,c12D21,c13D21;
wire signed [4:0] c10D31,c11D31,c12D31,c13D31;
wire signed [4:0] c10D41,c11D41,c12D41,c13D41;
wire signed [4:0] c10D51,c11D51,c12D51,c13D51;
wire signed [4:0] c10D61,c11D61,c12D61,c13D61;
wire signed [4:0] c10D71,c11D71,c12D71,c13D71;
wire signed [4:0] c10D81,c11D81,c12D81,c13D81;
wire signed [4:0] c10D91,c11D91,c12D91,c13D91;
wire signed [4:0] c10DA1,c11DA1,c12DA1,c13DA1;
wire signed [4:0] c10DB1,c11DB1,c12DB1,c13DB1;
wire signed [4:0] c10DC1,c11DC1,c12DC1,c13DC1;
wire signed [4:0] c10DD1,c11DD1,c12DD1,c13DD1;
wire signed [4:0] c10002,c11002,c12002,c13002;
wire signed [4:0] c10012,c11012,c12012,c13012;
wire signed [4:0] c10022,c11022,c12022,c13022;
wire signed [4:0] c10032,c11032,c12032,c13032;
wire signed [4:0] c10042,c11042,c12042,c13042;
wire signed [4:0] c10052,c11052,c12052,c13052;
wire signed [4:0] c10062,c11062,c12062,c13062;
wire signed [4:0] c10072,c11072,c12072,c13072;
wire signed [4:0] c10082,c11082,c12082,c13082;
wire signed [4:0] c10092,c11092,c12092,c13092;
wire signed [4:0] c100A2,c110A2,c120A2,c130A2;
wire signed [4:0] c100B2,c110B2,c120B2,c130B2;
wire signed [4:0] c100C2,c110C2,c120C2,c130C2;
wire signed [4:0] c100D2,c110D2,c120D2,c130D2;
wire signed [4:0] c10102,c11102,c12102,c13102;
wire signed [4:0] c10112,c11112,c12112,c13112;
wire signed [4:0] c10122,c11122,c12122,c13122;
wire signed [4:0] c10132,c11132,c12132,c13132;
wire signed [4:0] c10142,c11142,c12142,c13142;
wire signed [4:0] c10152,c11152,c12152,c13152;
wire signed [4:0] c10162,c11162,c12162,c13162;
wire signed [4:0] c10172,c11172,c12172,c13172;
wire signed [4:0] c10182,c11182,c12182,c13182;
wire signed [4:0] c10192,c11192,c12192,c13192;
wire signed [4:0] c101A2,c111A2,c121A2,c131A2;
wire signed [4:0] c101B2,c111B2,c121B2,c131B2;
wire signed [4:0] c101C2,c111C2,c121C2,c131C2;
wire signed [4:0] c101D2,c111D2,c121D2,c131D2;
wire signed [4:0] c10202,c11202,c12202,c13202;
wire signed [4:0] c10212,c11212,c12212,c13212;
wire signed [4:0] c10222,c11222,c12222,c13222;
wire signed [4:0] c10232,c11232,c12232,c13232;
wire signed [4:0] c10242,c11242,c12242,c13242;
wire signed [4:0] c10252,c11252,c12252,c13252;
wire signed [4:0] c10262,c11262,c12262,c13262;
wire signed [4:0] c10272,c11272,c12272,c13272;
wire signed [4:0] c10282,c11282,c12282,c13282;
wire signed [4:0] c10292,c11292,c12292,c13292;
wire signed [4:0] c102A2,c112A2,c122A2,c132A2;
wire signed [4:0] c102B2,c112B2,c122B2,c132B2;
wire signed [4:0] c102C2,c112C2,c122C2,c132C2;
wire signed [4:0] c102D2,c112D2,c122D2,c132D2;
wire signed [4:0] c10302,c11302,c12302,c13302;
wire signed [4:0] c10312,c11312,c12312,c13312;
wire signed [4:0] c10322,c11322,c12322,c13322;
wire signed [4:0] c10332,c11332,c12332,c13332;
wire signed [4:0] c10342,c11342,c12342,c13342;
wire signed [4:0] c10352,c11352,c12352,c13352;
wire signed [4:0] c10362,c11362,c12362,c13362;
wire signed [4:0] c10372,c11372,c12372,c13372;
wire signed [4:0] c10382,c11382,c12382,c13382;
wire signed [4:0] c10392,c11392,c12392,c13392;
wire signed [4:0] c103A2,c113A2,c123A2,c133A2;
wire signed [4:0] c103B2,c113B2,c123B2,c133B2;
wire signed [4:0] c103C2,c113C2,c123C2,c133C2;
wire signed [4:0] c103D2,c113D2,c123D2,c133D2;
wire signed [4:0] c10402,c11402,c12402,c13402;
wire signed [4:0] c10412,c11412,c12412,c13412;
wire signed [4:0] c10422,c11422,c12422,c13422;
wire signed [4:0] c10432,c11432,c12432,c13432;
wire signed [4:0] c10442,c11442,c12442,c13442;
wire signed [4:0] c10452,c11452,c12452,c13452;
wire signed [4:0] c10462,c11462,c12462,c13462;
wire signed [4:0] c10472,c11472,c12472,c13472;
wire signed [4:0] c10482,c11482,c12482,c13482;
wire signed [4:0] c10492,c11492,c12492,c13492;
wire signed [4:0] c104A2,c114A2,c124A2,c134A2;
wire signed [4:0] c104B2,c114B2,c124B2,c134B2;
wire signed [4:0] c104C2,c114C2,c124C2,c134C2;
wire signed [4:0] c104D2,c114D2,c124D2,c134D2;
wire signed [4:0] c10502,c11502,c12502,c13502;
wire signed [4:0] c10512,c11512,c12512,c13512;
wire signed [4:0] c10522,c11522,c12522,c13522;
wire signed [4:0] c10532,c11532,c12532,c13532;
wire signed [4:0] c10542,c11542,c12542,c13542;
wire signed [4:0] c10552,c11552,c12552,c13552;
wire signed [4:0] c10562,c11562,c12562,c13562;
wire signed [4:0] c10572,c11572,c12572,c13572;
wire signed [4:0] c10582,c11582,c12582,c13582;
wire signed [4:0] c10592,c11592,c12592,c13592;
wire signed [4:0] c105A2,c115A2,c125A2,c135A2;
wire signed [4:0] c105B2,c115B2,c125B2,c135B2;
wire signed [4:0] c105C2,c115C2,c125C2,c135C2;
wire signed [4:0] c105D2,c115D2,c125D2,c135D2;
wire signed [4:0] c10602,c11602,c12602,c13602;
wire signed [4:0] c10612,c11612,c12612,c13612;
wire signed [4:0] c10622,c11622,c12622,c13622;
wire signed [4:0] c10632,c11632,c12632,c13632;
wire signed [4:0] c10642,c11642,c12642,c13642;
wire signed [4:0] c10652,c11652,c12652,c13652;
wire signed [4:0] c10662,c11662,c12662,c13662;
wire signed [4:0] c10672,c11672,c12672,c13672;
wire signed [4:0] c10682,c11682,c12682,c13682;
wire signed [4:0] c10692,c11692,c12692,c13692;
wire signed [4:0] c106A2,c116A2,c126A2,c136A2;
wire signed [4:0] c106B2,c116B2,c126B2,c136B2;
wire signed [4:0] c106C2,c116C2,c126C2,c136C2;
wire signed [4:0] c106D2,c116D2,c126D2,c136D2;
wire signed [4:0] c10702,c11702,c12702,c13702;
wire signed [4:0] c10712,c11712,c12712,c13712;
wire signed [4:0] c10722,c11722,c12722,c13722;
wire signed [4:0] c10732,c11732,c12732,c13732;
wire signed [4:0] c10742,c11742,c12742,c13742;
wire signed [4:0] c10752,c11752,c12752,c13752;
wire signed [4:0] c10762,c11762,c12762,c13762;
wire signed [4:0] c10772,c11772,c12772,c13772;
wire signed [4:0] c10782,c11782,c12782,c13782;
wire signed [4:0] c10792,c11792,c12792,c13792;
wire signed [4:0] c107A2,c117A2,c127A2,c137A2;
wire signed [4:0] c107B2,c117B2,c127B2,c137B2;
wire signed [4:0] c107C2,c117C2,c127C2,c137C2;
wire signed [4:0] c107D2,c117D2,c127D2,c137D2;
wire signed [4:0] c10802,c11802,c12802,c13802;
wire signed [4:0] c10812,c11812,c12812,c13812;
wire signed [4:0] c10822,c11822,c12822,c13822;
wire signed [4:0] c10832,c11832,c12832,c13832;
wire signed [4:0] c10842,c11842,c12842,c13842;
wire signed [4:0] c10852,c11852,c12852,c13852;
wire signed [4:0] c10862,c11862,c12862,c13862;
wire signed [4:0] c10872,c11872,c12872,c13872;
wire signed [4:0] c10882,c11882,c12882,c13882;
wire signed [4:0] c10892,c11892,c12892,c13892;
wire signed [4:0] c108A2,c118A2,c128A2,c138A2;
wire signed [4:0] c108B2,c118B2,c128B2,c138B2;
wire signed [4:0] c108C2,c118C2,c128C2,c138C2;
wire signed [4:0] c108D2,c118D2,c128D2,c138D2;
wire signed [4:0] c10902,c11902,c12902,c13902;
wire signed [4:0] c10912,c11912,c12912,c13912;
wire signed [4:0] c10922,c11922,c12922,c13922;
wire signed [4:0] c10932,c11932,c12932,c13932;
wire signed [4:0] c10942,c11942,c12942,c13942;
wire signed [4:0] c10952,c11952,c12952,c13952;
wire signed [4:0] c10962,c11962,c12962,c13962;
wire signed [4:0] c10972,c11972,c12972,c13972;
wire signed [4:0] c10982,c11982,c12982,c13982;
wire signed [4:0] c10992,c11992,c12992,c13992;
wire signed [4:0] c109A2,c119A2,c129A2,c139A2;
wire signed [4:0] c109B2,c119B2,c129B2,c139B2;
wire signed [4:0] c109C2,c119C2,c129C2,c139C2;
wire signed [4:0] c109D2,c119D2,c129D2,c139D2;
wire signed [4:0] c10A02,c11A02,c12A02,c13A02;
wire signed [4:0] c10A12,c11A12,c12A12,c13A12;
wire signed [4:0] c10A22,c11A22,c12A22,c13A22;
wire signed [4:0] c10A32,c11A32,c12A32,c13A32;
wire signed [4:0] c10A42,c11A42,c12A42,c13A42;
wire signed [4:0] c10A52,c11A52,c12A52,c13A52;
wire signed [4:0] c10A62,c11A62,c12A62,c13A62;
wire signed [4:0] c10A72,c11A72,c12A72,c13A72;
wire signed [4:0] c10A82,c11A82,c12A82,c13A82;
wire signed [4:0] c10A92,c11A92,c12A92,c13A92;
wire signed [4:0] c10AA2,c11AA2,c12AA2,c13AA2;
wire signed [4:0] c10AB2,c11AB2,c12AB2,c13AB2;
wire signed [4:0] c10AC2,c11AC2,c12AC2,c13AC2;
wire signed [4:0] c10AD2,c11AD2,c12AD2,c13AD2;
wire signed [4:0] c10B02,c11B02,c12B02,c13B02;
wire signed [4:0] c10B12,c11B12,c12B12,c13B12;
wire signed [4:0] c10B22,c11B22,c12B22,c13B22;
wire signed [4:0] c10B32,c11B32,c12B32,c13B32;
wire signed [4:0] c10B42,c11B42,c12B42,c13B42;
wire signed [4:0] c10B52,c11B52,c12B52,c13B52;
wire signed [4:0] c10B62,c11B62,c12B62,c13B62;
wire signed [4:0] c10B72,c11B72,c12B72,c13B72;
wire signed [4:0] c10B82,c11B82,c12B82,c13B82;
wire signed [4:0] c10B92,c11B92,c12B92,c13B92;
wire signed [4:0] c10BA2,c11BA2,c12BA2,c13BA2;
wire signed [4:0] c10BB2,c11BB2,c12BB2,c13BB2;
wire signed [4:0] c10BC2,c11BC2,c12BC2,c13BC2;
wire signed [4:0] c10BD2,c11BD2,c12BD2,c13BD2;
wire signed [4:0] c10C02,c11C02,c12C02,c13C02;
wire signed [4:0] c10C12,c11C12,c12C12,c13C12;
wire signed [4:0] c10C22,c11C22,c12C22,c13C22;
wire signed [4:0] c10C32,c11C32,c12C32,c13C32;
wire signed [4:0] c10C42,c11C42,c12C42,c13C42;
wire signed [4:0] c10C52,c11C52,c12C52,c13C52;
wire signed [4:0] c10C62,c11C62,c12C62,c13C62;
wire signed [4:0] c10C72,c11C72,c12C72,c13C72;
wire signed [4:0] c10C82,c11C82,c12C82,c13C82;
wire signed [4:0] c10C92,c11C92,c12C92,c13C92;
wire signed [4:0] c10CA2,c11CA2,c12CA2,c13CA2;
wire signed [4:0] c10CB2,c11CB2,c12CB2,c13CB2;
wire signed [4:0] c10CC2,c11CC2,c12CC2,c13CC2;
wire signed [4:0] c10CD2,c11CD2,c12CD2,c13CD2;
wire signed [4:0] c10D02,c11D02,c12D02,c13D02;
wire signed [4:0] c10D12,c11D12,c12D12,c13D12;
wire signed [4:0] c10D22,c11D22,c12D22,c13D22;
wire signed [4:0] c10D32,c11D32,c12D32,c13D32;
wire signed [4:0] c10D42,c11D42,c12D42,c13D42;
wire signed [4:0] c10D52,c11D52,c12D52,c13D52;
wire signed [4:0] c10D62,c11D62,c12D62,c13D62;
wire signed [4:0] c10D72,c11D72,c12D72,c13D72;
wire signed [4:0] c10D82,c11D82,c12D82,c13D82;
wire signed [4:0] c10D92,c11D92,c12D92,c13D92;
wire signed [4:0] c10DA2,c11DA2,c12DA2,c13DA2;
wire signed [4:0] c10DB2,c11DB2,c12DB2,c13DB2;
wire signed [4:0] c10DC2,c11DC2,c12DC2,c13DC2;
wire signed [4:0] c10DD2,c11DD2,c12DD2,c13DD2;
wire signed [4:0] c10003,c11003,c12003,c13003;
wire signed [4:0] c10013,c11013,c12013,c13013;
wire signed [4:0] c10023,c11023,c12023,c13023;
wire signed [4:0] c10033,c11033,c12033,c13033;
wire signed [4:0] c10043,c11043,c12043,c13043;
wire signed [4:0] c10053,c11053,c12053,c13053;
wire signed [4:0] c10063,c11063,c12063,c13063;
wire signed [4:0] c10073,c11073,c12073,c13073;
wire signed [4:0] c10083,c11083,c12083,c13083;
wire signed [4:0] c10093,c11093,c12093,c13093;
wire signed [4:0] c100A3,c110A3,c120A3,c130A3;
wire signed [4:0] c100B3,c110B3,c120B3,c130B3;
wire signed [4:0] c100C3,c110C3,c120C3,c130C3;
wire signed [4:0] c100D3,c110D3,c120D3,c130D3;
wire signed [4:0] c10103,c11103,c12103,c13103;
wire signed [4:0] c10113,c11113,c12113,c13113;
wire signed [4:0] c10123,c11123,c12123,c13123;
wire signed [4:0] c10133,c11133,c12133,c13133;
wire signed [4:0] c10143,c11143,c12143,c13143;
wire signed [4:0] c10153,c11153,c12153,c13153;
wire signed [4:0] c10163,c11163,c12163,c13163;
wire signed [4:0] c10173,c11173,c12173,c13173;
wire signed [4:0] c10183,c11183,c12183,c13183;
wire signed [4:0] c10193,c11193,c12193,c13193;
wire signed [4:0] c101A3,c111A3,c121A3,c131A3;
wire signed [4:0] c101B3,c111B3,c121B3,c131B3;
wire signed [4:0] c101C3,c111C3,c121C3,c131C3;
wire signed [4:0] c101D3,c111D3,c121D3,c131D3;
wire signed [4:0] c10203,c11203,c12203,c13203;
wire signed [4:0] c10213,c11213,c12213,c13213;
wire signed [4:0] c10223,c11223,c12223,c13223;
wire signed [4:0] c10233,c11233,c12233,c13233;
wire signed [4:0] c10243,c11243,c12243,c13243;
wire signed [4:0] c10253,c11253,c12253,c13253;
wire signed [4:0] c10263,c11263,c12263,c13263;
wire signed [4:0] c10273,c11273,c12273,c13273;
wire signed [4:0] c10283,c11283,c12283,c13283;
wire signed [4:0] c10293,c11293,c12293,c13293;
wire signed [4:0] c102A3,c112A3,c122A3,c132A3;
wire signed [4:0] c102B3,c112B3,c122B3,c132B3;
wire signed [4:0] c102C3,c112C3,c122C3,c132C3;
wire signed [4:0] c102D3,c112D3,c122D3,c132D3;
wire signed [4:0] c10303,c11303,c12303,c13303;
wire signed [4:0] c10313,c11313,c12313,c13313;
wire signed [4:0] c10323,c11323,c12323,c13323;
wire signed [4:0] c10333,c11333,c12333,c13333;
wire signed [4:0] c10343,c11343,c12343,c13343;
wire signed [4:0] c10353,c11353,c12353,c13353;
wire signed [4:0] c10363,c11363,c12363,c13363;
wire signed [4:0] c10373,c11373,c12373,c13373;
wire signed [4:0] c10383,c11383,c12383,c13383;
wire signed [4:0] c10393,c11393,c12393,c13393;
wire signed [4:0] c103A3,c113A3,c123A3,c133A3;
wire signed [4:0] c103B3,c113B3,c123B3,c133B3;
wire signed [4:0] c103C3,c113C3,c123C3,c133C3;
wire signed [4:0] c103D3,c113D3,c123D3,c133D3;
wire signed [4:0] c10403,c11403,c12403,c13403;
wire signed [4:0] c10413,c11413,c12413,c13413;
wire signed [4:0] c10423,c11423,c12423,c13423;
wire signed [4:0] c10433,c11433,c12433,c13433;
wire signed [4:0] c10443,c11443,c12443,c13443;
wire signed [4:0] c10453,c11453,c12453,c13453;
wire signed [4:0] c10463,c11463,c12463,c13463;
wire signed [4:0] c10473,c11473,c12473,c13473;
wire signed [4:0] c10483,c11483,c12483,c13483;
wire signed [4:0] c10493,c11493,c12493,c13493;
wire signed [4:0] c104A3,c114A3,c124A3,c134A3;
wire signed [4:0] c104B3,c114B3,c124B3,c134B3;
wire signed [4:0] c104C3,c114C3,c124C3,c134C3;
wire signed [4:0] c104D3,c114D3,c124D3,c134D3;
wire signed [4:0] c10503,c11503,c12503,c13503;
wire signed [4:0] c10513,c11513,c12513,c13513;
wire signed [4:0] c10523,c11523,c12523,c13523;
wire signed [4:0] c10533,c11533,c12533,c13533;
wire signed [4:0] c10543,c11543,c12543,c13543;
wire signed [4:0] c10553,c11553,c12553,c13553;
wire signed [4:0] c10563,c11563,c12563,c13563;
wire signed [4:0] c10573,c11573,c12573,c13573;
wire signed [4:0] c10583,c11583,c12583,c13583;
wire signed [4:0] c10593,c11593,c12593,c13593;
wire signed [4:0] c105A3,c115A3,c125A3,c135A3;
wire signed [4:0] c105B3,c115B3,c125B3,c135B3;
wire signed [4:0] c105C3,c115C3,c125C3,c135C3;
wire signed [4:0] c105D3,c115D3,c125D3,c135D3;
wire signed [4:0] c10603,c11603,c12603,c13603;
wire signed [4:0] c10613,c11613,c12613,c13613;
wire signed [4:0] c10623,c11623,c12623,c13623;
wire signed [4:0] c10633,c11633,c12633,c13633;
wire signed [4:0] c10643,c11643,c12643,c13643;
wire signed [4:0] c10653,c11653,c12653,c13653;
wire signed [4:0] c10663,c11663,c12663,c13663;
wire signed [4:0] c10673,c11673,c12673,c13673;
wire signed [4:0] c10683,c11683,c12683,c13683;
wire signed [4:0] c10693,c11693,c12693,c13693;
wire signed [4:0] c106A3,c116A3,c126A3,c136A3;
wire signed [4:0] c106B3,c116B3,c126B3,c136B3;
wire signed [4:0] c106C3,c116C3,c126C3,c136C3;
wire signed [4:0] c106D3,c116D3,c126D3,c136D3;
wire signed [4:0] c10703,c11703,c12703,c13703;
wire signed [4:0] c10713,c11713,c12713,c13713;
wire signed [4:0] c10723,c11723,c12723,c13723;
wire signed [4:0] c10733,c11733,c12733,c13733;
wire signed [4:0] c10743,c11743,c12743,c13743;
wire signed [4:0] c10753,c11753,c12753,c13753;
wire signed [4:0] c10763,c11763,c12763,c13763;
wire signed [4:0] c10773,c11773,c12773,c13773;
wire signed [4:0] c10783,c11783,c12783,c13783;
wire signed [4:0] c10793,c11793,c12793,c13793;
wire signed [4:0] c107A3,c117A3,c127A3,c137A3;
wire signed [4:0] c107B3,c117B3,c127B3,c137B3;
wire signed [4:0] c107C3,c117C3,c127C3,c137C3;
wire signed [4:0] c107D3,c117D3,c127D3,c137D3;
wire signed [4:0] c10803,c11803,c12803,c13803;
wire signed [4:0] c10813,c11813,c12813,c13813;
wire signed [4:0] c10823,c11823,c12823,c13823;
wire signed [4:0] c10833,c11833,c12833,c13833;
wire signed [4:0] c10843,c11843,c12843,c13843;
wire signed [4:0] c10853,c11853,c12853,c13853;
wire signed [4:0] c10863,c11863,c12863,c13863;
wire signed [4:0] c10873,c11873,c12873,c13873;
wire signed [4:0] c10883,c11883,c12883,c13883;
wire signed [4:0] c10893,c11893,c12893,c13893;
wire signed [4:0] c108A3,c118A3,c128A3,c138A3;
wire signed [4:0] c108B3,c118B3,c128B3,c138B3;
wire signed [4:0] c108C3,c118C3,c128C3,c138C3;
wire signed [4:0] c108D3,c118D3,c128D3,c138D3;
wire signed [4:0] c10903,c11903,c12903,c13903;
wire signed [4:0] c10913,c11913,c12913,c13913;
wire signed [4:0] c10923,c11923,c12923,c13923;
wire signed [4:0] c10933,c11933,c12933,c13933;
wire signed [4:0] c10943,c11943,c12943,c13943;
wire signed [4:0] c10953,c11953,c12953,c13953;
wire signed [4:0] c10963,c11963,c12963,c13963;
wire signed [4:0] c10973,c11973,c12973,c13973;
wire signed [4:0] c10983,c11983,c12983,c13983;
wire signed [4:0] c10993,c11993,c12993,c13993;
wire signed [4:0] c109A3,c119A3,c129A3,c139A3;
wire signed [4:0] c109B3,c119B3,c129B3,c139B3;
wire signed [4:0] c109C3,c119C3,c129C3,c139C3;
wire signed [4:0] c109D3,c119D3,c129D3,c139D3;
wire signed [4:0] c10A03,c11A03,c12A03,c13A03;
wire signed [4:0] c10A13,c11A13,c12A13,c13A13;
wire signed [4:0] c10A23,c11A23,c12A23,c13A23;
wire signed [4:0] c10A33,c11A33,c12A33,c13A33;
wire signed [4:0] c10A43,c11A43,c12A43,c13A43;
wire signed [4:0] c10A53,c11A53,c12A53,c13A53;
wire signed [4:0] c10A63,c11A63,c12A63,c13A63;
wire signed [4:0] c10A73,c11A73,c12A73,c13A73;
wire signed [4:0] c10A83,c11A83,c12A83,c13A83;
wire signed [4:0] c10A93,c11A93,c12A93,c13A93;
wire signed [4:0] c10AA3,c11AA3,c12AA3,c13AA3;
wire signed [4:0] c10AB3,c11AB3,c12AB3,c13AB3;
wire signed [4:0] c10AC3,c11AC3,c12AC3,c13AC3;
wire signed [4:0] c10AD3,c11AD3,c12AD3,c13AD3;
wire signed [4:0] c10B03,c11B03,c12B03,c13B03;
wire signed [4:0] c10B13,c11B13,c12B13,c13B13;
wire signed [4:0] c10B23,c11B23,c12B23,c13B23;
wire signed [4:0] c10B33,c11B33,c12B33,c13B33;
wire signed [4:0] c10B43,c11B43,c12B43,c13B43;
wire signed [4:0] c10B53,c11B53,c12B53,c13B53;
wire signed [4:0] c10B63,c11B63,c12B63,c13B63;
wire signed [4:0] c10B73,c11B73,c12B73,c13B73;
wire signed [4:0] c10B83,c11B83,c12B83,c13B83;
wire signed [4:0] c10B93,c11B93,c12B93,c13B93;
wire signed [4:0] c10BA3,c11BA3,c12BA3,c13BA3;
wire signed [4:0] c10BB3,c11BB3,c12BB3,c13BB3;
wire signed [4:0] c10BC3,c11BC3,c12BC3,c13BC3;
wire signed [4:0] c10BD3,c11BD3,c12BD3,c13BD3;
wire signed [4:0] c10C03,c11C03,c12C03,c13C03;
wire signed [4:0] c10C13,c11C13,c12C13,c13C13;
wire signed [4:0] c10C23,c11C23,c12C23,c13C23;
wire signed [4:0] c10C33,c11C33,c12C33,c13C33;
wire signed [4:0] c10C43,c11C43,c12C43,c13C43;
wire signed [4:0] c10C53,c11C53,c12C53,c13C53;
wire signed [4:0] c10C63,c11C63,c12C63,c13C63;
wire signed [4:0] c10C73,c11C73,c12C73,c13C73;
wire signed [4:0] c10C83,c11C83,c12C83,c13C83;
wire signed [4:0] c10C93,c11C93,c12C93,c13C93;
wire signed [4:0] c10CA3,c11CA3,c12CA3,c13CA3;
wire signed [4:0] c10CB3,c11CB3,c12CB3,c13CB3;
wire signed [4:0] c10CC3,c11CC3,c12CC3,c13CC3;
wire signed [4:0] c10CD3,c11CD3,c12CD3,c13CD3;
wire signed [4:0] c10D03,c11D03,c12D03,c13D03;
wire signed [4:0] c10D13,c11D13,c12D13,c13D13;
wire signed [4:0] c10D23,c11D23,c12D23,c13D23;
wire signed [4:0] c10D33,c11D33,c12D33,c13D33;
wire signed [4:0] c10D43,c11D43,c12D43,c13D43;
wire signed [4:0] c10D53,c11D53,c12D53,c13D53;
wire signed [4:0] c10D63,c11D63,c12D63,c13D63;
wire signed [4:0] c10D73,c11D73,c12D73,c13D73;
wire signed [4:0] c10D83,c11D83,c12D83,c13D83;
wire signed [4:0] c10D93,c11D93,c12D93,c13D93;
wire signed [4:0] c10DA3,c11DA3,c12DA3,c13DA3;
wire signed [4:0] c10DB3,c11DB3,c12DB3,c13DB3;
wire signed [4:0] c10DC3,c11DC3,c12DC3,c13DC3;
wire signed [4:0] c10DD3,c11DD3,c12DD3,c13DD3;
wire signed [4:0] c10004,c11004,c12004,c13004;
wire signed [4:0] c10014,c11014,c12014,c13014;
wire signed [4:0] c10024,c11024,c12024,c13024;
wire signed [4:0] c10034,c11034,c12034,c13034;
wire signed [4:0] c10044,c11044,c12044,c13044;
wire signed [4:0] c10054,c11054,c12054,c13054;
wire signed [4:0] c10064,c11064,c12064,c13064;
wire signed [4:0] c10074,c11074,c12074,c13074;
wire signed [4:0] c10084,c11084,c12084,c13084;
wire signed [4:0] c10094,c11094,c12094,c13094;
wire signed [4:0] c100A4,c110A4,c120A4,c130A4;
wire signed [4:0] c100B4,c110B4,c120B4,c130B4;
wire signed [4:0] c100C4,c110C4,c120C4,c130C4;
wire signed [4:0] c100D4,c110D4,c120D4,c130D4;
wire signed [4:0] c10104,c11104,c12104,c13104;
wire signed [4:0] c10114,c11114,c12114,c13114;
wire signed [4:0] c10124,c11124,c12124,c13124;
wire signed [4:0] c10134,c11134,c12134,c13134;
wire signed [4:0] c10144,c11144,c12144,c13144;
wire signed [4:0] c10154,c11154,c12154,c13154;
wire signed [4:0] c10164,c11164,c12164,c13164;
wire signed [4:0] c10174,c11174,c12174,c13174;
wire signed [4:0] c10184,c11184,c12184,c13184;
wire signed [4:0] c10194,c11194,c12194,c13194;
wire signed [4:0] c101A4,c111A4,c121A4,c131A4;
wire signed [4:0] c101B4,c111B4,c121B4,c131B4;
wire signed [4:0] c101C4,c111C4,c121C4,c131C4;
wire signed [4:0] c101D4,c111D4,c121D4,c131D4;
wire signed [4:0] c10204,c11204,c12204,c13204;
wire signed [4:0] c10214,c11214,c12214,c13214;
wire signed [4:0] c10224,c11224,c12224,c13224;
wire signed [4:0] c10234,c11234,c12234,c13234;
wire signed [4:0] c10244,c11244,c12244,c13244;
wire signed [4:0] c10254,c11254,c12254,c13254;
wire signed [4:0] c10264,c11264,c12264,c13264;
wire signed [4:0] c10274,c11274,c12274,c13274;
wire signed [4:0] c10284,c11284,c12284,c13284;
wire signed [4:0] c10294,c11294,c12294,c13294;
wire signed [4:0] c102A4,c112A4,c122A4,c132A4;
wire signed [4:0] c102B4,c112B4,c122B4,c132B4;
wire signed [4:0] c102C4,c112C4,c122C4,c132C4;
wire signed [4:0] c102D4,c112D4,c122D4,c132D4;
wire signed [4:0] c10304,c11304,c12304,c13304;
wire signed [4:0] c10314,c11314,c12314,c13314;
wire signed [4:0] c10324,c11324,c12324,c13324;
wire signed [4:0] c10334,c11334,c12334,c13334;
wire signed [4:0] c10344,c11344,c12344,c13344;
wire signed [4:0] c10354,c11354,c12354,c13354;
wire signed [4:0] c10364,c11364,c12364,c13364;
wire signed [4:0] c10374,c11374,c12374,c13374;
wire signed [4:0] c10384,c11384,c12384,c13384;
wire signed [4:0] c10394,c11394,c12394,c13394;
wire signed [4:0] c103A4,c113A4,c123A4,c133A4;
wire signed [4:0] c103B4,c113B4,c123B4,c133B4;
wire signed [4:0] c103C4,c113C4,c123C4,c133C4;
wire signed [4:0] c103D4,c113D4,c123D4,c133D4;
wire signed [4:0] c10404,c11404,c12404,c13404;
wire signed [4:0] c10414,c11414,c12414,c13414;
wire signed [4:0] c10424,c11424,c12424,c13424;
wire signed [4:0] c10434,c11434,c12434,c13434;
wire signed [4:0] c10444,c11444,c12444,c13444;
wire signed [4:0] c10454,c11454,c12454,c13454;
wire signed [4:0] c10464,c11464,c12464,c13464;
wire signed [4:0] c10474,c11474,c12474,c13474;
wire signed [4:0] c10484,c11484,c12484,c13484;
wire signed [4:0] c10494,c11494,c12494,c13494;
wire signed [4:0] c104A4,c114A4,c124A4,c134A4;
wire signed [4:0] c104B4,c114B4,c124B4,c134B4;
wire signed [4:0] c104C4,c114C4,c124C4,c134C4;
wire signed [4:0] c104D4,c114D4,c124D4,c134D4;
wire signed [4:0] c10504,c11504,c12504,c13504;
wire signed [4:0] c10514,c11514,c12514,c13514;
wire signed [4:0] c10524,c11524,c12524,c13524;
wire signed [4:0] c10534,c11534,c12534,c13534;
wire signed [4:0] c10544,c11544,c12544,c13544;
wire signed [4:0] c10554,c11554,c12554,c13554;
wire signed [4:0] c10564,c11564,c12564,c13564;
wire signed [4:0] c10574,c11574,c12574,c13574;
wire signed [4:0] c10584,c11584,c12584,c13584;
wire signed [4:0] c10594,c11594,c12594,c13594;
wire signed [4:0] c105A4,c115A4,c125A4,c135A4;
wire signed [4:0] c105B4,c115B4,c125B4,c135B4;
wire signed [4:0] c105C4,c115C4,c125C4,c135C4;
wire signed [4:0] c105D4,c115D4,c125D4,c135D4;
wire signed [4:0] c10604,c11604,c12604,c13604;
wire signed [4:0] c10614,c11614,c12614,c13614;
wire signed [4:0] c10624,c11624,c12624,c13624;
wire signed [4:0] c10634,c11634,c12634,c13634;
wire signed [4:0] c10644,c11644,c12644,c13644;
wire signed [4:0] c10654,c11654,c12654,c13654;
wire signed [4:0] c10664,c11664,c12664,c13664;
wire signed [4:0] c10674,c11674,c12674,c13674;
wire signed [4:0] c10684,c11684,c12684,c13684;
wire signed [4:0] c10694,c11694,c12694,c13694;
wire signed [4:0] c106A4,c116A4,c126A4,c136A4;
wire signed [4:0] c106B4,c116B4,c126B4,c136B4;
wire signed [4:0] c106C4,c116C4,c126C4,c136C4;
wire signed [4:0] c106D4,c116D4,c126D4,c136D4;
wire signed [4:0] c10704,c11704,c12704,c13704;
wire signed [4:0] c10714,c11714,c12714,c13714;
wire signed [4:0] c10724,c11724,c12724,c13724;
wire signed [4:0] c10734,c11734,c12734,c13734;
wire signed [4:0] c10744,c11744,c12744,c13744;
wire signed [4:0] c10754,c11754,c12754,c13754;
wire signed [4:0] c10764,c11764,c12764,c13764;
wire signed [4:0] c10774,c11774,c12774,c13774;
wire signed [4:0] c10784,c11784,c12784,c13784;
wire signed [4:0] c10794,c11794,c12794,c13794;
wire signed [4:0] c107A4,c117A4,c127A4,c137A4;
wire signed [4:0] c107B4,c117B4,c127B4,c137B4;
wire signed [4:0] c107C4,c117C4,c127C4,c137C4;
wire signed [4:0] c107D4,c117D4,c127D4,c137D4;
wire signed [4:0] c10804,c11804,c12804,c13804;
wire signed [4:0] c10814,c11814,c12814,c13814;
wire signed [4:0] c10824,c11824,c12824,c13824;
wire signed [4:0] c10834,c11834,c12834,c13834;
wire signed [4:0] c10844,c11844,c12844,c13844;
wire signed [4:0] c10854,c11854,c12854,c13854;
wire signed [4:0] c10864,c11864,c12864,c13864;
wire signed [4:0] c10874,c11874,c12874,c13874;
wire signed [4:0] c10884,c11884,c12884,c13884;
wire signed [4:0] c10894,c11894,c12894,c13894;
wire signed [4:0] c108A4,c118A4,c128A4,c138A4;
wire signed [4:0] c108B4,c118B4,c128B4,c138B4;
wire signed [4:0] c108C4,c118C4,c128C4,c138C4;
wire signed [4:0] c108D4,c118D4,c128D4,c138D4;
wire signed [4:0] c10904,c11904,c12904,c13904;
wire signed [4:0] c10914,c11914,c12914,c13914;
wire signed [4:0] c10924,c11924,c12924,c13924;
wire signed [4:0] c10934,c11934,c12934,c13934;
wire signed [4:0] c10944,c11944,c12944,c13944;
wire signed [4:0] c10954,c11954,c12954,c13954;
wire signed [4:0] c10964,c11964,c12964,c13964;
wire signed [4:0] c10974,c11974,c12974,c13974;
wire signed [4:0] c10984,c11984,c12984,c13984;
wire signed [4:0] c10994,c11994,c12994,c13994;
wire signed [4:0] c109A4,c119A4,c129A4,c139A4;
wire signed [4:0] c109B4,c119B4,c129B4,c139B4;
wire signed [4:0] c109C4,c119C4,c129C4,c139C4;
wire signed [4:0] c109D4,c119D4,c129D4,c139D4;
wire signed [4:0] c10A04,c11A04,c12A04,c13A04;
wire signed [4:0] c10A14,c11A14,c12A14,c13A14;
wire signed [4:0] c10A24,c11A24,c12A24,c13A24;
wire signed [4:0] c10A34,c11A34,c12A34,c13A34;
wire signed [4:0] c10A44,c11A44,c12A44,c13A44;
wire signed [4:0] c10A54,c11A54,c12A54,c13A54;
wire signed [4:0] c10A64,c11A64,c12A64,c13A64;
wire signed [4:0] c10A74,c11A74,c12A74,c13A74;
wire signed [4:0] c10A84,c11A84,c12A84,c13A84;
wire signed [4:0] c10A94,c11A94,c12A94,c13A94;
wire signed [4:0] c10AA4,c11AA4,c12AA4,c13AA4;
wire signed [4:0] c10AB4,c11AB4,c12AB4,c13AB4;
wire signed [4:0] c10AC4,c11AC4,c12AC4,c13AC4;
wire signed [4:0] c10AD4,c11AD4,c12AD4,c13AD4;
wire signed [4:0] c10B04,c11B04,c12B04,c13B04;
wire signed [4:0] c10B14,c11B14,c12B14,c13B14;
wire signed [4:0] c10B24,c11B24,c12B24,c13B24;
wire signed [4:0] c10B34,c11B34,c12B34,c13B34;
wire signed [4:0] c10B44,c11B44,c12B44,c13B44;
wire signed [4:0] c10B54,c11B54,c12B54,c13B54;
wire signed [4:0] c10B64,c11B64,c12B64,c13B64;
wire signed [4:0] c10B74,c11B74,c12B74,c13B74;
wire signed [4:0] c10B84,c11B84,c12B84,c13B84;
wire signed [4:0] c10B94,c11B94,c12B94,c13B94;
wire signed [4:0] c10BA4,c11BA4,c12BA4,c13BA4;
wire signed [4:0] c10BB4,c11BB4,c12BB4,c13BB4;
wire signed [4:0] c10BC4,c11BC4,c12BC4,c13BC4;
wire signed [4:0] c10BD4,c11BD4,c12BD4,c13BD4;
wire signed [4:0] c10C04,c11C04,c12C04,c13C04;
wire signed [4:0] c10C14,c11C14,c12C14,c13C14;
wire signed [4:0] c10C24,c11C24,c12C24,c13C24;
wire signed [4:0] c10C34,c11C34,c12C34,c13C34;
wire signed [4:0] c10C44,c11C44,c12C44,c13C44;
wire signed [4:0] c10C54,c11C54,c12C54,c13C54;
wire signed [4:0] c10C64,c11C64,c12C64,c13C64;
wire signed [4:0] c10C74,c11C74,c12C74,c13C74;
wire signed [4:0] c10C84,c11C84,c12C84,c13C84;
wire signed [4:0] c10C94,c11C94,c12C94,c13C94;
wire signed [4:0] c10CA4,c11CA4,c12CA4,c13CA4;
wire signed [4:0] c10CB4,c11CB4,c12CB4,c13CB4;
wire signed [4:0] c10CC4,c11CC4,c12CC4,c13CC4;
wire signed [4:0] c10CD4,c11CD4,c12CD4,c13CD4;
wire signed [4:0] c10D04,c11D04,c12D04,c13D04;
wire signed [4:0] c10D14,c11D14,c12D14,c13D14;
wire signed [4:0] c10D24,c11D24,c12D24,c13D24;
wire signed [4:0] c10D34,c11D34,c12D34,c13D34;
wire signed [4:0] c10D44,c11D44,c12D44,c13D44;
wire signed [4:0] c10D54,c11D54,c12D54,c13D54;
wire signed [4:0] c10D64,c11D64,c12D64,c13D64;
wire signed [4:0] c10D74,c11D74,c12D74,c13D74;
wire signed [4:0] c10D84,c11D84,c12D84,c13D84;
wire signed [4:0] c10D94,c11D94,c12D94,c13D94;
wire signed [4:0] c10DA4,c11DA4,c12DA4,c13DA4;
wire signed [4:0] c10DB4,c11DB4,c12DB4,c13DB4;
wire signed [4:0] c10DC4,c11DC4,c12DC4,c13DC4;
wire signed [4:0] c10DD4,c11DD4,c12DD4,c13DD4;
wire signed [4:0] c10005,c11005,c12005,c13005;
wire signed [4:0] c10015,c11015,c12015,c13015;
wire signed [4:0] c10025,c11025,c12025,c13025;
wire signed [4:0] c10035,c11035,c12035,c13035;
wire signed [4:0] c10045,c11045,c12045,c13045;
wire signed [4:0] c10055,c11055,c12055,c13055;
wire signed [4:0] c10065,c11065,c12065,c13065;
wire signed [4:0] c10075,c11075,c12075,c13075;
wire signed [4:0] c10085,c11085,c12085,c13085;
wire signed [4:0] c10095,c11095,c12095,c13095;
wire signed [4:0] c100A5,c110A5,c120A5,c130A5;
wire signed [4:0] c100B5,c110B5,c120B5,c130B5;
wire signed [4:0] c100C5,c110C5,c120C5,c130C5;
wire signed [4:0] c100D5,c110D5,c120D5,c130D5;
wire signed [4:0] c10105,c11105,c12105,c13105;
wire signed [4:0] c10115,c11115,c12115,c13115;
wire signed [4:0] c10125,c11125,c12125,c13125;
wire signed [4:0] c10135,c11135,c12135,c13135;
wire signed [4:0] c10145,c11145,c12145,c13145;
wire signed [4:0] c10155,c11155,c12155,c13155;
wire signed [4:0] c10165,c11165,c12165,c13165;
wire signed [4:0] c10175,c11175,c12175,c13175;
wire signed [4:0] c10185,c11185,c12185,c13185;
wire signed [4:0] c10195,c11195,c12195,c13195;
wire signed [4:0] c101A5,c111A5,c121A5,c131A5;
wire signed [4:0] c101B5,c111B5,c121B5,c131B5;
wire signed [4:0] c101C5,c111C5,c121C5,c131C5;
wire signed [4:0] c101D5,c111D5,c121D5,c131D5;
wire signed [4:0] c10205,c11205,c12205,c13205;
wire signed [4:0] c10215,c11215,c12215,c13215;
wire signed [4:0] c10225,c11225,c12225,c13225;
wire signed [4:0] c10235,c11235,c12235,c13235;
wire signed [4:0] c10245,c11245,c12245,c13245;
wire signed [4:0] c10255,c11255,c12255,c13255;
wire signed [4:0] c10265,c11265,c12265,c13265;
wire signed [4:0] c10275,c11275,c12275,c13275;
wire signed [4:0] c10285,c11285,c12285,c13285;
wire signed [4:0] c10295,c11295,c12295,c13295;
wire signed [4:0] c102A5,c112A5,c122A5,c132A5;
wire signed [4:0] c102B5,c112B5,c122B5,c132B5;
wire signed [4:0] c102C5,c112C5,c122C5,c132C5;
wire signed [4:0] c102D5,c112D5,c122D5,c132D5;
wire signed [4:0] c10305,c11305,c12305,c13305;
wire signed [4:0] c10315,c11315,c12315,c13315;
wire signed [4:0] c10325,c11325,c12325,c13325;
wire signed [4:0] c10335,c11335,c12335,c13335;
wire signed [4:0] c10345,c11345,c12345,c13345;
wire signed [4:0] c10355,c11355,c12355,c13355;
wire signed [4:0] c10365,c11365,c12365,c13365;
wire signed [4:0] c10375,c11375,c12375,c13375;
wire signed [4:0] c10385,c11385,c12385,c13385;
wire signed [4:0] c10395,c11395,c12395,c13395;
wire signed [4:0] c103A5,c113A5,c123A5,c133A5;
wire signed [4:0] c103B5,c113B5,c123B5,c133B5;
wire signed [4:0] c103C5,c113C5,c123C5,c133C5;
wire signed [4:0] c103D5,c113D5,c123D5,c133D5;
wire signed [4:0] c10405,c11405,c12405,c13405;
wire signed [4:0] c10415,c11415,c12415,c13415;
wire signed [4:0] c10425,c11425,c12425,c13425;
wire signed [4:0] c10435,c11435,c12435,c13435;
wire signed [4:0] c10445,c11445,c12445,c13445;
wire signed [4:0] c10455,c11455,c12455,c13455;
wire signed [4:0] c10465,c11465,c12465,c13465;
wire signed [4:0] c10475,c11475,c12475,c13475;
wire signed [4:0] c10485,c11485,c12485,c13485;
wire signed [4:0] c10495,c11495,c12495,c13495;
wire signed [4:0] c104A5,c114A5,c124A5,c134A5;
wire signed [4:0] c104B5,c114B5,c124B5,c134B5;
wire signed [4:0] c104C5,c114C5,c124C5,c134C5;
wire signed [4:0] c104D5,c114D5,c124D5,c134D5;
wire signed [4:0] c10505,c11505,c12505,c13505;
wire signed [4:0] c10515,c11515,c12515,c13515;
wire signed [4:0] c10525,c11525,c12525,c13525;
wire signed [4:0] c10535,c11535,c12535,c13535;
wire signed [4:0] c10545,c11545,c12545,c13545;
wire signed [4:0] c10555,c11555,c12555,c13555;
wire signed [4:0] c10565,c11565,c12565,c13565;
wire signed [4:0] c10575,c11575,c12575,c13575;
wire signed [4:0] c10585,c11585,c12585,c13585;
wire signed [4:0] c10595,c11595,c12595,c13595;
wire signed [4:0] c105A5,c115A5,c125A5,c135A5;
wire signed [4:0] c105B5,c115B5,c125B5,c135B5;
wire signed [4:0] c105C5,c115C5,c125C5,c135C5;
wire signed [4:0] c105D5,c115D5,c125D5,c135D5;
wire signed [4:0] c10605,c11605,c12605,c13605;
wire signed [4:0] c10615,c11615,c12615,c13615;
wire signed [4:0] c10625,c11625,c12625,c13625;
wire signed [4:0] c10635,c11635,c12635,c13635;
wire signed [4:0] c10645,c11645,c12645,c13645;
wire signed [4:0] c10655,c11655,c12655,c13655;
wire signed [4:0] c10665,c11665,c12665,c13665;
wire signed [4:0] c10675,c11675,c12675,c13675;
wire signed [4:0] c10685,c11685,c12685,c13685;
wire signed [4:0] c10695,c11695,c12695,c13695;
wire signed [4:0] c106A5,c116A5,c126A5,c136A5;
wire signed [4:0] c106B5,c116B5,c126B5,c136B5;
wire signed [4:0] c106C5,c116C5,c126C5,c136C5;
wire signed [4:0] c106D5,c116D5,c126D5,c136D5;
wire signed [4:0] c10705,c11705,c12705,c13705;
wire signed [4:0] c10715,c11715,c12715,c13715;
wire signed [4:0] c10725,c11725,c12725,c13725;
wire signed [4:0] c10735,c11735,c12735,c13735;
wire signed [4:0] c10745,c11745,c12745,c13745;
wire signed [4:0] c10755,c11755,c12755,c13755;
wire signed [4:0] c10765,c11765,c12765,c13765;
wire signed [4:0] c10775,c11775,c12775,c13775;
wire signed [4:0] c10785,c11785,c12785,c13785;
wire signed [4:0] c10795,c11795,c12795,c13795;
wire signed [4:0] c107A5,c117A5,c127A5,c137A5;
wire signed [4:0] c107B5,c117B5,c127B5,c137B5;
wire signed [4:0] c107C5,c117C5,c127C5,c137C5;
wire signed [4:0] c107D5,c117D5,c127D5,c137D5;
wire signed [4:0] c10805,c11805,c12805,c13805;
wire signed [4:0] c10815,c11815,c12815,c13815;
wire signed [4:0] c10825,c11825,c12825,c13825;
wire signed [4:0] c10835,c11835,c12835,c13835;
wire signed [4:0] c10845,c11845,c12845,c13845;
wire signed [4:0] c10855,c11855,c12855,c13855;
wire signed [4:0] c10865,c11865,c12865,c13865;
wire signed [4:0] c10875,c11875,c12875,c13875;
wire signed [4:0] c10885,c11885,c12885,c13885;
wire signed [4:0] c10895,c11895,c12895,c13895;
wire signed [4:0] c108A5,c118A5,c128A5,c138A5;
wire signed [4:0] c108B5,c118B5,c128B5,c138B5;
wire signed [4:0] c108C5,c118C5,c128C5,c138C5;
wire signed [4:0] c108D5,c118D5,c128D5,c138D5;
wire signed [4:0] c10905,c11905,c12905,c13905;
wire signed [4:0] c10915,c11915,c12915,c13915;
wire signed [4:0] c10925,c11925,c12925,c13925;
wire signed [4:0] c10935,c11935,c12935,c13935;
wire signed [4:0] c10945,c11945,c12945,c13945;
wire signed [4:0] c10955,c11955,c12955,c13955;
wire signed [4:0] c10965,c11965,c12965,c13965;
wire signed [4:0] c10975,c11975,c12975,c13975;
wire signed [4:0] c10985,c11985,c12985,c13985;
wire signed [4:0] c10995,c11995,c12995,c13995;
wire signed [4:0] c109A5,c119A5,c129A5,c139A5;
wire signed [4:0] c109B5,c119B5,c129B5,c139B5;
wire signed [4:0] c109C5,c119C5,c129C5,c139C5;
wire signed [4:0] c109D5,c119D5,c129D5,c139D5;
wire signed [4:0] c10A05,c11A05,c12A05,c13A05;
wire signed [4:0] c10A15,c11A15,c12A15,c13A15;
wire signed [4:0] c10A25,c11A25,c12A25,c13A25;
wire signed [4:0] c10A35,c11A35,c12A35,c13A35;
wire signed [4:0] c10A45,c11A45,c12A45,c13A45;
wire signed [4:0] c10A55,c11A55,c12A55,c13A55;
wire signed [4:0] c10A65,c11A65,c12A65,c13A65;
wire signed [4:0] c10A75,c11A75,c12A75,c13A75;
wire signed [4:0] c10A85,c11A85,c12A85,c13A85;
wire signed [4:0] c10A95,c11A95,c12A95,c13A95;
wire signed [4:0] c10AA5,c11AA5,c12AA5,c13AA5;
wire signed [4:0] c10AB5,c11AB5,c12AB5,c13AB5;
wire signed [4:0] c10AC5,c11AC5,c12AC5,c13AC5;
wire signed [4:0] c10AD5,c11AD5,c12AD5,c13AD5;
wire signed [4:0] c10B05,c11B05,c12B05,c13B05;
wire signed [4:0] c10B15,c11B15,c12B15,c13B15;
wire signed [4:0] c10B25,c11B25,c12B25,c13B25;
wire signed [4:0] c10B35,c11B35,c12B35,c13B35;
wire signed [4:0] c10B45,c11B45,c12B45,c13B45;
wire signed [4:0] c10B55,c11B55,c12B55,c13B55;
wire signed [4:0] c10B65,c11B65,c12B65,c13B65;
wire signed [4:0] c10B75,c11B75,c12B75,c13B75;
wire signed [4:0] c10B85,c11B85,c12B85,c13B85;
wire signed [4:0] c10B95,c11B95,c12B95,c13B95;
wire signed [4:0] c10BA5,c11BA5,c12BA5,c13BA5;
wire signed [4:0] c10BB5,c11BB5,c12BB5,c13BB5;
wire signed [4:0] c10BC5,c11BC5,c12BC5,c13BC5;
wire signed [4:0] c10BD5,c11BD5,c12BD5,c13BD5;
wire signed [4:0] c10C05,c11C05,c12C05,c13C05;
wire signed [4:0] c10C15,c11C15,c12C15,c13C15;
wire signed [4:0] c10C25,c11C25,c12C25,c13C25;
wire signed [4:0] c10C35,c11C35,c12C35,c13C35;
wire signed [4:0] c10C45,c11C45,c12C45,c13C45;
wire signed [4:0] c10C55,c11C55,c12C55,c13C55;
wire signed [4:0] c10C65,c11C65,c12C65,c13C65;
wire signed [4:0] c10C75,c11C75,c12C75,c13C75;
wire signed [4:0] c10C85,c11C85,c12C85,c13C85;
wire signed [4:0] c10C95,c11C95,c12C95,c13C95;
wire signed [4:0] c10CA5,c11CA5,c12CA5,c13CA5;
wire signed [4:0] c10CB5,c11CB5,c12CB5,c13CB5;
wire signed [4:0] c10CC5,c11CC5,c12CC5,c13CC5;
wire signed [4:0] c10CD5,c11CD5,c12CD5,c13CD5;
wire signed [4:0] c10D05,c11D05,c12D05,c13D05;
wire signed [4:0] c10D15,c11D15,c12D15,c13D15;
wire signed [4:0] c10D25,c11D25,c12D25,c13D25;
wire signed [4:0] c10D35,c11D35,c12D35,c13D35;
wire signed [4:0] c10D45,c11D45,c12D45,c13D45;
wire signed [4:0] c10D55,c11D55,c12D55,c13D55;
wire signed [4:0] c10D65,c11D65,c12D65,c13D65;
wire signed [4:0] c10D75,c11D75,c12D75,c13D75;
wire signed [4:0] c10D85,c11D85,c12D85,c13D85;
wire signed [4:0] c10D95,c11D95,c12D95,c13D95;
wire signed [4:0] c10DA5,c11DA5,c12DA5,c13DA5;
wire signed [4:0] c10DB5,c11DB5,c12DB5,c13DB5;
wire signed [4:0] c10DC5,c11DC5,c12DC5,c13DC5;
wire signed [4:0] c10DD5,c11DD5,c12DD5,c13DD5;
wire signed [4:0] c10006,c11006,c12006,c13006;
wire signed [4:0] c10016,c11016,c12016,c13016;
wire signed [4:0] c10026,c11026,c12026,c13026;
wire signed [4:0] c10036,c11036,c12036,c13036;
wire signed [4:0] c10046,c11046,c12046,c13046;
wire signed [4:0] c10056,c11056,c12056,c13056;
wire signed [4:0] c10066,c11066,c12066,c13066;
wire signed [4:0] c10076,c11076,c12076,c13076;
wire signed [4:0] c10086,c11086,c12086,c13086;
wire signed [4:0] c10096,c11096,c12096,c13096;
wire signed [4:0] c100A6,c110A6,c120A6,c130A6;
wire signed [4:0] c100B6,c110B6,c120B6,c130B6;
wire signed [4:0] c100C6,c110C6,c120C6,c130C6;
wire signed [4:0] c100D6,c110D6,c120D6,c130D6;
wire signed [4:0] c10106,c11106,c12106,c13106;
wire signed [4:0] c10116,c11116,c12116,c13116;
wire signed [4:0] c10126,c11126,c12126,c13126;
wire signed [4:0] c10136,c11136,c12136,c13136;
wire signed [4:0] c10146,c11146,c12146,c13146;
wire signed [4:0] c10156,c11156,c12156,c13156;
wire signed [4:0] c10166,c11166,c12166,c13166;
wire signed [4:0] c10176,c11176,c12176,c13176;
wire signed [4:0] c10186,c11186,c12186,c13186;
wire signed [4:0] c10196,c11196,c12196,c13196;
wire signed [4:0] c101A6,c111A6,c121A6,c131A6;
wire signed [4:0] c101B6,c111B6,c121B6,c131B6;
wire signed [4:0] c101C6,c111C6,c121C6,c131C6;
wire signed [4:0] c101D6,c111D6,c121D6,c131D6;
wire signed [4:0] c10206,c11206,c12206,c13206;
wire signed [4:0] c10216,c11216,c12216,c13216;
wire signed [4:0] c10226,c11226,c12226,c13226;
wire signed [4:0] c10236,c11236,c12236,c13236;
wire signed [4:0] c10246,c11246,c12246,c13246;
wire signed [4:0] c10256,c11256,c12256,c13256;
wire signed [4:0] c10266,c11266,c12266,c13266;
wire signed [4:0] c10276,c11276,c12276,c13276;
wire signed [4:0] c10286,c11286,c12286,c13286;
wire signed [4:0] c10296,c11296,c12296,c13296;
wire signed [4:0] c102A6,c112A6,c122A6,c132A6;
wire signed [4:0] c102B6,c112B6,c122B6,c132B6;
wire signed [4:0] c102C6,c112C6,c122C6,c132C6;
wire signed [4:0] c102D6,c112D6,c122D6,c132D6;
wire signed [4:0] c10306,c11306,c12306,c13306;
wire signed [4:0] c10316,c11316,c12316,c13316;
wire signed [4:0] c10326,c11326,c12326,c13326;
wire signed [4:0] c10336,c11336,c12336,c13336;
wire signed [4:0] c10346,c11346,c12346,c13346;
wire signed [4:0] c10356,c11356,c12356,c13356;
wire signed [4:0] c10366,c11366,c12366,c13366;
wire signed [4:0] c10376,c11376,c12376,c13376;
wire signed [4:0] c10386,c11386,c12386,c13386;
wire signed [4:0] c10396,c11396,c12396,c13396;
wire signed [4:0] c103A6,c113A6,c123A6,c133A6;
wire signed [4:0] c103B6,c113B6,c123B6,c133B6;
wire signed [4:0] c103C6,c113C6,c123C6,c133C6;
wire signed [4:0] c103D6,c113D6,c123D6,c133D6;
wire signed [4:0] c10406,c11406,c12406,c13406;
wire signed [4:0] c10416,c11416,c12416,c13416;
wire signed [4:0] c10426,c11426,c12426,c13426;
wire signed [4:0] c10436,c11436,c12436,c13436;
wire signed [4:0] c10446,c11446,c12446,c13446;
wire signed [4:0] c10456,c11456,c12456,c13456;
wire signed [4:0] c10466,c11466,c12466,c13466;
wire signed [4:0] c10476,c11476,c12476,c13476;
wire signed [4:0] c10486,c11486,c12486,c13486;
wire signed [4:0] c10496,c11496,c12496,c13496;
wire signed [4:0] c104A6,c114A6,c124A6,c134A6;
wire signed [4:0] c104B6,c114B6,c124B6,c134B6;
wire signed [4:0] c104C6,c114C6,c124C6,c134C6;
wire signed [4:0] c104D6,c114D6,c124D6,c134D6;
wire signed [4:0] c10506,c11506,c12506,c13506;
wire signed [4:0] c10516,c11516,c12516,c13516;
wire signed [4:0] c10526,c11526,c12526,c13526;
wire signed [4:0] c10536,c11536,c12536,c13536;
wire signed [4:0] c10546,c11546,c12546,c13546;
wire signed [4:0] c10556,c11556,c12556,c13556;
wire signed [4:0] c10566,c11566,c12566,c13566;
wire signed [4:0] c10576,c11576,c12576,c13576;
wire signed [4:0] c10586,c11586,c12586,c13586;
wire signed [4:0] c10596,c11596,c12596,c13596;
wire signed [4:0] c105A6,c115A6,c125A6,c135A6;
wire signed [4:0] c105B6,c115B6,c125B6,c135B6;
wire signed [4:0] c105C6,c115C6,c125C6,c135C6;
wire signed [4:0] c105D6,c115D6,c125D6,c135D6;
wire signed [4:0] c10606,c11606,c12606,c13606;
wire signed [4:0] c10616,c11616,c12616,c13616;
wire signed [4:0] c10626,c11626,c12626,c13626;
wire signed [4:0] c10636,c11636,c12636,c13636;
wire signed [4:0] c10646,c11646,c12646,c13646;
wire signed [4:0] c10656,c11656,c12656,c13656;
wire signed [4:0] c10666,c11666,c12666,c13666;
wire signed [4:0] c10676,c11676,c12676,c13676;
wire signed [4:0] c10686,c11686,c12686,c13686;
wire signed [4:0] c10696,c11696,c12696,c13696;
wire signed [4:0] c106A6,c116A6,c126A6,c136A6;
wire signed [4:0] c106B6,c116B6,c126B6,c136B6;
wire signed [4:0] c106C6,c116C6,c126C6,c136C6;
wire signed [4:0] c106D6,c116D6,c126D6,c136D6;
wire signed [4:0] c10706,c11706,c12706,c13706;
wire signed [4:0] c10716,c11716,c12716,c13716;
wire signed [4:0] c10726,c11726,c12726,c13726;
wire signed [4:0] c10736,c11736,c12736,c13736;
wire signed [4:0] c10746,c11746,c12746,c13746;
wire signed [4:0] c10756,c11756,c12756,c13756;
wire signed [4:0] c10766,c11766,c12766,c13766;
wire signed [4:0] c10776,c11776,c12776,c13776;
wire signed [4:0] c10786,c11786,c12786,c13786;
wire signed [4:0] c10796,c11796,c12796,c13796;
wire signed [4:0] c107A6,c117A6,c127A6,c137A6;
wire signed [4:0] c107B6,c117B6,c127B6,c137B6;
wire signed [4:0] c107C6,c117C6,c127C6,c137C6;
wire signed [4:0] c107D6,c117D6,c127D6,c137D6;
wire signed [4:0] c10806,c11806,c12806,c13806;
wire signed [4:0] c10816,c11816,c12816,c13816;
wire signed [4:0] c10826,c11826,c12826,c13826;
wire signed [4:0] c10836,c11836,c12836,c13836;
wire signed [4:0] c10846,c11846,c12846,c13846;
wire signed [4:0] c10856,c11856,c12856,c13856;
wire signed [4:0] c10866,c11866,c12866,c13866;
wire signed [4:0] c10876,c11876,c12876,c13876;
wire signed [4:0] c10886,c11886,c12886,c13886;
wire signed [4:0] c10896,c11896,c12896,c13896;
wire signed [4:0] c108A6,c118A6,c128A6,c138A6;
wire signed [4:0] c108B6,c118B6,c128B6,c138B6;
wire signed [4:0] c108C6,c118C6,c128C6,c138C6;
wire signed [4:0] c108D6,c118D6,c128D6,c138D6;
wire signed [4:0] c10906,c11906,c12906,c13906;
wire signed [4:0] c10916,c11916,c12916,c13916;
wire signed [4:0] c10926,c11926,c12926,c13926;
wire signed [4:0] c10936,c11936,c12936,c13936;
wire signed [4:0] c10946,c11946,c12946,c13946;
wire signed [4:0] c10956,c11956,c12956,c13956;
wire signed [4:0] c10966,c11966,c12966,c13966;
wire signed [4:0] c10976,c11976,c12976,c13976;
wire signed [4:0] c10986,c11986,c12986,c13986;
wire signed [4:0] c10996,c11996,c12996,c13996;
wire signed [4:0] c109A6,c119A6,c129A6,c139A6;
wire signed [4:0] c109B6,c119B6,c129B6,c139B6;
wire signed [4:0] c109C6,c119C6,c129C6,c139C6;
wire signed [4:0] c109D6,c119D6,c129D6,c139D6;
wire signed [4:0] c10A06,c11A06,c12A06,c13A06;
wire signed [4:0] c10A16,c11A16,c12A16,c13A16;
wire signed [4:0] c10A26,c11A26,c12A26,c13A26;
wire signed [4:0] c10A36,c11A36,c12A36,c13A36;
wire signed [4:0] c10A46,c11A46,c12A46,c13A46;
wire signed [4:0] c10A56,c11A56,c12A56,c13A56;
wire signed [4:0] c10A66,c11A66,c12A66,c13A66;
wire signed [4:0] c10A76,c11A76,c12A76,c13A76;
wire signed [4:0] c10A86,c11A86,c12A86,c13A86;
wire signed [4:0] c10A96,c11A96,c12A96,c13A96;
wire signed [4:0] c10AA6,c11AA6,c12AA6,c13AA6;
wire signed [4:0] c10AB6,c11AB6,c12AB6,c13AB6;
wire signed [4:0] c10AC6,c11AC6,c12AC6,c13AC6;
wire signed [4:0] c10AD6,c11AD6,c12AD6,c13AD6;
wire signed [4:0] c10B06,c11B06,c12B06,c13B06;
wire signed [4:0] c10B16,c11B16,c12B16,c13B16;
wire signed [4:0] c10B26,c11B26,c12B26,c13B26;
wire signed [4:0] c10B36,c11B36,c12B36,c13B36;
wire signed [4:0] c10B46,c11B46,c12B46,c13B46;
wire signed [4:0] c10B56,c11B56,c12B56,c13B56;
wire signed [4:0] c10B66,c11B66,c12B66,c13B66;
wire signed [4:0] c10B76,c11B76,c12B76,c13B76;
wire signed [4:0] c10B86,c11B86,c12B86,c13B86;
wire signed [4:0] c10B96,c11B96,c12B96,c13B96;
wire signed [4:0] c10BA6,c11BA6,c12BA6,c13BA6;
wire signed [4:0] c10BB6,c11BB6,c12BB6,c13BB6;
wire signed [4:0] c10BC6,c11BC6,c12BC6,c13BC6;
wire signed [4:0] c10BD6,c11BD6,c12BD6,c13BD6;
wire signed [4:0] c10C06,c11C06,c12C06,c13C06;
wire signed [4:0] c10C16,c11C16,c12C16,c13C16;
wire signed [4:0] c10C26,c11C26,c12C26,c13C26;
wire signed [4:0] c10C36,c11C36,c12C36,c13C36;
wire signed [4:0] c10C46,c11C46,c12C46,c13C46;
wire signed [4:0] c10C56,c11C56,c12C56,c13C56;
wire signed [4:0] c10C66,c11C66,c12C66,c13C66;
wire signed [4:0] c10C76,c11C76,c12C76,c13C76;
wire signed [4:0] c10C86,c11C86,c12C86,c13C86;
wire signed [4:0] c10C96,c11C96,c12C96,c13C96;
wire signed [4:0] c10CA6,c11CA6,c12CA6,c13CA6;
wire signed [4:0] c10CB6,c11CB6,c12CB6,c13CB6;
wire signed [4:0] c10CC6,c11CC6,c12CC6,c13CC6;
wire signed [4:0] c10CD6,c11CD6,c12CD6,c13CD6;
wire signed [4:0] c10D06,c11D06,c12D06,c13D06;
wire signed [4:0] c10D16,c11D16,c12D16,c13D16;
wire signed [4:0] c10D26,c11D26,c12D26,c13D26;
wire signed [4:0] c10D36,c11D36,c12D36,c13D36;
wire signed [4:0] c10D46,c11D46,c12D46,c13D46;
wire signed [4:0] c10D56,c11D56,c12D56,c13D56;
wire signed [4:0] c10D66,c11D66,c12D66,c13D66;
wire signed [4:0] c10D76,c11D76,c12D76,c13D76;
wire signed [4:0] c10D86,c11D86,c12D86,c13D86;
wire signed [4:0] c10D96,c11D96,c12D96,c13D96;
wire signed [4:0] c10DA6,c11DA6,c12DA6,c13DA6;
wire signed [4:0] c10DB6,c11DB6,c12DB6,c13DB6;
wire signed [4:0] c10DC6,c11DC6,c12DC6,c13DC6;
wire signed [4:0] c10DD6,c11DD6,c12DD6,c13DD6;
wire signed [4:0] c10007,c11007,c12007,c13007;
wire signed [4:0] c10017,c11017,c12017,c13017;
wire signed [4:0] c10027,c11027,c12027,c13027;
wire signed [4:0] c10037,c11037,c12037,c13037;
wire signed [4:0] c10047,c11047,c12047,c13047;
wire signed [4:0] c10057,c11057,c12057,c13057;
wire signed [4:0] c10067,c11067,c12067,c13067;
wire signed [4:0] c10077,c11077,c12077,c13077;
wire signed [4:0] c10087,c11087,c12087,c13087;
wire signed [4:0] c10097,c11097,c12097,c13097;
wire signed [4:0] c100A7,c110A7,c120A7,c130A7;
wire signed [4:0] c100B7,c110B7,c120B7,c130B7;
wire signed [4:0] c100C7,c110C7,c120C7,c130C7;
wire signed [4:0] c100D7,c110D7,c120D7,c130D7;
wire signed [4:0] c10107,c11107,c12107,c13107;
wire signed [4:0] c10117,c11117,c12117,c13117;
wire signed [4:0] c10127,c11127,c12127,c13127;
wire signed [4:0] c10137,c11137,c12137,c13137;
wire signed [4:0] c10147,c11147,c12147,c13147;
wire signed [4:0] c10157,c11157,c12157,c13157;
wire signed [4:0] c10167,c11167,c12167,c13167;
wire signed [4:0] c10177,c11177,c12177,c13177;
wire signed [4:0] c10187,c11187,c12187,c13187;
wire signed [4:0] c10197,c11197,c12197,c13197;
wire signed [4:0] c101A7,c111A7,c121A7,c131A7;
wire signed [4:0] c101B7,c111B7,c121B7,c131B7;
wire signed [4:0] c101C7,c111C7,c121C7,c131C7;
wire signed [4:0] c101D7,c111D7,c121D7,c131D7;
wire signed [4:0] c10207,c11207,c12207,c13207;
wire signed [4:0] c10217,c11217,c12217,c13217;
wire signed [4:0] c10227,c11227,c12227,c13227;
wire signed [4:0] c10237,c11237,c12237,c13237;
wire signed [4:0] c10247,c11247,c12247,c13247;
wire signed [4:0] c10257,c11257,c12257,c13257;
wire signed [4:0] c10267,c11267,c12267,c13267;
wire signed [4:0] c10277,c11277,c12277,c13277;
wire signed [4:0] c10287,c11287,c12287,c13287;
wire signed [4:0] c10297,c11297,c12297,c13297;
wire signed [4:0] c102A7,c112A7,c122A7,c132A7;
wire signed [4:0] c102B7,c112B7,c122B7,c132B7;
wire signed [4:0] c102C7,c112C7,c122C7,c132C7;
wire signed [4:0] c102D7,c112D7,c122D7,c132D7;
wire signed [4:0] c10307,c11307,c12307,c13307;
wire signed [4:0] c10317,c11317,c12317,c13317;
wire signed [4:0] c10327,c11327,c12327,c13327;
wire signed [4:0] c10337,c11337,c12337,c13337;
wire signed [4:0] c10347,c11347,c12347,c13347;
wire signed [4:0] c10357,c11357,c12357,c13357;
wire signed [4:0] c10367,c11367,c12367,c13367;
wire signed [4:0] c10377,c11377,c12377,c13377;
wire signed [4:0] c10387,c11387,c12387,c13387;
wire signed [4:0] c10397,c11397,c12397,c13397;
wire signed [4:0] c103A7,c113A7,c123A7,c133A7;
wire signed [4:0] c103B7,c113B7,c123B7,c133B7;
wire signed [4:0] c103C7,c113C7,c123C7,c133C7;
wire signed [4:0] c103D7,c113D7,c123D7,c133D7;
wire signed [4:0] c10407,c11407,c12407,c13407;
wire signed [4:0] c10417,c11417,c12417,c13417;
wire signed [4:0] c10427,c11427,c12427,c13427;
wire signed [4:0] c10437,c11437,c12437,c13437;
wire signed [4:0] c10447,c11447,c12447,c13447;
wire signed [4:0] c10457,c11457,c12457,c13457;
wire signed [4:0] c10467,c11467,c12467,c13467;
wire signed [4:0] c10477,c11477,c12477,c13477;
wire signed [4:0] c10487,c11487,c12487,c13487;
wire signed [4:0] c10497,c11497,c12497,c13497;
wire signed [4:0] c104A7,c114A7,c124A7,c134A7;
wire signed [4:0] c104B7,c114B7,c124B7,c134B7;
wire signed [4:0] c104C7,c114C7,c124C7,c134C7;
wire signed [4:0] c104D7,c114D7,c124D7,c134D7;
wire signed [4:0] c10507,c11507,c12507,c13507;
wire signed [4:0] c10517,c11517,c12517,c13517;
wire signed [4:0] c10527,c11527,c12527,c13527;
wire signed [4:0] c10537,c11537,c12537,c13537;
wire signed [4:0] c10547,c11547,c12547,c13547;
wire signed [4:0] c10557,c11557,c12557,c13557;
wire signed [4:0] c10567,c11567,c12567,c13567;
wire signed [4:0] c10577,c11577,c12577,c13577;
wire signed [4:0] c10587,c11587,c12587,c13587;
wire signed [4:0] c10597,c11597,c12597,c13597;
wire signed [4:0] c105A7,c115A7,c125A7,c135A7;
wire signed [4:0] c105B7,c115B7,c125B7,c135B7;
wire signed [4:0] c105C7,c115C7,c125C7,c135C7;
wire signed [4:0] c105D7,c115D7,c125D7,c135D7;
wire signed [4:0] c10607,c11607,c12607,c13607;
wire signed [4:0] c10617,c11617,c12617,c13617;
wire signed [4:0] c10627,c11627,c12627,c13627;
wire signed [4:0] c10637,c11637,c12637,c13637;
wire signed [4:0] c10647,c11647,c12647,c13647;
wire signed [4:0] c10657,c11657,c12657,c13657;
wire signed [4:0] c10667,c11667,c12667,c13667;
wire signed [4:0] c10677,c11677,c12677,c13677;
wire signed [4:0] c10687,c11687,c12687,c13687;
wire signed [4:0] c10697,c11697,c12697,c13697;
wire signed [4:0] c106A7,c116A7,c126A7,c136A7;
wire signed [4:0] c106B7,c116B7,c126B7,c136B7;
wire signed [4:0] c106C7,c116C7,c126C7,c136C7;
wire signed [4:0] c106D7,c116D7,c126D7,c136D7;
wire signed [4:0] c10707,c11707,c12707,c13707;
wire signed [4:0] c10717,c11717,c12717,c13717;
wire signed [4:0] c10727,c11727,c12727,c13727;
wire signed [4:0] c10737,c11737,c12737,c13737;
wire signed [4:0] c10747,c11747,c12747,c13747;
wire signed [4:0] c10757,c11757,c12757,c13757;
wire signed [4:0] c10767,c11767,c12767,c13767;
wire signed [4:0] c10777,c11777,c12777,c13777;
wire signed [4:0] c10787,c11787,c12787,c13787;
wire signed [4:0] c10797,c11797,c12797,c13797;
wire signed [4:0] c107A7,c117A7,c127A7,c137A7;
wire signed [4:0] c107B7,c117B7,c127B7,c137B7;
wire signed [4:0] c107C7,c117C7,c127C7,c137C7;
wire signed [4:0] c107D7,c117D7,c127D7,c137D7;
wire signed [4:0] c10807,c11807,c12807,c13807;
wire signed [4:0] c10817,c11817,c12817,c13817;
wire signed [4:0] c10827,c11827,c12827,c13827;
wire signed [4:0] c10837,c11837,c12837,c13837;
wire signed [4:0] c10847,c11847,c12847,c13847;
wire signed [4:0] c10857,c11857,c12857,c13857;
wire signed [4:0] c10867,c11867,c12867,c13867;
wire signed [4:0] c10877,c11877,c12877,c13877;
wire signed [4:0] c10887,c11887,c12887,c13887;
wire signed [4:0] c10897,c11897,c12897,c13897;
wire signed [4:0] c108A7,c118A7,c128A7,c138A7;
wire signed [4:0] c108B7,c118B7,c128B7,c138B7;
wire signed [4:0] c108C7,c118C7,c128C7,c138C7;
wire signed [4:0] c108D7,c118D7,c128D7,c138D7;
wire signed [4:0] c10907,c11907,c12907,c13907;
wire signed [4:0] c10917,c11917,c12917,c13917;
wire signed [4:0] c10927,c11927,c12927,c13927;
wire signed [4:0] c10937,c11937,c12937,c13937;
wire signed [4:0] c10947,c11947,c12947,c13947;
wire signed [4:0] c10957,c11957,c12957,c13957;
wire signed [4:0] c10967,c11967,c12967,c13967;
wire signed [4:0] c10977,c11977,c12977,c13977;
wire signed [4:0] c10987,c11987,c12987,c13987;
wire signed [4:0] c10997,c11997,c12997,c13997;
wire signed [4:0] c109A7,c119A7,c129A7,c139A7;
wire signed [4:0] c109B7,c119B7,c129B7,c139B7;
wire signed [4:0] c109C7,c119C7,c129C7,c139C7;
wire signed [4:0] c109D7,c119D7,c129D7,c139D7;
wire signed [4:0] c10A07,c11A07,c12A07,c13A07;
wire signed [4:0] c10A17,c11A17,c12A17,c13A17;
wire signed [4:0] c10A27,c11A27,c12A27,c13A27;
wire signed [4:0] c10A37,c11A37,c12A37,c13A37;
wire signed [4:0] c10A47,c11A47,c12A47,c13A47;
wire signed [4:0] c10A57,c11A57,c12A57,c13A57;
wire signed [4:0] c10A67,c11A67,c12A67,c13A67;
wire signed [4:0] c10A77,c11A77,c12A77,c13A77;
wire signed [4:0] c10A87,c11A87,c12A87,c13A87;
wire signed [4:0] c10A97,c11A97,c12A97,c13A97;
wire signed [4:0] c10AA7,c11AA7,c12AA7,c13AA7;
wire signed [4:0] c10AB7,c11AB7,c12AB7,c13AB7;
wire signed [4:0] c10AC7,c11AC7,c12AC7,c13AC7;
wire signed [4:0] c10AD7,c11AD7,c12AD7,c13AD7;
wire signed [4:0] c10B07,c11B07,c12B07,c13B07;
wire signed [4:0] c10B17,c11B17,c12B17,c13B17;
wire signed [4:0] c10B27,c11B27,c12B27,c13B27;
wire signed [4:0] c10B37,c11B37,c12B37,c13B37;
wire signed [4:0] c10B47,c11B47,c12B47,c13B47;
wire signed [4:0] c10B57,c11B57,c12B57,c13B57;
wire signed [4:0] c10B67,c11B67,c12B67,c13B67;
wire signed [4:0] c10B77,c11B77,c12B77,c13B77;
wire signed [4:0] c10B87,c11B87,c12B87,c13B87;
wire signed [4:0] c10B97,c11B97,c12B97,c13B97;
wire signed [4:0] c10BA7,c11BA7,c12BA7,c13BA7;
wire signed [4:0] c10BB7,c11BB7,c12BB7,c13BB7;
wire signed [4:0] c10BC7,c11BC7,c12BC7,c13BC7;
wire signed [4:0] c10BD7,c11BD7,c12BD7,c13BD7;
wire signed [4:0] c10C07,c11C07,c12C07,c13C07;
wire signed [4:0] c10C17,c11C17,c12C17,c13C17;
wire signed [4:0] c10C27,c11C27,c12C27,c13C27;
wire signed [4:0] c10C37,c11C37,c12C37,c13C37;
wire signed [4:0] c10C47,c11C47,c12C47,c13C47;
wire signed [4:0] c10C57,c11C57,c12C57,c13C57;
wire signed [4:0] c10C67,c11C67,c12C67,c13C67;
wire signed [4:0] c10C77,c11C77,c12C77,c13C77;
wire signed [4:0] c10C87,c11C87,c12C87,c13C87;
wire signed [4:0] c10C97,c11C97,c12C97,c13C97;
wire signed [4:0] c10CA7,c11CA7,c12CA7,c13CA7;
wire signed [4:0] c10CB7,c11CB7,c12CB7,c13CB7;
wire signed [4:0] c10CC7,c11CC7,c12CC7,c13CC7;
wire signed [4:0] c10CD7,c11CD7,c12CD7,c13CD7;
wire signed [4:0] c10D07,c11D07,c12D07,c13D07;
wire signed [4:0] c10D17,c11D17,c12D17,c13D17;
wire signed [4:0] c10D27,c11D27,c12D27,c13D27;
wire signed [4:0] c10D37,c11D37,c12D37,c13D37;
wire signed [4:0] c10D47,c11D47,c12D47,c13D47;
wire signed [4:0] c10D57,c11D57,c12D57,c13D57;
wire signed [4:0] c10D67,c11D67,c12D67,c13D67;
wire signed [4:0] c10D77,c11D77,c12D77,c13D77;
wire signed [4:0] c10D87,c11D87,c12D87,c13D87;
wire signed [4:0] c10D97,c11D97,c12D97,c13D97;
wire signed [4:0] c10DA7,c11DA7,c12DA7,c13DA7;
wire signed [4:0] c10DB7,c11DB7,c12DB7,c13DB7;
wire signed [4:0] c10DC7,c11DC7,c12DC7,c13DC7;
wire signed [4:0] c10DD7,c11DD7,c12DD7,c13DD7;
wire signed [6:0] C1000;
wire A1000;
wire signed [6:0] C1010;
wire A1010;
wire signed [6:0] C1020;
wire A1020;
wire signed [6:0] C1030;
wire A1030;
wire signed [6:0] C1040;
wire A1040;
wire signed [6:0] C1050;
wire A1050;
wire signed [6:0] C1060;
wire A1060;
wire signed [6:0] C1070;
wire A1070;
wire signed [6:0] C1080;
wire A1080;
wire signed [6:0] C1090;
wire A1090;
wire signed [6:0] C10A0;
wire A10A0;
wire signed [6:0] C10B0;
wire A10B0;
wire signed [6:0] C10C0;
wire A10C0;
wire signed [6:0] C10D0;
wire A10D0;
wire signed [6:0] C1100;
wire A1100;
wire signed [6:0] C1110;
wire A1110;
wire signed [6:0] C1120;
wire A1120;
wire signed [6:0] C1130;
wire A1130;
wire signed [6:0] C1140;
wire A1140;
wire signed [6:0] C1150;
wire A1150;
wire signed [6:0] C1160;
wire A1160;
wire signed [6:0] C1170;
wire A1170;
wire signed [6:0] C1180;
wire A1180;
wire signed [6:0] C1190;
wire A1190;
wire signed [6:0] C11A0;
wire A11A0;
wire signed [6:0] C11B0;
wire A11B0;
wire signed [6:0] C11C0;
wire A11C0;
wire signed [6:0] C11D0;
wire A11D0;
wire signed [6:0] C1200;
wire A1200;
wire signed [6:0] C1210;
wire A1210;
wire signed [6:0] C1220;
wire A1220;
wire signed [6:0] C1230;
wire A1230;
wire signed [6:0] C1240;
wire A1240;
wire signed [6:0] C1250;
wire A1250;
wire signed [6:0] C1260;
wire A1260;
wire signed [6:0] C1270;
wire A1270;
wire signed [6:0] C1280;
wire A1280;
wire signed [6:0] C1290;
wire A1290;
wire signed [6:0] C12A0;
wire A12A0;
wire signed [6:0] C12B0;
wire A12B0;
wire signed [6:0] C12C0;
wire A12C0;
wire signed [6:0] C12D0;
wire A12D0;
wire signed [6:0] C1300;
wire A1300;
wire signed [6:0] C1310;
wire A1310;
wire signed [6:0] C1320;
wire A1320;
wire signed [6:0] C1330;
wire A1330;
wire signed [6:0] C1340;
wire A1340;
wire signed [6:0] C1350;
wire A1350;
wire signed [6:0] C1360;
wire A1360;
wire signed [6:0] C1370;
wire A1370;
wire signed [6:0] C1380;
wire A1380;
wire signed [6:0] C1390;
wire A1390;
wire signed [6:0] C13A0;
wire A13A0;
wire signed [6:0] C13B0;
wire A13B0;
wire signed [6:0] C13C0;
wire A13C0;
wire signed [6:0] C13D0;
wire A13D0;
wire signed [6:0] C1400;
wire A1400;
wire signed [6:0] C1410;
wire A1410;
wire signed [6:0] C1420;
wire A1420;
wire signed [6:0] C1430;
wire A1430;
wire signed [6:0] C1440;
wire A1440;
wire signed [6:0] C1450;
wire A1450;
wire signed [6:0] C1460;
wire A1460;
wire signed [6:0] C1470;
wire A1470;
wire signed [6:0] C1480;
wire A1480;
wire signed [6:0] C1490;
wire A1490;
wire signed [6:0] C14A0;
wire A14A0;
wire signed [6:0] C14B0;
wire A14B0;
wire signed [6:0] C14C0;
wire A14C0;
wire signed [6:0] C14D0;
wire A14D0;
wire signed [6:0] C1500;
wire A1500;
wire signed [6:0] C1510;
wire A1510;
wire signed [6:0] C1520;
wire A1520;
wire signed [6:0] C1530;
wire A1530;
wire signed [6:0] C1540;
wire A1540;
wire signed [6:0] C1550;
wire A1550;
wire signed [6:0] C1560;
wire A1560;
wire signed [6:0] C1570;
wire A1570;
wire signed [6:0] C1580;
wire A1580;
wire signed [6:0] C1590;
wire A1590;
wire signed [6:0] C15A0;
wire A15A0;
wire signed [6:0] C15B0;
wire A15B0;
wire signed [6:0] C15C0;
wire A15C0;
wire signed [6:0] C15D0;
wire A15D0;
wire signed [6:0] C1600;
wire A1600;
wire signed [6:0] C1610;
wire A1610;
wire signed [6:0] C1620;
wire A1620;
wire signed [6:0] C1630;
wire A1630;
wire signed [6:0] C1640;
wire A1640;
wire signed [6:0] C1650;
wire A1650;
wire signed [6:0] C1660;
wire A1660;
wire signed [6:0] C1670;
wire A1670;
wire signed [6:0] C1680;
wire A1680;
wire signed [6:0] C1690;
wire A1690;
wire signed [6:0] C16A0;
wire A16A0;
wire signed [6:0] C16B0;
wire A16B0;
wire signed [6:0] C16C0;
wire A16C0;
wire signed [6:0] C16D0;
wire A16D0;
wire signed [6:0] C1700;
wire A1700;
wire signed [6:0] C1710;
wire A1710;
wire signed [6:0] C1720;
wire A1720;
wire signed [6:0] C1730;
wire A1730;
wire signed [6:0] C1740;
wire A1740;
wire signed [6:0] C1750;
wire A1750;
wire signed [6:0] C1760;
wire A1760;
wire signed [6:0] C1770;
wire A1770;
wire signed [6:0] C1780;
wire A1780;
wire signed [6:0] C1790;
wire A1790;
wire signed [6:0] C17A0;
wire A17A0;
wire signed [6:0] C17B0;
wire A17B0;
wire signed [6:0] C17C0;
wire A17C0;
wire signed [6:0] C17D0;
wire A17D0;
wire signed [6:0] C1800;
wire A1800;
wire signed [6:0] C1810;
wire A1810;
wire signed [6:0] C1820;
wire A1820;
wire signed [6:0] C1830;
wire A1830;
wire signed [6:0] C1840;
wire A1840;
wire signed [6:0] C1850;
wire A1850;
wire signed [6:0] C1860;
wire A1860;
wire signed [6:0] C1870;
wire A1870;
wire signed [6:0] C1880;
wire A1880;
wire signed [6:0] C1890;
wire A1890;
wire signed [6:0] C18A0;
wire A18A0;
wire signed [6:0] C18B0;
wire A18B0;
wire signed [6:0] C18C0;
wire A18C0;
wire signed [6:0] C18D0;
wire A18D0;
wire signed [6:0] C1900;
wire A1900;
wire signed [6:0] C1910;
wire A1910;
wire signed [6:0] C1920;
wire A1920;
wire signed [6:0] C1930;
wire A1930;
wire signed [6:0] C1940;
wire A1940;
wire signed [6:0] C1950;
wire A1950;
wire signed [6:0] C1960;
wire A1960;
wire signed [6:0] C1970;
wire A1970;
wire signed [6:0] C1980;
wire A1980;
wire signed [6:0] C1990;
wire A1990;
wire signed [6:0] C19A0;
wire A19A0;
wire signed [6:0] C19B0;
wire A19B0;
wire signed [6:0] C19C0;
wire A19C0;
wire signed [6:0] C19D0;
wire A19D0;
wire signed [6:0] C1A00;
wire A1A00;
wire signed [6:0] C1A10;
wire A1A10;
wire signed [6:0] C1A20;
wire A1A20;
wire signed [6:0] C1A30;
wire A1A30;
wire signed [6:0] C1A40;
wire A1A40;
wire signed [6:0] C1A50;
wire A1A50;
wire signed [6:0] C1A60;
wire A1A60;
wire signed [6:0] C1A70;
wire A1A70;
wire signed [6:0] C1A80;
wire A1A80;
wire signed [6:0] C1A90;
wire A1A90;
wire signed [6:0] C1AA0;
wire A1AA0;
wire signed [6:0] C1AB0;
wire A1AB0;
wire signed [6:0] C1AC0;
wire A1AC0;
wire signed [6:0] C1AD0;
wire A1AD0;
wire signed [6:0] C1B00;
wire A1B00;
wire signed [6:0] C1B10;
wire A1B10;
wire signed [6:0] C1B20;
wire A1B20;
wire signed [6:0] C1B30;
wire A1B30;
wire signed [6:0] C1B40;
wire A1B40;
wire signed [6:0] C1B50;
wire A1B50;
wire signed [6:0] C1B60;
wire A1B60;
wire signed [6:0] C1B70;
wire A1B70;
wire signed [6:0] C1B80;
wire A1B80;
wire signed [6:0] C1B90;
wire A1B90;
wire signed [6:0] C1BA0;
wire A1BA0;
wire signed [6:0] C1BB0;
wire A1BB0;
wire signed [6:0] C1BC0;
wire A1BC0;
wire signed [6:0] C1BD0;
wire A1BD0;
wire signed [6:0] C1C00;
wire A1C00;
wire signed [6:0] C1C10;
wire A1C10;
wire signed [6:0] C1C20;
wire A1C20;
wire signed [6:0] C1C30;
wire A1C30;
wire signed [6:0] C1C40;
wire A1C40;
wire signed [6:0] C1C50;
wire A1C50;
wire signed [6:0] C1C60;
wire A1C60;
wire signed [6:0] C1C70;
wire A1C70;
wire signed [6:0] C1C80;
wire A1C80;
wire signed [6:0] C1C90;
wire A1C90;
wire signed [6:0] C1CA0;
wire A1CA0;
wire signed [6:0] C1CB0;
wire A1CB0;
wire signed [6:0] C1CC0;
wire A1CC0;
wire signed [6:0] C1CD0;
wire A1CD0;
wire signed [6:0] C1D00;
wire A1D00;
wire signed [6:0] C1D10;
wire A1D10;
wire signed [6:0] C1D20;
wire A1D20;
wire signed [6:0] C1D30;
wire A1D30;
wire signed [6:0] C1D40;
wire A1D40;
wire signed [6:0] C1D50;
wire A1D50;
wire signed [6:0] C1D60;
wire A1D60;
wire signed [6:0] C1D70;
wire A1D70;
wire signed [6:0] C1D80;
wire A1D80;
wire signed [6:0] C1D90;
wire A1D90;
wire signed [6:0] C1DA0;
wire A1DA0;
wire signed [6:0] C1DB0;
wire A1DB0;
wire signed [6:0] C1DC0;
wire A1DC0;
wire signed [6:0] C1DD0;
wire A1DD0;
wire signed [6:0] C1001;
wire A1001;
wire signed [6:0] C1011;
wire A1011;
wire signed [6:0] C1021;
wire A1021;
wire signed [6:0] C1031;
wire A1031;
wire signed [6:0] C1041;
wire A1041;
wire signed [6:0] C1051;
wire A1051;
wire signed [6:0] C1061;
wire A1061;
wire signed [6:0] C1071;
wire A1071;
wire signed [6:0] C1081;
wire A1081;
wire signed [6:0] C1091;
wire A1091;
wire signed [6:0] C10A1;
wire A10A1;
wire signed [6:0] C10B1;
wire A10B1;
wire signed [6:0] C10C1;
wire A10C1;
wire signed [6:0] C10D1;
wire A10D1;
wire signed [6:0] C1101;
wire A1101;
wire signed [6:0] C1111;
wire A1111;
wire signed [6:0] C1121;
wire A1121;
wire signed [6:0] C1131;
wire A1131;
wire signed [6:0] C1141;
wire A1141;
wire signed [6:0] C1151;
wire A1151;
wire signed [6:0] C1161;
wire A1161;
wire signed [6:0] C1171;
wire A1171;
wire signed [6:0] C1181;
wire A1181;
wire signed [6:0] C1191;
wire A1191;
wire signed [6:0] C11A1;
wire A11A1;
wire signed [6:0] C11B1;
wire A11B1;
wire signed [6:0] C11C1;
wire A11C1;
wire signed [6:0] C11D1;
wire A11D1;
wire signed [6:0] C1201;
wire A1201;
wire signed [6:0] C1211;
wire A1211;
wire signed [6:0] C1221;
wire A1221;
wire signed [6:0] C1231;
wire A1231;
wire signed [6:0] C1241;
wire A1241;
wire signed [6:0] C1251;
wire A1251;
wire signed [6:0] C1261;
wire A1261;
wire signed [6:0] C1271;
wire A1271;
wire signed [6:0] C1281;
wire A1281;
wire signed [6:0] C1291;
wire A1291;
wire signed [6:0] C12A1;
wire A12A1;
wire signed [6:0] C12B1;
wire A12B1;
wire signed [6:0] C12C1;
wire A12C1;
wire signed [6:0] C12D1;
wire A12D1;
wire signed [6:0] C1301;
wire A1301;
wire signed [6:0] C1311;
wire A1311;
wire signed [6:0] C1321;
wire A1321;
wire signed [6:0] C1331;
wire A1331;
wire signed [6:0] C1341;
wire A1341;
wire signed [6:0] C1351;
wire A1351;
wire signed [6:0] C1361;
wire A1361;
wire signed [6:0] C1371;
wire A1371;
wire signed [6:0] C1381;
wire A1381;
wire signed [6:0] C1391;
wire A1391;
wire signed [6:0] C13A1;
wire A13A1;
wire signed [6:0] C13B1;
wire A13B1;
wire signed [6:0] C13C1;
wire A13C1;
wire signed [6:0] C13D1;
wire A13D1;
wire signed [6:0] C1401;
wire A1401;
wire signed [6:0] C1411;
wire A1411;
wire signed [6:0] C1421;
wire A1421;
wire signed [6:0] C1431;
wire A1431;
wire signed [6:0] C1441;
wire A1441;
wire signed [6:0] C1451;
wire A1451;
wire signed [6:0] C1461;
wire A1461;
wire signed [6:0] C1471;
wire A1471;
wire signed [6:0] C1481;
wire A1481;
wire signed [6:0] C1491;
wire A1491;
wire signed [6:0] C14A1;
wire A14A1;
wire signed [6:0] C14B1;
wire A14B1;
wire signed [6:0] C14C1;
wire A14C1;
wire signed [6:0] C14D1;
wire A14D1;
wire signed [6:0] C1501;
wire A1501;
wire signed [6:0] C1511;
wire A1511;
wire signed [6:0] C1521;
wire A1521;
wire signed [6:0] C1531;
wire A1531;
wire signed [6:0] C1541;
wire A1541;
wire signed [6:0] C1551;
wire A1551;
wire signed [6:0] C1561;
wire A1561;
wire signed [6:0] C1571;
wire A1571;
wire signed [6:0] C1581;
wire A1581;
wire signed [6:0] C1591;
wire A1591;
wire signed [6:0] C15A1;
wire A15A1;
wire signed [6:0] C15B1;
wire A15B1;
wire signed [6:0] C15C1;
wire A15C1;
wire signed [6:0] C15D1;
wire A15D1;
wire signed [6:0] C1601;
wire A1601;
wire signed [6:0] C1611;
wire A1611;
wire signed [6:0] C1621;
wire A1621;
wire signed [6:0] C1631;
wire A1631;
wire signed [6:0] C1641;
wire A1641;
wire signed [6:0] C1651;
wire A1651;
wire signed [6:0] C1661;
wire A1661;
wire signed [6:0] C1671;
wire A1671;
wire signed [6:0] C1681;
wire A1681;
wire signed [6:0] C1691;
wire A1691;
wire signed [6:0] C16A1;
wire A16A1;
wire signed [6:0] C16B1;
wire A16B1;
wire signed [6:0] C16C1;
wire A16C1;
wire signed [6:0] C16D1;
wire A16D1;
wire signed [6:0] C1701;
wire A1701;
wire signed [6:0] C1711;
wire A1711;
wire signed [6:0] C1721;
wire A1721;
wire signed [6:0] C1731;
wire A1731;
wire signed [6:0] C1741;
wire A1741;
wire signed [6:0] C1751;
wire A1751;
wire signed [6:0] C1761;
wire A1761;
wire signed [6:0] C1771;
wire A1771;
wire signed [6:0] C1781;
wire A1781;
wire signed [6:0] C1791;
wire A1791;
wire signed [6:0] C17A1;
wire A17A1;
wire signed [6:0] C17B1;
wire A17B1;
wire signed [6:0] C17C1;
wire A17C1;
wire signed [6:0] C17D1;
wire A17D1;
wire signed [6:0] C1801;
wire A1801;
wire signed [6:0] C1811;
wire A1811;
wire signed [6:0] C1821;
wire A1821;
wire signed [6:0] C1831;
wire A1831;
wire signed [6:0] C1841;
wire A1841;
wire signed [6:0] C1851;
wire A1851;
wire signed [6:0] C1861;
wire A1861;
wire signed [6:0] C1871;
wire A1871;
wire signed [6:0] C1881;
wire A1881;
wire signed [6:0] C1891;
wire A1891;
wire signed [6:0] C18A1;
wire A18A1;
wire signed [6:0] C18B1;
wire A18B1;
wire signed [6:0] C18C1;
wire A18C1;
wire signed [6:0] C18D1;
wire A18D1;
wire signed [6:0] C1901;
wire A1901;
wire signed [6:0] C1911;
wire A1911;
wire signed [6:0] C1921;
wire A1921;
wire signed [6:0] C1931;
wire A1931;
wire signed [6:0] C1941;
wire A1941;
wire signed [6:0] C1951;
wire A1951;
wire signed [6:0] C1961;
wire A1961;
wire signed [6:0] C1971;
wire A1971;
wire signed [6:0] C1981;
wire A1981;
wire signed [6:0] C1991;
wire A1991;
wire signed [6:0] C19A1;
wire A19A1;
wire signed [6:0] C19B1;
wire A19B1;
wire signed [6:0] C19C1;
wire A19C1;
wire signed [6:0] C19D1;
wire A19D1;
wire signed [6:0] C1A01;
wire A1A01;
wire signed [6:0] C1A11;
wire A1A11;
wire signed [6:0] C1A21;
wire A1A21;
wire signed [6:0] C1A31;
wire A1A31;
wire signed [6:0] C1A41;
wire A1A41;
wire signed [6:0] C1A51;
wire A1A51;
wire signed [6:0] C1A61;
wire A1A61;
wire signed [6:0] C1A71;
wire A1A71;
wire signed [6:0] C1A81;
wire A1A81;
wire signed [6:0] C1A91;
wire A1A91;
wire signed [6:0] C1AA1;
wire A1AA1;
wire signed [6:0] C1AB1;
wire A1AB1;
wire signed [6:0] C1AC1;
wire A1AC1;
wire signed [6:0] C1AD1;
wire A1AD1;
wire signed [6:0] C1B01;
wire A1B01;
wire signed [6:0] C1B11;
wire A1B11;
wire signed [6:0] C1B21;
wire A1B21;
wire signed [6:0] C1B31;
wire A1B31;
wire signed [6:0] C1B41;
wire A1B41;
wire signed [6:0] C1B51;
wire A1B51;
wire signed [6:0] C1B61;
wire A1B61;
wire signed [6:0] C1B71;
wire A1B71;
wire signed [6:0] C1B81;
wire A1B81;
wire signed [6:0] C1B91;
wire A1B91;
wire signed [6:0] C1BA1;
wire A1BA1;
wire signed [6:0] C1BB1;
wire A1BB1;
wire signed [6:0] C1BC1;
wire A1BC1;
wire signed [6:0] C1BD1;
wire A1BD1;
wire signed [6:0] C1C01;
wire A1C01;
wire signed [6:0] C1C11;
wire A1C11;
wire signed [6:0] C1C21;
wire A1C21;
wire signed [6:0] C1C31;
wire A1C31;
wire signed [6:0] C1C41;
wire A1C41;
wire signed [6:0] C1C51;
wire A1C51;
wire signed [6:0] C1C61;
wire A1C61;
wire signed [6:0] C1C71;
wire A1C71;
wire signed [6:0] C1C81;
wire A1C81;
wire signed [6:0] C1C91;
wire A1C91;
wire signed [6:0] C1CA1;
wire A1CA1;
wire signed [6:0] C1CB1;
wire A1CB1;
wire signed [6:0] C1CC1;
wire A1CC1;
wire signed [6:0] C1CD1;
wire A1CD1;
wire signed [6:0] C1D01;
wire A1D01;
wire signed [6:0] C1D11;
wire A1D11;
wire signed [6:0] C1D21;
wire A1D21;
wire signed [6:0] C1D31;
wire A1D31;
wire signed [6:0] C1D41;
wire A1D41;
wire signed [6:0] C1D51;
wire A1D51;
wire signed [6:0] C1D61;
wire A1D61;
wire signed [6:0] C1D71;
wire A1D71;
wire signed [6:0] C1D81;
wire A1D81;
wire signed [6:0] C1D91;
wire A1D91;
wire signed [6:0] C1DA1;
wire A1DA1;
wire signed [6:0] C1DB1;
wire A1DB1;
wire signed [6:0] C1DC1;
wire A1DC1;
wire signed [6:0] C1DD1;
wire A1DD1;
wire signed [6:0] C1002;
wire A1002;
wire signed [6:0] C1012;
wire A1012;
wire signed [6:0] C1022;
wire A1022;
wire signed [6:0] C1032;
wire A1032;
wire signed [6:0] C1042;
wire A1042;
wire signed [6:0] C1052;
wire A1052;
wire signed [6:0] C1062;
wire A1062;
wire signed [6:0] C1072;
wire A1072;
wire signed [6:0] C1082;
wire A1082;
wire signed [6:0] C1092;
wire A1092;
wire signed [6:0] C10A2;
wire A10A2;
wire signed [6:0] C10B2;
wire A10B2;
wire signed [6:0] C10C2;
wire A10C2;
wire signed [6:0] C10D2;
wire A10D2;
wire signed [6:0] C1102;
wire A1102;
wire signed [6:0] C1112;
wire A1112;
wire signed [6:0] C1122;
wire A1122;
wire signed [6:0] C1132;
wire A1132;
wire signed [6:0] C1142;
wire A1142;
wire signed [6:0] C1152;
wire A1152;
wire signed [6:0] C1162;
wire A1162;
wire signed [6:0] C1172;
wire A1172;
wire signed [6:0] C1182;
wire A1182;
wire signed [6:0] C1192;
wire A1192;
wire signed [6:0] C11A2;
wire A11A2;
wire signed [6:0] C11B2;
wire A11B2;
wire signed [6:0] C11C2;
wire A11C2;
wire signed [6:0] C11D2;
wire A11D2;
wire signed [6:0] C1202;
wire A1202;
wire signed [6:0] C1212;
wire A1212;
wire signed [6:0] C1222;
wire A1222;
wire signed [6:0] C1232;
wire A1232;
wire signed [6:0] C1242;
wire A1242;
wire signed [6:0] C1252;
wire A1252;
wire signed [6:0] C1262;
wire A1262;
wire signed [6:0] C1272;
wire A1272;
wire signed [6:0] C1282;
wire A1282;
wire signed [6:0] C1292;
wire A1292;
wire signed [6:0] C12A2;
wire A12A2;
wire signed [6:0] C12B2;
wire A12B2;
wire signed [6:0] C12C2;
wire A12C2;
wire signed [6:0] C12D2;
wire A12D2;
wire signed [6:0] C1302;
wire A1302;
wire signed [6:0] C1312;
wire A1312;
wire signed [6:0] C1322;
wire A1322;
wire signed [6:0] C1332;
wire A1332;
wire signed [6:0] C1342;
wire A1342;
wire signed [6:0] C1352;
wire A1352;
wire signed [6:0] C1362;
wire A1362;
wire signed [6:0] C1372;
wire A1372;
wire signed [6:0] C1382;
wire A1382;
wire signed [6:0] C1392;
wire A1392;
wire signed [6:0] C13A2;
wire A13A2;
wire signed [6:0] C13B2;
wire A13B2;
wire signed [6:0] C13C2;
wire A13C2;
wire signed [6:0] C13D2;
wire A13D2;
wire signed [6:0] C1402;
wire A1402;
wire signed [6:0] C1412;
wire A1412;
wire signed [6:0] C1422;
wire A1422;
wire signed [6:0] C1432;
wire A1432;
wire signed [6:0] C1442;
wire A1442;
wire signed [6:0] C1452;
wire A1452;
wire signed [6:0] C1462;
wire A1462;
wire signed [6:0] C1472;
wire A1472;
wire signed [6:0] C1482;
wire A1482;
wire signed [6:0] C1492;
wire A1492;
wire signed [6:0] C14A2;
wire A14A2;
wire signed [6:0] C14B2;
wire A14B2;
wire signed [6:0] C14C2;
wire A14C2;
wire signed [6:0] C14D2;
wire A14D2;
wire signed [6:0] C1502;
wire A1502;
wire signed [6:0] C1512;
wire A1512;
wire signed [6:0] C1522;
wire A1522;
wire signed [6:0] C1532;
wire A1532;
wire signed [6:0] C1542;
wire A1542;
wire signed [6:0] C1552;
wire A1552;
wire signed [6:0] C1562;
wire A1562;
wire signed [6:0] C1572;
wire A1572;
wire signed [6:0] C1582;
wire A1582;
wire signed [6:0] C1592;
wire A1592;
wire signed [6:0] C15A2;
wire A15A2;
wire signed [6:0] C15B2;
wire A15B2;
wire signed [6:0] C15C2;
wire A15C2;
wire signed [6:0] C15D2;
wire A15D2;
wire signed [6:0] C1602;
wire A1602;
wire signed [6:0] C1612;
wire A1612;
wire signed [6:0] C1622;
wire A1622;
wire signed [6:0] C1632;
wire A1632;
wire signed [6:0] C1642;
wire A1642;
wire signed [6:0] C1652;
wire A1652;
wire signed [6:0] C1662;
wire A1662;
wire signed [6:0] C1672;
wire A1672;
wire signed [6:0] C1682;
wire A1682;
wire signed [6:0] C1692;
wire A1692;
wire signed [6:0] C16A2;
wire A16A2;
wire signed [6:0] C16B2;
wire A16B2;
wire signed [6:0] C16C2;
wire A16C2;
wire signed [6:0] C16D2;
wire A16D2;
wire signed [6:0] C1702;
wire A1702;
wire signed [6:0] C1712;
wire A1712;
wire signed [6:0] C1722;
wire A1722;
wire signed [6:0] C1732;
wire A1732;
wire signed [6:0] C1742;
wire A1742;
wire signed [6:0] C1752;
wire A1752;
wire signed [6:0] C1762;
wire A1762;
wire signed [6:0] C1772;
wire A1772;
wire signed [6:0] C1782;
wire A1782;
wire signed [6:0] C1792;
wire A1792;
wire signed [6:0] C17A2;
wire A17A2;
wire signed [6:0] C17B2;
wire A17B2;
wire signed [6:0] C17C2;
wire A17C2;
wire signed [6:0] C17D2;
wire A17D2;
wire signed [6:0] C1802;
wire A1802;
wire signed [6:0] C1812;
wire A1812;
wire signed [6:0] C1822;
wire A1822;
wire signed [6:0] C1832;
wire A1832;
wire signed [6:0] C1842;
wire A1842;
wire signed [6:0] C1852;
wire A1852;
wire signed [6:0] C1862;
wire A1862;
wire signed [6:0] C1872;
wire A1872;
wire signed [6:0] C1882;
wire A1882;
wire signed [6:0] C1892;
wire A1892;
wire signed [6:0] C18A2;
wire A18A2;
wire signed [6:0] C18B2;
wire A18B2;
wire signed [6:0] C18C2;
wire A18C2;
wire signed [6:0] C18D2;
wire A18D2;
wire signed [6:0] C1902;
wire A1902;
wire signed [6:0] C1912;
wire A1912;
wire signed [6:0] C1922;
wire A1922;
wire signed [6:0] C1932;
wire A1932;
wire signed [6:0] C1942;
wire A1942;
wire signed [6:0] C1952;
wire A1952;
wire signed [6:0] C1962;
wire A1962;
wire signed [6:0] C1972;
wire A1972;
wire signed [6:0] C1982;
wire A1982;
wire signed [6:0] C1992;
wire A1992;
wire signed [6:0] C19A2;
wire A19A2;
wire signed [6:0] C19B2;
wire A19B2;
wire signed [6:0] C19C2;
wire A19C2;
wire signed [6:0] C19D2;
wire A19D2;
wire signed [6:0] C1A02;
wire A1A02;
wire signed [6:0] C1A12;
wire A1A12;
wire signed [6:0] C1A22;
wire A1A22;
wire signed [6:0] C1A32;
wire A1A32;
wire signed [6:0] C1A42;
wire A1A42;
wire signed [6:0] C1A52;
wire A1A52;
wire signed [6:0] C1A62;
wire A1A62;
wire signed [6:0] C1A72;
wire A1A72;
wire signed [6:0] C1A82;
wire A1A82;
wire signed [6:0] C1A92;
wire A1A92;
wire signed [6:0] C1AA2;
wire A1AA2;
wire signed [6:0] C1AB2;
wire A1AB2;
wire signed [6:0] C1AC2;
wire A1AC2;
wire signed [6:0] C1AD2;
wire A1AD2;
wire signed [6:0] C1B02;
wire A1B02;
wire signed [6:0] C1B12;
wire A1B12;
wire signed [6:0] C1B22;
wire A1B22;
wire signed [6:0] C1B32;
wire A1B32;
wire signed [6:0] C1B42;
wire A1B42;
wire signed [6:0] C1B52;
wire A1B52;
wire signed [6:0] C1B62;
wire A1B62;
wire signed [6:0] C1B72;
wire A1B72;
wire signed [6:0] C1B82;
wire A1B82;
wire signed [6:0] C1B92;
wire A1B92;
wire signed [6:0] C1BA2;
wire A1BA2;
wire signed [6:0] C1BB2;
wire A1BB2;
wire signed [6:0] C1BC2;
wire A1BC2;
wire signed [6:0] C1BD2;
wire A1BD2;
wire signed [6:0] C1C02;
wire A1C02;
wire signed [6:0] C1C12;
wire A1C12;
wire signed [6:0] C1C22;
wire A1C22;
wire signed [6:0] C1C32;
wire A1C32;
wire signed [6:0] C1C42;
wire A1C42;
wire signed [6:0] C1C52;
wire A1C52;
wire signed [6:0] C1C62;
wire A1C62;
wire signed [6:0] C1C72;
wire A1C72;
wire signed [6:0] C1C82;
wire A1C82;
wire signed [6:0] C1C92;
wire A1C92;
wire signed [6:0] C1CA2;
wire A1CA2;
wire signed [6:0] C1CB2;
wire A1CB2;
wire signed [6:0] C1CC2;
wire A1CC2;
wire signed [6:0] C1CD2;
wire A1CD2;
wire signed [6:0] C1D02;
wire A1D02;
wire signed [6:0] C1D12;
wire A1D12;
wire signed [6:0] C1D22;
wire A1D22;
wire signed [6:0] C1D32;
wire A1D32;
wire signed [6:0] C1D42;
wire A1D42;
wire signed [6:0] C1D52;
wire A1D52;
wire signed [6:0] C1D62;
wire A1D62;
wire signed [6:0] C1D72;
wire A1D72;
wire signed [6:0] C1D82;
wire A1D82;
wire signed [6:0] C1D92;
wire A1D92;
wire signed [6:0] C1DA2;
wire A1DA2;
wire signed [6:0] C1DB2;
wire A1DB2;
wire signed [6:0] C1DC2;
wire A1DC2;
wire signed [6:0] C1DD2;
wire A1DD2;
wire signed [6:0] C1003;
wire A1003;
wire signed [6:0] C1013;
wire A1013;
wire signed [6:0] C1023;
wire A1023;
wire signed [6:0] C1033;
wire A1033;
wire signed [6:0] C1043;
wire A1043;
wire signed [6:0] C1053;
wire A1053;
wire signed [6:0] C1063;
wire A1063;
wire signed [6:0] C1073;
wire A1073;
wire signed [6:0] C1083;
wire A1083;
wire signed [6:0] C1093;
wire A1093;
wire signed [6:0] C10A3;
wire A10A3;
wire signed [6:0] C10B3;
wire A10B3;
wire signed [6:0] C10C3;
wire A10C3;
wire signed [6:0] C10D3;
wire A10D3;
wire signed [6:0] C1103;
wire A1103;
wire signed [6:0] C1113;
wire A1113;
wire signed [6:0] C1123;
wire A1123;
wire signed [6:0] C1133;
wire A1133;
wire signed [6:0] C1143;
wire A1143;
wire signed [6:0] C1153;
wire A1153;
wire signed [6:0] C1163;
wire A1163;
wire signed [6:0] C1173;
wire A1173;
wire signed [6:0] C1183;
wire A1183;
wire signed [6:0] C1193;
wire A1193;
wire signed [6:0] C11A3;
wire A11A3;
wire signed [6:0] C11B3;
wire A11B3;
wire signed [6:0] C11C3;
wire A11C3;
wire signed [6:0] C11D3;
wire A11D3;
wire signed [6:0] C1203;
wire A1203;
wire signed [6:0] C1213;
wire A1213;
wire signed [6:0] C1223;
wire A1223;
wire signed [6:0] C1233;
wire A1233;
wire signed [6:0] C1243;
wire A1243;
wire signed [6:0] C1253;
wire A1253;
wire signed [6:0] C1263;
wire A1263;
wire signed [6:0] C1273;
wire A1273;
wire signed [6:0] C1283;
wire A1283;
wire signed [6:0] C1293;
wire A1293;
wire signed [6:0] C12A3;
wire A12A3;
wire signed [6:0] C12B3;
wire A12B3;
wire signed [6:0] C12C3;
wire A12C3;
wire signed [6:0] C12D3;
wire A12D3;
wire signed [6:0] C1303;
wire A1303;
wire signed [6:0] C1313;
wire A1313;
wire signed [6:0] C1323;
wire A1323;
wire signed [6:0] C1333;
wire A1333;
wire signed [6:0] C1343;
wire A1343;
wire signed [6:0] C1353;
wire A1353;
wire signed [6:0] C1363;
wire A1363;
wire signed [6:0] C1373;
wire A1373;
wire signed [6:0] C1383;
wire A1383;
wire signed [6:0] C1393;
wire A1393;
wire signed [6:0] C13A3;
wire A13A3;
wire signed [6:0] C13B3;
wire A13B3;
wire signed [6:0] C13C3;
wire A13C3;
wire signed [6:0] C13D3;
wire A13D3;
wire signed [6:0] C1403;
wire A1403;
wire signed [6:0] C1413;
wire A1413;
wire signed [6:0] C1423;
wire A1423;
wire signed [6:0] C1433;
wire A1433;
wire signed [6:0] C1443;
wire A1443;
wire signed [6:0] C1453;
wire A1453;
wire signed [6:0] C1463;
wire A1463;
wire signed [6:0] C1473;
wire A1473;
wire signed [6:0] C1483;
wire A1483;
wire signed [6:0] C1493;
wire A1493;
wire signed [6:0] C14A3;
wire A14A3;
wire signed [6:0] C14B3;
wire A14B3;
wire signed [6:0] C14C3;
wire A14C3;
wire signed [6:0] C14D3;
wire A14D3;
wire signed [6:0] C1503;
wire A1503;
wire signed [6:0] C1513;
wire A1513;
wire signed [6:0] C1523;
wire A1523;
wire signed [6:0] C1533;
wire A1533;
wire signed [6:0] C1543;
wire A1543;
wire signed [6:0] C1553;
wire A1553;
wire signed [6:0] C1563;
wire A1563;
wire signed [6:0] C1573;
wire A1573;
wire signed [6:0] C1583;
wire A1583;
wire signed [6:0] C1593;
wire A1593;
wire signed [6:0] C15A3;
wire A15A3;
wire signed [6:0] C15B3;
wire A15B3;
wire signed [6:0] C15C3;
wire A15C3;
wire signed [6:0] C15D3;
wire A15D3;
wire signed [6:0] C1603;
wire A1603;
wire signed [6:0] C1613;
wire A1613;
wire signed [6:0] C1623;
wire A1623;
wire signed [6:0] C1633;
wire A1633;
wire signed [6:0] C1643;
wire A1643;
wire signed [6:0] C1653;
wire A1653;
wire signed [6:0] C1663;
wire A1663;
wire signed [6:0] C1673;
wire A1673;
wire signed [6:0] C1683;
wire A1683;
wire signed [6:0] C1693;
wire A1693;
wire signed [6:0] C16A3;
wire A16A3;
wire signed [6:0] C16B3;
wire A16B3;
wire signed [6:0] C16C3;
wire A16C3;
wire signed [6:0] C16D3;
wire A16D3;
wire signed [6:0] C1703;
wire A1703;
wire signed [6:0] C1713;
wire A1713;
wire signed [6:0] C1723;
wire A1723;
wire signed [6:0] C1733;
wire A1733;
wire signed [6:0] C1743;
wire A1743;
wire signed [6:0] C1753;
wire A1753;
wire signed [6:0] C1763;
wire A1763;
wire signed [6:0] C1773;
wire A1773;
wire signed [6:0] C1783;
wire A1783;
wire signed [6:0] C1793;
wire A1793;
wire signed [6:0] C17A3;
wire A17A3;
wire signed [6:0] C17B3;
wire A17B3;
wire signed [6:0] C17C3;
wire A17C3;
wire signed [6:0] C17D3;
wire A17D3;
wire signed [6:0] C1803;
wire A1803;
wire signed [6:0] C1813;
wire A1813;
wire signed [6:0] C1823;
wire A1823;
wire signed [6:0] C1833;
wire A1833;
wire signed [6:0] C1843;
wire A1843;
wire signed [6:0] C1853;
wire A1853;
wire signed [6:0] C1863;
wire A1863;
wire signed [6:0] C1873;
wire A1873;
wire signed [6:0] C1883;
wire A1883;
wire signed [6:0] C1893;
wire A1893;
wire signed [6:0] C18A3;
wire A18A3;
wire signed [6:0] C18B3;
wire A18B3;
wire signed [6:0] C18C3;
wire A18C3;
wire signed [6:0] C18D3;
wire A18D3;
wire signed [6:0] C1903;
wire A1903;
wire signed [6:0] C1913;
wire A1913;
wire signed [6:0] C1923;
wire A1923;
wire signed [6:0] C1933;
wire A1933;
wire signed [6:0] C1943;
wire A1943;
wire signed [6:0] C1953;
wire A1953;
wire signed [6:0] C1963;
wire A1963;
wire signed [6:0] C1973;
wire A1973;
wire signed [6:0] C1983;
wire A1983;
wire signed [6:0] C1993;
wire A1993;
wire signed [6:0] C19A3;
wire A19A3;
wire signed [6:0] C19B3;
wire A19B3;
wire signed [6:0] C19C3;
wire A19C3;
wire signed [6:0] C19D3;
wire A19D3;
wire signed [6:0] C1A03;
wire A1A03;
wire signed [6:0] C1A13;
wire A1A13;
wire signed [6:0] C1A23;
wire A1A23;
wire signed [6:0] C1A33;
wire A1A33;
wire signed [6:0] C1A43;
wire A1A43;
wire signed [6:0] C1A53;
wire A1A53;
wire signed [6:0] C1A63;
wire A1A63;
wire signed [6:0] C1A73;
wire A1A73;
wire signed [6:0] C1A83;
wire A1A83;
wire signed [6:0] C1A93;
wire A1A93;
wire signed [6:0] C1AA3;
wire A1AA3;
wire signed [6:0] C1AB3;
wire A1AB3;
wire signed [6:0] C1AC3;
wire A1AC3;
wire signed [6:0] C1AD3;
wire A1AD3;
wire signed [6:0] C1B03;
wire A1B03;
wire signed [6:0] C1B13;
wire A1B13;
wire signed [6:0] C1B23;
wire A1B23;
wire signed [6:0] C1B33;
wire A1B33;
wire signed [6:0] C1B43;
wire A1B43;
wire signed [6:0] C1B53;
wire A1B53;
wire signed [6:0] C1B63;
wire A1B63;
wire signed [6:0] C1B73;
wire A1B73;
wire signed [6:0] C1B83;
wire A1B83;
wire signed [6:0] C1B93;
wire A1B93;
wire signed [6:0] C1BA3;
wire A1BA3;
wire signed [6:0] C1BB3;
wire A1BB3;
wire signed [6:0] C1BC3;
wire A1BC3;
wire signed [6:0] C1BD3;
wire A1BD3;
wire signed [6:0] C1C03;
wire A1C03;
wire signed [6:0] C1C13;
wire A1C13;
wire signed [6:0] C1C23;
wire A1C23;
wire signed [6:0] C1C33;
wire A1C33;
wire signed [6:0] C1C43;
wire A1C43;
wire signed [6:0] C1C53;
wire A1C53;
wire signed [6:0] C1C63;
wire A1C63;
wire signed [6:0] C1C73;
wire A1C73;
wire signed [6:0] C1C83;
wire A1C83;
wire signed [6:0] C1C93;
wire A1C93;
wire signed [6:0] C1CA3;
wire A1CA3;
wire signed [6:0] C1CB3;
wire A1CB3;
wire signed [6:0] C1CC3;
wire A1CC3;
wire signed [6:0] C1CD3;
wire A1CD3;
wire signed [6:0] C1D03;
wire A1D03;
wire signed [6:0] C1D13;
wire A1D13;
wire signed [6:0] C1D23;
wire A1D23;
wire signed [6:0] C1D33;
wire A1D33;
wire signed [6:0] C1D43;
wire A1D43;
wire signed [6:0] C1D53;
wire A1D53;
wire signed [6:0] C1D63;
wire A1D63;
wire signed [6:0] C1D73;
wire A1D73;
wire signed [6:0] C1D83;
wire A1D83;
wire signed [6:0] C1D93;
wire A1D93;
wire signed [6:0] C1DA3;
wire A1DA3;
wire signed [6:0] C1DB3;
wire A1DB3;
wire signed [6:0] C1DC3;
wire A1DC3;
wire signed [6:0] C1DD3;
wire A1DD3;
wire signed [6:0] C1004;
wire A1004;
wire signed [6:0] C1014;
wire A1014;
wire signed [6:0] C1024;
wire A1024;
wire signed [6:0] C1034;
wire A1034;
wire signed [6:0] C1044;
wire A1044;
wire signed [6:0] C1054;
wire A1054;
wire signed [6:0] C1064;
wire A1064;
wire signed [6:0] C1074;
wire A1074;
wire signed [6:0] C1084;
wire A1084;
wire signed [6:0] C1094;
wire A1094;
wire signed [6:0] C10A4;
wire A10A4;
wire signed [6:0] C10B4;
wire A10B4;
wire signed [6:0] C10C4;
wire A10C4;
wire signed [6:0] C10D4;
wire A10D4;
wire signed [6:0] C1104;
wire A1104;
wire signed [6:0] C1114;
wire A1114;
wire signed [6:0] C1124;
wire A1124;
wire signed [6:0] C1134;
wire A1134;
wire signed [6:0] C1144;
wire A1144;
wire signed [6:0] C1154;
wire A1154;
wire signed [6:0] C1164;
wire A1164;
wire signed [6:0] C1174;
wire A1174;
wire signed [6:0] C1184;
wire A1184;
wire signed [6:0] C1194;
wire A1194;
wire signed [6:0] C11A4;
wire A11A4;
wire signed [6:0] C11B4;
wire A11B4;
wire signed [6:0] C11C4;
wire A11C4;
wire signed [6:0] C11D4;
wire A11D4;
wire signed [6:0] C1204;
wire A1204;
wire signed [6:0] C1214;
wire A1214;
wire signed [6:0] C1224;
wire A1224;
wire signed [6:0] C1234;
wire A1234;
wire signed [6:0] C1244;
wire A1244;
wire signed [6:0] C1254;
wire A1254;
wire signed [6:0] C1264;
wire A1264;
wire signed [6:0] C1274;
wire A1274;
wire signed [6:0] C1284;
wire A1284;
wire signed [6:0] C1294;
wire A1294;
wire signed [6:0] C12A4;
wire A12A4;
wire signed [6:0] C12B4;
wire A12B4;
wire signed [6:0] C12C4;
wire A12C4;
wire signed [6:0] C12D4;
wire A12D4;
wire signed [6:0] C1304;
wire A1304;
wire signed [6:0] C1314;
wire A1314;
wire signed [6:0] C1324;
wire A1324;
wire signed [6:0] C1334;
wire A1334;
wire signed [6:0] C1344;
wire A1344;
wire signed [6:0] C1354;
wire A1354;
wire signed [6:0] C1364;
wire A1364;
wire signed [6:0] C1374;
wire A1374;
wire signed [6:0] C1384;
wire A1384;
wire signed [6:0] C1394;
wire A1394;
wire signed [6:0] C13A4;
wire A13A4;
wire signed [6:0] C13B4;
wire A13B4;
wire signed [6:0] C13C4;
wire A13C4;
wire signed [6:0] C13D4;
wire A13D4;
wire signed [6:0] C1404;
wire A1404;
wire signed [6:0] C1414;
wire A1414;
wire signed [6:0] C1424;
wire A1424;
wire signed [6:0] C1434;
wire A1434;
wire signed [6:0] C1444;
wire A1444;
wire signed [6:0] C1454;
wire A1454;
wire signed [6:0] C1464;
wire A1464;
wire signed [6:0] C1474;
wire A1474;
wire signed [6:0] C1484;
wire A1484;
wire signed [6:0] C1494;
wire A1494;
wire signed [6:0] C14A4;
wire A14A4;
wire signed [6:0] C14B4;
wire A14B4;
wire signed [6:0] C14C4;
wire A14C4;
wire signed [6:0] C14D4;
wire A14D4;
wire signed [6:0] C1504;
wire A1504;
wire signed [6:0] C1514;
wire A1514;
wire signed [6:0] C1524;
wire A1524;
wire signed [6:0] C1534;
wire A1534;
wire signed [6:0] C1544;
wire A1544;
wire signed [6:0] C1554;
wire A1554;
wire signed [6:0] C1564;
wire A1564;
wire signed [6:0] C1574;
wire A1574;
wire signed [6:0] C1584;
wire A1584;
wire signed [6:0] C1594;
wire A1594;
wire signed [6:0] C15A4;
wire A15A4;
wire signed [6:0] C15B4;
wire A15B4;
wire signed [6:0] C15C4;
wire A15C4;
wire signed [6:0] C15D4;
wire A15D4;
wire signed [6:0] C1604;
wire A1604;
wire signed [6:0] C1614;
wire A1614;
wire signed [6:0] C1624;
wire A1624;
wire signed [6:0] C1634;
wire A1634;
wire signed [6:0] C1644;
wire A1644;
wire signed [6:0] C1654;
wire A1654;
wire signed [6:0] C1664;
wire A1664;
wire signed [6:0] C1674;
wire A1674;
wire signed [6:0] C1684;
wire A1684;
wire signed [6:0] C1694;
wire A1694;
wire signed [6:0] C16A4;
wire A16A4;
wire signed [6:0] C16B4;
wire A16B4;
wire signed [6:0] C16C4;
wire A16C4;
wire signed [6:0] C16D4;
wire A16D4;
wire signed [6:0] C1704;
wire A1704;
wire signed [6:0] C1714;
wire A1714;
wire signed [6:0] C1724;
wire A1724;
wire signed [6:0] C1734;
wire A1734;
wire signed [6:0] C1744;
wire A1744;
wire signed [6:0] C1754;
wire A1754;
wire signed [6:0] C1764;
wire A1764;
wire signed [6:0] C1774;
wire A1774;
wire signed [6:0] C1784;
wire A1784;
wire signed [6:0] C1794;
wire A1794;
wire signed [6:0] C17A4;
wire A17A4;
wire signed [6:0] C17B4;
wire A17B4;
wire signed [6:0] C17C4;
wire A17C4;
wire signed [6:0] C17D4;
wire A17D4;
wire signed [6:0] C1804;
wire A1804;
wire signed [6:0] C1814;
wire A1814;
wire signed [6:0] C1824;
wire A1824;
wire signed [6:0] C1834;
wire A1834;
wire signed [6:0] C1844;
wire A1844;
wire signed [6:0] C1854;
wire A1854;
wire signed [6:0] C1864;
wire A1864;
wire signed [6:0] C1874;
wire A1874;
wire signed [6:0] C1884;
wire A1884;
wire signed [6:0] C1894;
wire A1894;
wire signed [6:0] C18A4;
wire A18A4;
wire signed [6:0] C18B4;
wire A18B4;
wire signed [6:0] C18C4;
wire A18C4;
wire signed [6:0] C18D4;
wire A18D4;
wire signed [6:0] C1904;
wire A1904;
wire signed [6:0] C1914;
wire A1914;
wire signed [6:0] C1924;
wire A1924;
wire signed [6:0] C1934;
wire A1934;
wire signed [6:0] C1944;
wire A1944;
wire signed [6:0] C1954;
wire A1954;
wire signed [6:0] C1964;
wire A1964;
wire signed [6:0] C1974;
wire A1974;
wire signed [6:0] C1984;
wire A1984;
wire signed [6:0] C1994;
wire A1994;
wire signed [6:0] C19A4;
wire A19A4;
wire signed [6:0] C19B4;
wire A19B4;
wire signed [6:0] C19C4;
wire A19C4;
wire signed [6:0] C19D4;
wire A19D4;
wire signed [6:0] C1A04;
wire A1A04;
wire signed [6:0] C1A14;
wire A1A14;
wire signed [6:0] C1A24;
wire A1A24;
wire signed [6:0] C1A34;
wire A1A34;
wire signed [6:0] C1A44;
wire A1A44;
wire signed [6:0] C1A54;
wire A1A54;
wire signed [6:0] C1A64;
wire A1A64;
wire signed [6:0] C1A74;
wire A1A74;
wire signed [6:0] C1A84;
wire A1A84;
wire signed [6:0] C1A94;
wire A1A94;
wire signed [6:0] C1AA4;
wire A1AA4;
wire signed [6:0] C1AB4;
wire A1AB4;
wire signed [6:0] C1AC4;
wire A1AC4;
wire signed [6:0] C1AD4;
wire A1AD4;
wire signed [6:0] C1B04;
wire A1B04;
wire signed [6:0] C1B14;
wire A1B14;
wire signed [6:0] C1B24;
wire A1B24;
wire signed [6:0] C1B34;
wire A1B34;
wire signed [6:0] C1B44;
wire A1B44;
wire signed [6:0] C1B54;
wire A1B54;
wire signed [6:0] C1B64;
wire A1B64;
wire signed [6:0] C1B74;
wire A1B74;
wire signed [6:0] C1B84;
wire A1B84;
wire signed [6:0] C1B94;
wire A1B94;
wire signed [6:0] C1BA4;
wire A1BA4;
wire signed [6:0] C1BB4;
wire A1BB4;
wire signed [6:0] C1BC4;
wire A1BC4;
wire signed [6:0] C1BD4;
wire A1BD4;
wire signed [6:0] C1C04;
wire A1C04;
wire signed [6:0] C1C14;
wire A1C14;
wire signed [6:0] C1C24;
wire A1C24;
wire signed [6:0] C1C34;
wire A1C34;
wire signed [6:0] C1C44;
wire A1C44;
wire signed [6:0] C1C54;
wire A1C54;
wire signed [6:0] C1C64;
wire A1C64;
wire signed [6:0] C1C74;
wire A1C74;
wire signed [6:0] C1C84;
wire A1C84;
wire signed [6:0] C1C94;
wire A1C94;
wire signed [6:0] C1CA4;
wire A1CA4;
wire signed [6:0] C1CB4;
wire A1CB4;
wire signed [6:0] C1CC4;
wire A1CC4;
wire signed [6:0] C1CD4;
wire A1CD4;
wire signed [6:0] C1D04;
wire A1D04;
wire signed [6:0] C1D14;
wire A1D14;
wire signed [6:0] C1D24;
wire A1D24;
wire signed [6:0] C1D34;
wire A1D34;
wire signed [6:0] C1D44;
wire A1D44;
wire signed [6:0] C1D54;
wire A1D54;
wire signed [6:0] C1D64;
wire A1D64;
wire signed [6:0] C1D74;
wire A1D74;
wire signed [6:0] C1D84;
wire A1D84;
wire signed [6:0] C1D94;
wire A1D94;
wire signed [6:0] C1DA4;
wire A1DA4;
wire signed [6:0] C1DB4;
wire A1DB4;
wire signed [6:0] C1DC4;
wire A1DC4;
wire signed [6:0] C1DD4;
wire A1DD4;
wire signed [6:0] C1005;
wire A1005;
wire signed [6:0] C1015;
wire A1015;
wire signed [6:0] C1025;
wire A1025;
wire signed [6:0] C1035;
wire A1035;
wire signed [6:0] C1045;
wire A1045;
wire signed [6:0] C1055;
wire A1055;
wire signed [6:0] C1065;
wire A1065;
wire signed [6:0] C1075;
wire A1075;
wire signed [6:0] C1085;
wire A1085;
wire signed [6:0] C1095;
wire A1095;
wire signed [6:0] C10A5;
wire A10A5;
wire signed [6:0] C10B5;
wire A10B5;
wire signed [6:0] C10C5;
wire A10C5;
wire signed [6:0] C10D5;
wire A10D5;
wire signed [6:0] C1105;
wire A1105;
wire signed [6:0] C1115;
wire A1115;
wire signed [6:0] C1125;
wire A1125;
wire signed [6:0] C1135;
wire A1135;
wire signed [6:0] C1145;
wire A1145;
wire signed [6:0] C1155;
wire A1155;
wire signed [6:0] C1165;
wire A1165;
wire signed [6:0] C1175;
wire A1175;
wire signed [6:0] C1185;
wire A1185;
wire signed [6:0] C1195;
wire A1195;
wire signed [6:0] C11A5;
wire A11A5;
wire signed [6:0] C11B5;
wire A11B5;
wire signed [6:0] C11C5;
wire A11C5;
wire signed [6:0] C11D5;
wire A11D5;
wire signed [6:0] C1205;
wire A1205;
wire signed [6:0] C1215;
wire A1215;
wire signed [6:0] C1225;
wire A1225;
wire signed [6:0] C1235;
wire A1235;
wire signed [6:0] C1245;
wire A1245;
wire signed [6:0] C1255;
wire A1255;
wire signed [6:0] C1265;
wire A1265;
wire signed [6:0] C1275;
wire A1275;
wire signed [6:0] C1285;
wire A1285;
wire signed [6:0] C1295;
wire A1295;
wire signed [6:0] C12A5;
wire A12A5;
wire signed [6:0] C12B5;
wire A12B5;
wire signed [6:0] C12C5;
wire A12C5;
wire signed [6:0] C12D5;
wire A12D5;
wire signed [6:0] C1305;
wire A1305;
wire signed [6:0] C1315;
wire A1315;
wire signed [6:0] C1325;
wire A1325;
wire signed [6:0] C1335;
wire A1335;
wire signed [6:0] C1345;
wire A1345;
wire signed [6:0] C1355;
wire A1355;
wire signed [6:0] C1365;
wire A1365;
wire signed [6:0] C1375;
wire A1375;
wire signed [6:0] C1385;
wire A1385;
wire signed [6:0] C1395;
wire A1395;
wire signed [6:0] C13A5;
wire A13A5;
wire signed [6:0] C13B5;
wire A13B5;
wire signed [6:0] C13C5;
wire A13C5;
wire signed [6:0] C13D5;
wire A13D5;
wire signed [6:0] C1405;
wire A1405;
wire signed [6:0] C1415;
wire A1415;
wire signed [6:0] C1425;
wire A1425;
wire signed [6:0] C1435;
wire A1435;
wire signed [6:0] C1445;
wire A1445;
wire signed [6:0] C1455;
wire A1455;
wire signed [6:0] C1465;
wire A1465;
wire signed [6:0] C1475;
wire A1475;
wire signed [6:0] C1485;
wire A1485;
wire signed [6:0] C1495;
wire A1495;
wire signed [6:0] C14A5;
wire A14A5;
wire signed [6:0] C14B5;
wire A14B5;
wire signed [6:0] C14C5;
wire A14C5;
wire signed [6:0] C14D5;
wire A14D5;
wire signed [6:0] C1505;
wire A1505;
wire signed [6:0] C1515;
wire A1515;
wire signed [6:0] C1525;
wire A1525;
wire signed [6:0] C1535;
wire A1535;
wire signed [6:0] C1545;
wire A1545;
wire signed [6:0] C1555;
wire A1555;
wire signed [6:0] C1565;
wire A1565;
wire signed [6:0] C1575;
wire A1575;
wire signed [6:0] C1585;
wire A1585;
wire signed [6:0] C1595;
wire A1595;
wire signed [6:0] C15A5;
wire A15A5;
wire signed [6:0] C15B5;
wire A15B5;
wire signed [6:0] C15C5;
wire A15C5;
wire signed [6:0] C15D5;
wire A15D5;
wire signed [6:0] C1605;
wire A1605;
wire signed [6:0] C1615;
wire A1615;
wire signed [6:0] C1625;
wire A1625;
wire signed [6:0] C1635;
wire A1635;
wire signed [6:0] C1645;
wire A1645;
wire signed [6:0] C1655;
wire A1655;
wire signed [6:0] C1665;
wire A1665;
wire signed [6:0] C1675;
wire A1675;
wire signed [6:0] C1685;
wire A1685;
wire signed [6:0] C1695;
wire A1695;
wire signed [6:0] C16A5;
wire A16A5;
wire signed [6:0] C16B5;
wire A16B5;
wire signed [6:0] C16C5;
wire A16C5;
wire signed [6:0] C16D5;
wire A16D5;
wire signed [6:0] C1705;
wire A1705;
wire signed [6:0] C1715;
wire A1715;
wire signed [6:0] C1725;
wire A1725;
wire signed [6:0] C1735;
wire A1735;
wire signed [6:0] C1745;
wire A1745;
wire signed [6:0] C1755;
wire A1755;
wire signed [6:0] C1765;
wire A1765;
wire signed [6:0] C1775;
wire A1775;
wire signed [6:0] C1785;
wire A1785;
wire signed [6:0] C1795;
wire A1795;
wire signed [6:0] C17A5;
wire A17A5;
wire signed [6:0] C17B5;
wire A17B5;
wire signed [6:0] C17C5;
wire A17C5;
wire signed [6:0] C17D5;
wire A17D5;
wire signed [6:0] C1805;
wire A1805;
wire signed [6:0] C1815;
wire A1815;
wire signed [6:0] C1825;
wire A1825;
wire signed [6:0] C1835;
wire A1835;
wire signed [6:0] C1845;
wire A1845;
wire signed [6:0] C1855;
wire A1855;
wire signed [6:0] C1865;
wire A1865;
wire signed [6:0] C1875;
wire A1875;
wire signed [6:0] C1885;
wire A1885;
wire signed [6:0] C1895;
wire A1895;
wire signed [6:0] C18A5;
wire A18A5;
wire signed [6:0] C18B5;
wire A18B5;
wire signed [6:0] C18C5;
wire A18C5;
wire signed [6:0] C18D5;
wire A18D5;
wire signed [6:0] C1905;
wire A1905;
wire signed [6:0] C1915;
wire A1915;
wire signed [6:0] C1925;
wire A1925;
wire signed [6:0] C1935;
wire A1935;
wire signed [6:0] C1945;
wire A1945;
wire signed [6:0] C1955;
wire A1955;
wire signed [6:0] C1965;
wire A1965;
wire signed [6:0] C1975;
wire A1975;
wire signed [6:0] C1985;
wire A1985;
wire signed [6:0] C1995;
wire A1995;
wire signed [6:0] C19A5;
wire A19A5;
wire signed [6:0] C19B5;
wire A19B5;
wire signed [6:0] C19C5;
wire A19C5;
wire signed [6:0] C19D5;
wire A19D5;
wire signed [6:0] C1A05;
wire A1A05;
wire signed [6:0] C1A15;
wire A1A15;
wire signed [6:0] C1A25;
wire A1A25;
wire signed [6:0] C1A35;
wire A1A35;
wire signed [6:0] C1A45;
wire A1A45;
wire signed [6:0] C1A55;
wire A1A55;
wire signed [6:0] C1A65;
wire A1A65;
wire signed [6:0] C1A75;
wire A1A75;
wire signed [6:0] C1A85;
wire A1A85;
wire signed [6:0] C1A95;
wire A1A95;
wire signed [6:0] C1AA5;
wire A1AA5;
wire signed [6:0] C1AB5;
wire A1AB5;
wire signed [6:0] C1AC5;
wire A1AC5;
wire signed [6:0] C1AD5;
wire A1AD5;
wire signed [6:0] C1B05;
wire A1B05;
wire signed [6:0] C1B15;
wire A1B15;
wire signed [6:0] C1B25;
wire A1B25;
wire signed [6:0] C1B35;
wire A1B35;
wire signed [6:0] C1B45;
wire A1B45;
wire signed [6:0] C1B55;
wire A1B55;
wire signed [6:0] C1B65;
wire A1B65;
wire signed [6:0] C1B75;
wire A1B75;
wire signed [6:0] C1B85;
wire A1B85;
wire signed [6:0] C1B95;
wire A1B95;
wire signed [6:0] C1BA5;
wire A1BA5;
wire signed [6:0] C1BB5;
wire A1BB5;
wire signed [6:0] C1BC5;
wire A1BC5;
wire signed [6:0] C1BD5;
wire A1BD5;
wire signed [6:0] C1C05;
wire A1C05;
wire signed [6:0] C1C15;
wire A1C15;
wire signed [6:0] C1C25;
wire A1C25;
wire signed [6:0] C1C35;
wire A1C35;
wire signed [6:0] C1C45;
wire A1C45;
wire signed [6:0] C1C55;
wire A1C55;
wire signed [6:0] C1C65;
wire A1C65;
wire signed [6:0] C1C75;
wire A1C75;
wire signed [6:0] C1C85;
wire A1C85;
wire signed [6:0] C1C95;
wire A1C95;
wire signed [6:0] C1CA5;
wire A1CA5;
wire signed [6:0] C1CB5;
wire A1CB5;
wire signed [6:0] C1CC5;
wire A1CC5;
wire signed [6:0] C1CD5;
wire A1CD5;
wire signed [6:0] C1D05;
wire A1D05;
wire signed [6:0] C1D15;
wire A1D15;
wire signed [6:0] C1D25;
wire A1D25;
wire signed [6:0] C1D35;
wire A1D35;
wire signed [6:0] C1D45;
wire A1D45;
wire signed [6:0] C1D55;
wire A1D55;
wire signed [6:0] C1D65;
wire A1D65;
wire signed [6:0] C1D75;
wire A1D75;
wire signed [6:0] C1D85;
wire A1D85;
wire signed [6:0] C1D95;
wire A1D95;
wire signed [6:0] C1DA5;
wire A1DA5;
wire signed [6:0] C1DB5;
wire A1DB5;
wire signed [6:0] C1DC5;
wire A1DC5;
wire signed [6:0] C1DD5;
wire A1DD5;
wire signed [6:0] C1006;
wire A1006;
wire signed [6:0] C1016;
wire A1016;
wire signed [6:0] C1026;
wire A1026;
wire signed [6:0] C1036;
wire A1036;
wire signed [6:0] C1046;
wire A1046;
wire signed [6:0] C1056;
wire A1056;
wire signed [6:0] C1066;
wire A1066;
wire signed [6:0] C1076;
wire A1076;
wire signed [6:0] C1086;
wire A1086;
wire signed [6:0] C1096;
wire A1096;
wire signed [6:0] C10A6;
wire A10A6;
wire signed [6:0] C10B6;
wire A10B6;
wire signed [6:0] C10C6;
wire A10C6;
wire signed [6:0] C10D6;
wire A10D6;
wire signed [6:0] C1106;
wire A1106;
wire signed [6:0] C1116;
wire A1116;
wire signed [6:0] C1126;
wire A1126;
wire signed [6:0] C1136;
wire A1136;
wire signed [6:0] C1146;
wire A1146;
wire signed [6:0] C1156;
wire A1156;
wire signed [6:0] C1166;
wire A1166;
wire signed [6:0] C1176;
wire A1176;
wire signed [6:0] C1186;
wire A1186;
wire signed [6:0] C1196;
wire A1196;
wire signed [6:0] C11A6;
wire A11A6;
wire signed [6:0] C11B6;
wire A11B6;
wire signed [6:0] C11C6;
wire A11C6;
wire signed [6:0] C11D6;
wire A11D6;
wire signed [6:0] C1206;
wire A1206;
wire signed [6:0] C1216;
wire A1216;
wire signed [6:0] C1226;
wire A1226;
wire signed [6:0] C1236;
wire A1236;
wire signed [6:0] C1246;
wire A1246;
wire signed [6:0] C1256;
wire A1256;
wire signed [6:0] C1266;
wire A1266;
wire signed [6:0] C1276;
wire A1276;
wire signed [6:0] C1286;
wire A1286;
wire signed [6:0] C1296;
wire A1296;
wire signed [6:0] C12A6;
wire A12A6;
wire signed [6:0] C12B6;
wire A12B6;
wire signed [6:0] C12C6;
wire A12C6;
wire signed [6:0] C12D6;
wire A12D6;
wire signed [6:0] C1306;
wire A1306;
wire signed [6:0] C1316;
wire A1316;
wire signed [6:0] C1326;
wire A1326;
wire signed [6:0] C1336;
wire A1336;
wire signed [6:0] C1346;
wire A1346;
wire signed [6:0] C1356;
wire A1356;
wire signed [6:0] C1366;
wire A1366;
wire signed [6:0] C1376;
wire A1376;
wire signed [6:0] C1386;
wire A1386;
wire signed [6:0] C1396;
wire A1396;
wire signed [6:0] C13A6;
wire A13A6;
wire signed [6:0] C13B6;
wire A13B6;
wire signed [6:0] C13C6;
wire A13C6;
wire signed [6:0] C13D6;
wire A13D6;
wire signed [6:0] C1406;
wire A1406;
wire signed [6:0] C1416;
wire A1416;
wire signed [6:0] C1426;
wire A1426;
wire signed [6:0] C1436;
wire A1436;
wire signed [6:0] C1446;
wire A1446;
wire signed [6:0] C1456;
wire A1456;
wire signed [6:0] C1466;
wire A1466;
wire signed [6:0] C1476;
wire A1476;
wire signed [6:0] C1486;
wire A1486;
wire signed [6:0] C1496;
wire A1496;
wire signed [6:0] C14A6;
wire A14A6;
wire signed [6:0] C14B6;
wire A14B6;
wire signed [6:0] C14C6;
wire A14C6;
wire signed [6:0] C14D6;
wire A14D6;
wire signed [6:0] C1506;
wire A1506;
wire signed [6:0] C1516;
wire A1516;
wire signed [6:0] C1526;
wire A1526;
wire signed [6:0] C1536;
wire A1536;
wire signed [6:0] C1546;
wire A1546;
wire signed [6:0] C1556;
wire A1556;
wire signed [6:0] C1566;
wire A1566;
wire signed [6:0] C1576;
wire A1576;
wire signed [6:0] C1586;
wire A1586;
wire signed [6:0] C1596;
wire A1596;
wire signed [6:0] C15A6;
wire A15A6;
wire signed [6:0] C15B6;
wire A15B6;
wire signed [6:0] C15C6;
wire A15C6;
wire signed [6:0] C15D6;
wire A15D6;
wire signed [6:0] C1606;
wire A1606;
wire signed [6:0] C1616;
wire A1616;
wire signed [6:0] C1626;
wire A1626;
wire signed [6:0] C1636;
wire A1636;
wire signed [6:0] C1646;
wire A1646;
wire signed [6:0] C1656;
wire A1656;
wire signed [6:0] C1666;
wire A1666;
wire signed [6:0] C1676;
wire A1676;
wire signed [6:0] C1686;
wire A1686;
wire signed [6:0] C1696;
wire A1696;
wire signed [6:0] C16A6;
wire A16A6;
wire signed [6:0] C16B6;
wire A16B6;
wire signed [6:0] C16C6;
wire A16C6;
wire signed [6:0] C16D6;
wire A16D6;
wire signed [6:0] C1706;
wire A1706;
wire signed [6:0] C1716;
wire A1716;
wire signed [6:0] C1726;
wire A1726;
wire signed [6:0] C1736;
wire A1736;
wire signed [6:0] C1746;
wire A1746;
wire signed [6:0] C1756;
wire A1756;
wire signed [6:0] C1766;
wire A1766;
wire signed [6:0] C1776;
wire A1776;
wire signed [6:0] C1786;
wire A1786;
wire signed [6:0] C1796;
wire A1796;
wire signed [6:0] C17A6;
wire A17A6;
wire signed [6:0] C17B6;
wire A17B6;
wire signed [6:0] C17C6;
wire A17C6;
wire signed [6:0] C17D6;
wire A17D6;
wire signed [6:0] C1806;
wire A1806;
wire signed [6:0] C1816;
wire A1816;
wire signed [6:0] C1826;
wire A1826;
wire signed [6:0] C1836;
wire A1836;
wire signed [6:0] C1846;
wire A1846;
wire signed [6:0] C1856;
wire A1856;
wire signed [6:0] C1866;
wire A1866;
wire signed [6:0] C1876;
wire A1876;
wire signed [6:0] C1886;
wire A1886;
wire signed [6:0] C1896;
wire A1896;
wire signed [6:0] C18A6;
wire A18A6;
wire signed [6:0] C18B6;
wire A18B6;
wire signed [6:0] C18C6;
wire A18C6;
wire signed [6:0] C18D6;
wire A18D6;
wire signed [6:0] C1906;
wire A1906;
wire signed [6:0] C1916;
wire A1916;
wire signed [6:0] C1926;
wire A1926;
wire signed [6:0] C1936;
wire A1936;
wire signed [6:0] C1946;
wire A1946;
wire signed [6:0] C1956;
wire A1956;
wire signed [6:0] C1966;
wire A1966;
wire signed [6:0] C1976;
wire A1976;
wire signed [6:0] C1986;
wire A1986;
wire signed [6:0] C1996;
wire A1996;
wire signed [6:0] C19A6;
wire A19A6;
wire signed [6:0] C19B6;
wire A19B6;
wire signed [6:0] C19C6;
wire A19C6;
wire signed [6:0] C19D6;
wire A19D6;
wire signed [6:0] C1A06;
wire A1A06;
wire signed [6:0] C1A16;
wire A1A16;
wire signed [6:0] C1A26;
wire A1A26;
wire signed [6:0] C1A36;
wire A1A36;
wire signed [6:0] C1A46;
wire A1A46;
wire signed [6:0] C1A56;
wire A1A56;
wire signed [6:0] C1A66;
wire A1A66;
wire signed [6:0] C1A76;
wire A1A76;
wire signed [6:0] C1A86;
wire A1A86;
wire signed [6:0] C1A96;
wire A1A96;
wire signed [6:0] C1AA6;
wire A1AA6;
wire signed [6:0] C1AB6;
wire A1AB6;
wire signed [6:0] C1AC6;
wire A1AC6;
wire signed [6:0] C1AD6;
wire A1AD6;
wire signed [6:0] C1B06;
wire A1B06;
wire signed [6:0] C1B16;
wire A1B16;
wire signed [6:0] C1B26;
wire A1B26;
wire signed [6:0] C1B36;
wire A1B36;
wire signed [6:0] C1B46;
wire A1B46;
wire signed [6:0] C1B56;
wire A1B56;
wire signed [6:0] C1B66;
wire A1B66;
wire signed [6:0] C1B76;
wire A1B76;
wire signed [6:0] C1B86;
wire A1B86;
wire signed [6:0] C1B96;
wire A1B96;
wire signed [6:0] C1BA6;
wire A1BA6;
wire signed [6:0] C1BB6;
wire A1BB6;
wire signed [6:0] C1BC6;
wire A1BC6;
wire signed [6:0] C1BD6;
wire A1BD6;
wire signed [6:0] C1C06;
wire A1C06;
wire signed [6:0] C1C16;
wire A1C16;
wire signed [6:0] C1C26;
wire A1C26;
wire signed [6:0] C1C36;
wire A1C36;
wire signed [6:0] C1C46;
wire A1C46;
wire signed [6:0] C1C56;
wire A1C56;
wire signed [6:0] C1C66;
wire A1C66;
wire signed [6:0] C1C76;
wire A1C76;
wire signed [6:0] C1C86;
wire A1C86;
wire signed [6:0] C1C96;
wire A1C96;
wire signed [6:0] C1CA6;
wire A1CA6;
wire signed [6:0] C1CB6;
wire A1CB6;
wire signed [6:0] C1CC6;
wire A1CC6;
wire signed [6:0] C1CD6;
wire A1CD6;
wire signed [6:0] C1D06;
wire A1D06;
wire signed [6:0] C1D16;
wire A1D16;
wire signed [6:0] C1D26;
wire A1D26;
wire signed [6:0] C1D36;
wire A1D36;
wire signed [6:0] C1D46;
wire A1D46;
wire signed [6:0] C1D56;
wire A1D56;
wire signed [6:0] C1D66;
wire A1D66;
wire signed [6:0] C1D76;
wire A1D76;
wire signed [6:0] C1D86;
wire A1D86;
wire signed [6:0] C1D96;
wire A1D96;
wire signed [6:0] C1DA6;
wire A1DA6;
wire signed [6:0] C1DB6;
wire A1DB6;
wire signed [6:0] C1DC6;
wire A1DC6;
wire signed [6:0] C1DD6;
wire A1DD6;
wire signed [6:0] C1007;
wire A1007;
wire signed [6:0] C1017;
wire A1017;
wire signed [6:0] C1027;
wire A1027;
wire signed [6:0] C1037;
wire A1037;
wire signed [6:0] C1047;
wire A1047;
wire signed [6:0] C1057;
wire A1057;
wire signed [6:0] C1067;
wire A1067;
wire signed [6:0] C1077;
wire A1077;
wire signed [6:0] C1087;
wire A1087;
wire signed [6:0] C1097;
wire A1097;
wire signed [6:0] C10A7;
wire A10A7;
wire signed [6:0] C10B7;
wire A10B7;
wire signed [6:0] C10C7;
wire A10C7;
wire signed [6:0] C10D7;
wire A10D7;
wire signed [6:0] C1107;
wire A1107;
wire signed [6:0] C1117;
wire A1117;
wire signed [6:0] C1127;
wire A1127;
wire signed [6:0] C1137;
wire A1137;
wire signed [6:0] C1147;
wire A1147;
wire signed [6:0] C1157;
wire A1157;
wire signed [6:0] C1167;
wire A1167;
wire signed [6:0] C1177;
wire A1177;
wire signed [6:0] C1187;
wire A1187;
wire signed [6:0] C1197;
wire A1197;
wire signed [6:0] C11A7;
wire A11A7;
wire signed [6:0] C11B7;
wire A11B7;
wire signed [6:0] C11C7;
wire A11C7;
wire signed [6:0] C11D7;
wire A11D7;
wire signed [6:0] C1207;
wire A1207;
wire signed [6:0] C1217;
wire A1217;
wire signed [6:0] C1227;
wire A1227;
wire signed [6:0] C1237;
wire A1237;
wire signed [6:0] C1247;
wire A1247;
wire signed [6:0] C1257;
wire A1257;
wire signed [6:0] C1267;
wire A1267;
wire signed [6:0] C1277;
wire A1277;
wire signed [6:0] C1287;
wire A1287;
wire signed [6:0] C1297;
wire A1297;
wire signed [6:0] C12A7;
wire A12A7;
wire signed [6:0] C12B7;
wire A12B7;
wire signed [6:0] C12C7;
wire A12C7;
wire signed [6:0] C12D7;
wire A12D7;
wire signed [6:0] C1307;
wire A1307;
wire signed [6:0] C1317;
wire A1317;
wire signed [6:0] C1327;
wire A1327;
wire signed [6:0] C1337;
wire A1337;
wire signed [6:0] C1347;
wire A1347;
wire signed [6:0] C1357;
wire A1357;
wire signed [6:0] C1367;
wire A1367;
wire signed [6:0] C1377;
wire A1377;
wire signed [6:0] C1387;
wire A1387;
wire signed [6:0] C1397;
wire A1397;
wire signed [6:0] C13A7;
wire A13A7;
wire signed [6:0] C13B7;
wire A13B7;
wire signed [6:0] C13C7;
wire A13C7;
wire signed [6:0] C13D7;
wire A13D7;
wire signed [6:0] C1407;
wire A1407;
wire signed [6:0] C1417;
wire A1417;
wire signed [6:0] C1427;
wire A1427;
wire signed [6:0] C1437;
wire A1437;
wire signed [6:0] C1447;
wire A1447;
wire signed [6:0] C1457;
wire A1457;
wire signed [6:0] C1467;
wire A1467;
wire signed [6:0] C1477;
wire A1477;
wire signed [6:0] C1487;
wire A1487;
wire signed [6:0] C1497;
wire A1497;
wire signed [6:0] C14A7;
wire A14A7;
wire signed [6:0] C14B7;
wire A14B7;
wire signed [6:0] C14C7;
wire A14C7;
wire signed [6:0] C14D7;
wire A14D7;
wire signed [6:0] C1507;
wire A1507;
wire signed [6:0] C1517;
wire A1517;
wire signed [6:0] C1527;
wire A1527;
wire signed [6:0] C1537;
wire A1537;
wire signed [6:0] C1547;
wire A1547;
wire signed [6:0] C1557;
wire A1557;
wire signed [6:0] C1567;
wire A1567;
wire signed [6:0] C1577;
wire A1577;
wire signed [6:0] C1587;
wire A1587;
wire signed [6:0] C1597;
wire A1597;
wire signed [6:0] C15A7;
wire A15A7;
wire signed [6:0] C15B7;
wire A15B7;
wire signed [6:0] C15C7;
wire A15C7;
wire signed [6:0] C15D7;
wire A15D7;
wire signed [6:0] C1607;
wire A1607;
wire signed [6:0] C1617;
wire A1617;
wire signed [6:0] C1627;
wire A1627;
wire signed [6:0] C1637;
wire A1637;
wire signed [6:0] C1647;
wire A1647;
wire signed [6:0] C1657;
wire A1657;
wire signed [6:0] C1667;
wire A1667;
wire signed [6:0] C1677;
wire A1677;
wire signed [6:0] C1687;
wire A1687;
wire signed [6:0] C1697;
wire A1697;
wire signed [6:0] C16A7;
wire A16A7;
wire signed [6:0] C16B7;
wire A16B7;
wire signed [6:0] C16C7;
wire A16C7;
wire signed [6:0] C16D7;
wire A16D7;
wire signed [6:0] C1707;
wire A1707;
wire signed [6:0] C1717;
wire A1717;
wire signed [6:0] C1727;
wire A1727;
wire signed [6:0] C1737;
wire A1737;
wire signed [6:0] C1747;
wire A1747;
wire signed [6:0] C1757;
wire A1757;
wire signed [6:0] C1767;
wire A1767;
wire signed [6:0] C1777;
wire A1777;
wire signed [6:0] C1787;
wire A1787;
wire signed [6:0] C1797;
wire A1797;
wire signed [6:0] C17A7;
wire A17A7;
wire signed [6:0] C17B7;
wire A17B7;
wire signed [6:0] C17C7;
wire A17C7;
wire signed [6:0] C17D7;
wire A17D7;
wire signed [6:0] C1807;
wire A1807;
wire signed [6:0] C1817;
wire A1817;
wire signed [6:0] C1827;
wire A1827;
wire signed [6:0] C1837;
wire A1837;
wire signed [6:0] C1847;
wire A1847;
wire signed [6:0] C1857;
wire A1857;
wire signed [6:0] C1867;
wire A1867;
wire signed [6:0] C1877;
wire A1877;
wire signed [6:0] C1887;
wire A1887;
wire signed [6:0] C1897;
wire A1897;
wire signed [6:0] C18A7;
wire A18A7;
wire signed [6:0] C18B7;
wire A18B7;
wire signed [6:0] C18C7;
wire A18C7;
wire signed [6:0] C18D7;
wire A18D7;
wire signed [6:0] C1907;
wire A1907;
wire signed [6:0] C1917;
wire A1917;
wire signed [6:0] C1927;
wire A1927;
wire signed [6:0] C1937;
wire A1937;
wire signed [6:0] C1947;
wire A1947;
wire signed [6:0] C1957;
wire A1957;
wire signed [6:0] C1967;
wire A1967;
wire signed [6:0] C1977;
wire A1977;
wire signed [6:0] C1987;
wire A1987;
wire signed [6:0] C1997;
wire A1997;
wire signed [6:0] C19A7;
wire A19A7;
wire signed [6:0] C19B7;
wire A19B7;
wire signed [6:0] C19C7;
wire A19C7;
wire signed [6:0] C19D7;
wire A19D7;
wire signed [6:0] C1A07;
wire A1A07;
wire signed [6:0] C1A17;
wire A1A17;
wire signed [6:0] C1A27;
wire A1A27;
wire signed [6:0] C1A37;
wire A1A37;
wire signed [6:0] C1A47;
wire A1A47;
wire signed [6:0] C1A57;
wire A1A57;
wire signed [6:0] C1A67;
wire A1A67;
wire signed [6:0] C1A77;
wire A1A77;
wire signed [6:0] C1A87;
wire A1A87;
wire signed [6:0] C1A97;
wire A1A97;
wire signed [6:0] C1AA7;
wire A1AA7;
wire signed [6:0] C1AB7;
wire A1AB7;
wire signed [6:0] C1AC7;
wire A1AC7;
wire signed [6:0] C1AD7;
wire A1AD7;
wire signed [6:0] C1B07;
wire A1B07;
wire signed [6:0] C1B17;
wire A1B17;
wire signed [6:0] C1B27;
wire A1B27;
wire signed [6:0] C1B37;
wire A1B37;
wire signed [6:0] C1B47;
wire A1B47;
wire signed [6:0] C1B57;
wire A1B57;
wire signed [6:0] C1B67;
wire A1B67;
wire signed [6:0] C1B77;
wire A1B77;
wire signed [6:0] C1B87;
wire A1B87;
wire signed [6:0] C1B97;
wire A1B97;
wire signed [6:0] C1BA7;
wire A1BA7;
wire signed [6:0] C1BB7;
wire A1BB7;
wire signed [6:0] C1BC7;
wire A1BC7;
wire signed [6:0] C1BD7;
wire A1BD7;
wire signed [6:0] C1C07;
wire A1C07;
wire signed [6:0] C1C17;
wire A1C17;
wire signed [6:0] C1C27;
wire A1C27;
wire signed [6:0] C1C37;
wire A1C37;
wire signed [6:0] C1C47;
wire A1C47;
wire signed [6:0] C1C57;
wire A1C57;
wire signed [6:0] C1C67;
wire A1C67;
wire signed [6:0] C1C77;
wire A1C77;
wire signed [6:0] C1C87;
wire A1C87;
wire signed [6:0] C1C97;
wire A1C97;
wire signed [6:0] C1CA7;
wire A1CA7;
wire signed [6:0] C1CB7;
wire A1CB7;
wire signed [6:0] C1CC7;
wire A1CC7;
wire signed [6:0] C1CD7;
wire A1CD7;
wire signed [6:0] C1D07;
wire A1D07;
wire signed [6:0] C1D17;
wire A1D17;
wire signed [6:0] C1D27;
wire A1D27;
wire signed [6:0] C1D37;
wire A1D37;
wire signed [6:0] C1D47;
wire A1D47;
wire signed [6:0] C1D57;
wire A1D57;
wire signed [6:0] C1D67;
wire A1D67;
wire signed [6:0] C1D77;
wire A1D77;
wire signed [6:0] C1D87;
wire A1D87;
wire signed [6:0] C1D97;
wire A1D97;
wire signed [6:0] C1DA7;
wire A1DA7;
wire signed [6:0] C1DB7;
wire A1DB7;
wire signed [6:0] C1DC7;
wire A1DC7;
wire signed [6:0] C1DD7;
wire A1DD7;
DFF_save_fm DFF_P0(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1000));
DFF_save_fm DFF_P1(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1010));
DFF_save_fm DFF_P2(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1020));
DFF_save_fm DFF_P3(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1030));
DFF_save_fm DFF_P4(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1040));
DFF_save_fm DFF_P5(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1050));
DFF_save_fm DFF_P6(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1060));
DFF_save_fm DFF_P7(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1070));
DFF_save_fm DFF_P8(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1080));
DFF_save_fm DFF_P9(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1090));
DFF_save_fm DFF_P10(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10A0));
DFF_save_fm DFF_P11(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10B0));
DFF_save_fm DFF_P12(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10C0));
DFF_save_fm DFF_P13(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10D0));
DFF_save_fm DFF_P14(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10E0));
DFF_save_fm DFF_P15(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10F0));
DFF_save_fm DFF_P16(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1100));
DFF_save_fm DFF_P17(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1110));
DFF_save_fm DFF_P18(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1120));
DFF_save_fm DFF_P19(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1130));
DFF_save_fm DFF_P20(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1140));
DFF_save_fm DFF_P21(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1150));
DFF_save_fm DFF_P22(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1160));
DFF_save_fm DFF_P23(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1170));
DFF_save_fm DFF_P24(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1180));
DFF_save_fm DFF_P25(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1190));
DFF_save_fm DFF_P26(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11A0));
DFF_save_fm DFF_P27(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11B0));
DFF_save_fm DFF_P28(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11C0));
DFF_save_fm DFF_P29(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11D0));
DFF_save_fm DFF_P30(.clk(clk),.rstn(rstn),.reset_value(0),.q(P11E0));
DFF_save_fm DFF_P31(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11F0));
DFF_save_fm DFF_P32(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1200));
DFF_save_fm DFF_P33(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1210));
DFF_save_fm DFF_P34(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1220));
DFF_save_fm DFF_P35(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1230));
DFF_save_fm DFF_P36(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1240));
DFF_save_fm DFF_P37(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1250));
DFF_save_fm DFF_P38(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1260));
DFF_save_fm DFF_P39(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1270));
DFF_save_fm DFF_P40(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1280));
DFF_save_fm DFF_P41(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1290));
DFF_save_fm DFF_P42(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12A0));
DFF_save_fm DFF_P43(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12B0));
DFF_save_fm DFF_P44(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12C0));
DFF_save_fm DFF_P45(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12D0));
DFF_save_fm DFF_P46(.clk(clk),.rstn(rstn),.reset_value(0),.q(P12E0));
DFF_save_fm DFF_P47(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12F0));
DFF_save_fm DFF_P48(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1300));
DFF_save_fm DFF_P49(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1310));
DFF_save_fm DFF_P50(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1320));
DFF_save_fm DFF_P51(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1330));
DFF_save_fm DFF_P52(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1340));
DFF_save_fm DFF_P53(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1350));
DFF_save_fm DFF_P54(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1360));
DFF_save_fm DFF_P55(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1370));
DFF_save_fm DFF_P56(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1380));
DFF_save_fm DFF_P57(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1390));
DFF_save_fm DFF_P58(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13A0));
DFF_save_fm DFF_P59(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13B0));
DFF_save_fm DFF_P60(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13C0));
DFF_save_fm DFF_P61(.clk(clk),.rstn(rstn),.reset_value(0),.q(P13D0));
DFF_save_fm DFF_P62(.clk(clk),.rstn(rstn),.reset_value(0),.q(P13E0));
DFF_save_fm DFF_P63(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13F0));
DFF_save_fm DFF_P64(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1400));
DFF_save_fm DFF_P65(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1410));
DFF_save_fm DFF_P66(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1420));
DFF_save_fm DFF_P67(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1430));
DFF_save_fm DFF_P68(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1440));
DFF_save_fm DFF_P69(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1450));
DFF_save_fm DFF_P70(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1460));
DFF_save_fm DFF_P71(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1470));
DFF_save_fm DFF_P72(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1480));
DFF_save_fm DFF_P73(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1490));
DFF_save_fm DFF_P74(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14A0));
DFF_save_fm DFF_P75(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14B0));
DFF_save_fm DFF_P76(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14C0));
DFF_save_fm DFF_P77(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14D0));
DFF_save_fm DFF_P78(.clk(clk),.rstn(rstn),.reset_value(0),.q(P14E0));
DFF_save_fm DFF_P79(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14F0));
DFF_save_fm DFF_P80(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1500));
DFF_save_fm DFF_P81(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1510));
DFF_save_fm DFF_P82(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1520));
DFF_save_fm DFF_P83(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1530));
DFF_save_fm DFF_P84(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1540));
DFF_save_fm DFF_P85(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1550));
DFF_save_fm DFF_P86(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1560));
DFF_save_fm DFF_P87(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1570));
DFF_save_fm DFF_P88(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1580));
DFF_save_fm DFF_P89(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1590));
DFF_save_fm DFF_P90(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15A0));
DFF_save_fm DFF_P91(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15B0));
DFF_save_fm DFF_P92(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15C0));
DFF_save_fm DFF_P93(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15D0));
DFF_save_fm DFF_P94(.clk(clk),.rstn(rstn),.reset_value(0),.q(P15E0));
DFF_save_fm DFF_P95(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15F0));
DFF_save_fm DFF_P96(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1600));
DFF_save_fm DFF_P97(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1610));
DFF_save_fm DFF_P98(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1620));
DFF_save_fm DFF_P99(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1630));
DFF_save_fm DFF_P100(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1640));
DFF_save_fm DFF_P101(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1650));
DFF_save_fm DFF_P102(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1660));
DFF_save_fm DFF_P103(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1670));
DFF_save_fm DFF_P104(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1680));
DFF_save_fm DFF_P105(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1690));
DFF_save_fm DFF_P106(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16A0));
DFF_save_fm DFF_P107(.clk(clk),.rstn(rstn),.reset_value(0),.q(P16B0));
DFF_save_fm DFF_P108(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16C0));
DFF_save_fm DFF_P109(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16D0));
DFF_save_fm DFF_P110(.clk(clk),.rstn(rstn),.reset_value(0),.q(P16E0));
DFF_save_fm DFF_P111(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16F0));
DFF_save_fm DFF_P112(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1700));
DFF_save_fm DFF_P113(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1710));
DFF_save_fm DFF_P114(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1720));
DFF_save_fm DFF_P115(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1730));
DFF_save_fm DFF_P116(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1740));
DFF_save_fm DFF_P117(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1750));
DFF_save_fm DFF_P118(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1760));
DFF_save_fm DFF_P119(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1770));
DFF_save_fm DFF_P120(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1780));
DFF_save_fm DFF_P121(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1790));
DFF_save_fm DFF_P122(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17A0));
DFF_save_fm DFF_P123(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17B0));
DFF_save_fm DFF_P124(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17C0));
DFF_save_fm DFF_P125(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17D0));
DFF_save_fm DFF_P126(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17E0));
DFF_save_fm DFF_P127(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17F0));
DFF_save_fm DFF_P128(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1800));
DFF_save_fm DFF_P129(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1810));
DFF_save_fm DFF_P130(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1820));
DFF_save_fm DFF_P131(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1830));
DFF_save_fm DFF_P132(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1840));
DFF_save_fm DFF_P133(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1850));
DFF_save_fm DFF_P134(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1860));
DFF_save_fm DFF_P135(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1870));
DFF_save_fm DFF_P136(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1880));
DFF_save_fm DFF_P137(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1890));
DFF_save_fm DFF_P138(.clk(clk),.rstn(rstn),.reset_value(0),.q(P18A0));
DFF_save_fm DFF_P139(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18B0));
DFF_save_fm DFF_P140(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18C0));
DFF_save_fm DFF_P141(.clk(clk),.rstn(rstn),.reset_value(0),.q(P18D0));
DFF_save_fm DFF_P142(.clk(clk),.rstn(rstn),.reset_value(0),.q(P18E0));
DFF_save_fm DFF_P143(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18F0));
DFF_save_fm DFF_P144(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1900));
DFF_save_fm DFF_P145(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1910));
DFF_save_fm DFF_P146(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1920));
DFF_save_fm DFF_P147(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1930));
DFF_save_fm DFF_P148(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1940));
DFF_save_fm DFF_P149(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1950));
DFF_save_fm DFF_P150(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1960));
DFF_save_fm DFF_P151(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1970));
DFF_save_fm DFF_P152(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1980));
DFF_save_fm DFF_P153(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1990));
DFF_save_fm DFF_P154(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19A0));
DFF_save_fm DFF_P155(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19B0));
DFF_save_fm DFF_P156(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19C0));
DFF_save_fm DFF_P157(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19D0));
DFF_save_fm DFF_P158(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19E0));
DFF_save_fm DFF_P159(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19F0));
DFF_save_fm DFF_P160(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A00));
DFF_save_fm DFF_P161(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A10));
DFF_save_fm DFF_P162(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A20));
DFF_save_fm DFF_P163(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A30));
DFF_save_fm DFF_P164(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A40));
DFF_save_fm DFF_P165(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A50));
DFF_save_fm DFF_P166(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A60));
DFF_save_fm DFF_P167(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A70));
DFF_save_fm DFF_P168(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A80));
DFF_save_fm DFF_P169(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A90));
DFF_save_fm DFF_P170(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AA0));
DFF_save_fm DFF_P171(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AB0));
DFF_save_fm DFF_P172(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AC0));
DFF_save_fm DFF_P173(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AD0));
DFF_save_fm DFF_P174(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AE0));
DFF_save_fm DFF_P175(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AF0));
DFF_save_fm DFF_P176(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B00));
DFF_save_fm DFF_P177(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B10));
DFF_save_fm DFF_P178(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B20));
DFF_save_fm DFF_P179(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B30));
DFF_save_fm DFF_P180(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B40));
DFF_save_fm DFF_P181(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B50));
DFF_save_fm DFF_P182(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B60));
DFF_save_fm DFF_P183(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B70));
DFF_save_fm DFF_P184(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B80));
DFF_save_fm DFF_P185(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B90));
DFF_save_fm DFF_P186(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BA0));
DFF_save_fm DFF_P187(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BB0));
DFF_save_fm DFF_P188(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BC0));
DFF_save_fm DFF_P189(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BD0));
DFF_save_fm DFF_P190(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BE0));
DFF_save_fm DFF_P191(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BF0));
DFF_save_fm DFF_P192(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C00));
DFF_save_fm DFF_P193(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C10));
DFF_save_fm DFF_P194(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C20));
DFF_save_fm DFF_P195(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C30));
DFF_save_fm DFF_P196(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C40));
DFF_save_fm DFF_P197(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C50));
DFF_save_fm DFF_P198(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C60));
DFF_save_fm DFF_P199(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C70));
DFF_save_fm DFF_P200(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C80));
DFF_save_fm DFF_P201(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C90));
DFF_save_fm DFF_P202(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CA0));
DFF_save_fm DFF_P203(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CB0));
DFF_save_fm DFF_P204(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CC0));
DFF_save_fm DFF_P205(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CD0));
DFF_save_fm DFF_P206(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CE0));
DFF_save_fm DFF_P207(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CF0));
DFF_save_fm DFF_P208(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D00));
DFF_save_fm DFF_P209(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D10));
DFF_save_fm DFF_P210(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D20));
DFF_save_fm DFF_P211(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D30));
DFF_save_fm DFF_P212(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D40));
DFF_save_fm DFF_P213(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D50));
DFF_save_fm DFF_P214(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D60));
DFF_save_fm DFF_P215(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D70));
DFF_save_fm DFF_P216(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D80));
DFF_save_fm DFF_P217(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D90));
DFF_save_fm DFF_P218(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DA0));
DFF_save_fm DFF_P219(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DB0));
DFF_save_fm DFF_P220(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1DC0));
DFF_save_fm DFF_P221(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1DD0));
DFF_save_fm DFF_P222(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1DE0));
DFF_save_fm DFF_P223(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DF0));
DFF_save_fm DFF_P224(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E00));
DFF_save_fm DFF_P225(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E10));
DFF_save_fm DFF_P226(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E20));
DFF_save_fm DFF_P227(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E30));
DFF_save_fm DFF_P228(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E40));
DFF_save_fm DFF_P229(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E50));
DFF_save_fm DFF_P230(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E60));
DFF_save_fm DFF_P231(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E70));
DFF_save_fm DFF_P232(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E80));
DFF_save_fm DFF_P233(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E90));
DFF_save_fm DFF_P234(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EA0));
DFF_save_fm DFF_P235(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EB0));
DFF_save_fm DFF_P236(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EC0));
DFF_save_fm DFF_P237(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1ED0));
DFF_save_fm DFF_P238(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1EE0));
DFF_save_fm DFF_P239(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EF0));
DFF_save_fm DFF_P240(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F00));
DFF_save_fm DFF_P241(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F10));
DFF_save_fm DFF_P242(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F20));
DFF_save_fm DFF_P243(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F30));
DFF_save_fm DFF_P244(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F40));
DFF_save_fm DFF_P245(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F50));
DFF_save_fm DFF_P246(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F60));
DFF_save_fm DFF_P247(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F70));
DFF_save_fm DFF_P248(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F80));
DFF_save_fm DFF_P249(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F90));
DFF_save_fm DFF_P250(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FA0));
DFF_save_fm DFF_P251(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FB0));
DFF_save_fm DFF_P252(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FC0));
DFF_save_fm DFF_P253(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FD0));
DFF_save_fm DFF_P254(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FE0));
DFF_save_fm DFF_P255(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FF0));
DFF_save_fm DFF_P256(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1001));
DFF_save_fm DFF_P257(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1011));
DFF_save_fm DFF_P258(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1021));
DFF_save_fm DFF_P259(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1031));
DFF_save_fm DFF_P260(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1041));
DFF_save_fm DFF_P261(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1051));
DFF_save_fm DFF_P262(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1061));
DFF_save_fm DFF_P263(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1071));
DFF_save_fm DFF_P264(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1081));
DFF_save_fm DFF_P265(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1091));
DFF_save_fm DFF_P266(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10A1));
DFF_save_fm DFF_P267(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10B1));
DFF_save_fm DFF_P268(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10C1));
DFF_save_fm DFF_P269(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10D1));
DFF_save_fm DFF_P270(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10E1));
DFF_save_fm DFF_P271(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10F1));
DFF_save_fm DFF_P272(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1101));
DFF_save_fm DFF_P273(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1111));
DFF_save_fm DFF_P274(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1121));
DFF_save_fm DFF_P275(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1131));
DFF_save_fm DFF_P276(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1141));
DFF_save_fm DFF_P277(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1151));
DFF_save_fm DFF_P278(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1161));
DFF_save_fm DFF_P279(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1171));
DFF_save_fm DFF_P280(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1181));
DFF_save_fm DFF_P281(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1191));
DFF_save_fm DFF_P282(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11A1));
DFF_save_fm DFF_P283(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11B1));
DFF_save_fm DFF_P284(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11C1));
DFF_save_fm DFF_P285(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11D1));
DFF_save_fm DFF_P286(.clk(clk),.rstn(rstn),.reset_value(0),.q(P11E1));
DFF_save_fm DFF_P287(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11F1));
DFF_save_fm DFF_P288(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1201));
DFF_save_fm DFF_P289(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1211));
DFF_save_fm DFF_P290(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1221));
DFF_save_fm DFF_P291(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1231));
DFF_save_fm DFF_P292(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1241));
DFF_save_fm DFF_P293(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1251));
DFF_save_fm DFF_P294(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1261));
DFF_save_fm DFF_P295(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1271));
DFF_save_fm DFF_P296(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1281));
DFF_save_fm DFF_P297(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1291));
DFF_save_fm DFF_P298(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12A1));
DFF_save_fm DFF_P299(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12B1));
DFF_save_fm DFF_P300(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12C1));
DFF_save_fm DFF_P301(.clk(clk),.rstn(rstn),.reset_value(0),.q(P12D1));
DFF_save_fm DFF_P302(.clk(clk),.rstn(rstn),.reset_value(0),.q(P12E1));
DFF_save_fm DFF_P303(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12F1));
DFF_save_fm DFF_P304(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1301));
DFF_save_fm DFF_P305(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1311));
DFF_save_fm DFF_P306(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1321));
DFF_save_fm DFF_P307(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1331));
DFF_save_fm DFF_P308(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1341));
DFF_save_fm DFF_P309(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1351));
DFF_save_fm DFF_P310(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1361));
DFF_save_fm DFF_P311(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1371));
DFF_save_fm DFF_P312(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1381));
DFF_save_fm DFF_P313(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1391));
DFF_save_fm DFF_P314(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13A1));
DFF_save_fm DFF_P315(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13B1));
DFF_save_fm DFF_P316(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13C1));
DFF_save_fm DFF_P317(.clk(clk),.rstn(rstn),.reset_value(0),.q(P13D1));
DFF_save_fm DFF_P318(.clk(clk),.rstn(rstn),.reset_value(0),.q(P13E1));
DFF_save_fm DFF_P319(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13F1));
DFF_save_fm DFF_P320(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1401));
DFF_save_fm DFF_P321(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1411));
DFF_save_fm DFF_P322(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1421));
DFF_save_fm DFF_P323(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1431));
DFF_save_fm DFF_P324(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1441));
DFF_save_fm DFF_P325(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1451));
DFF_save_fm DFF_P326(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1461));
DFF_save_fm DFF_P327(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1471));
DFF_save_fm DFF_P328(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1481));
DFF_save_fm DFF_P329(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1491));
DFF_save_fm DFF_P330(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14A1));
DFF_save_fm DFF_P331(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14B1));
DFF_save_fm DFF_P332(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14C1));
DFF_save_fm DFF_P333(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14D1));
DFF_save_fm DFF_P334(.clk(clk),.rstn(rstn),.reset_value(0),.q(P14E1));
DFF_save_fm DFF_P335(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14F1));
DFF_save_fm DFF_P336(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1501));
DFF_save_fm DFF_P337(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1511));
DFF_save_fm DFF_P338(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1521));
DFF_save_fm DFF_P339(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1531));
DFF_save_fm DFF_P340(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1541));
DFF_save_fm DFF_P341(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1551));
DFF_save_fm DFF_P342(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1561));
DFF_save_fm DFF_P343(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1571));
DFF_save_fm DFF_P344(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1581));
DFF_save_fm DFF_P345(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1591));
DFF_save_fm DFF_P346(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15A1));
DFF_save_fm DFF_P347(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15B1));
DFF_save_fm DFF_P348(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15C1));
DFF_save_fm DFF_P349(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15D1));
DFF_save_fm DFF_P350(.clk(clk),.rstn(rstn),.reset_value(0),.q(P15E1));
DFF_save_fm DFF_P351(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15F1));
DFF_save_fm DFF_P352(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1601));
DFF_save_fm DFF_P353(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1611));
DFF_save_fm DFF_P354(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1621));
DFF_save_fm DFF_P355(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1631));
DFF_save_fm DFF_P356(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1641));
DFF_save_fm DFF_P357(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1651));
DFF_save_fm DFF_P358(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1661));
DFF_save_fm DFF_P359(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1671));
DFF_save_fm DFF_P360(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1681));
DFF_save_fm DFF_P361(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1691));
DFF_save_fm DFF_P362(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16A1));
DFF_save_fm DFF_P363(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16B1));
DFF_save_fm DFF_P364(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16C1));
DFF_save_fm DFF_P365(.clk(clk),.rstn(rstn),.reset_value(0),.q(P16D1));
DFF_save_fm DFF_P366(.clk(clk),.rstn(rstn),.reset_value(0),.q(P16E1));
DFF_save_fm DFF_P367(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16F1));
DFF_save_fm DFF_P368(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1701));
DFF_save_fm DFF_P369(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1711));
DFF_save_fm DFF_P370(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1721));
DFF_save_fm DFF_P371(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1731));
DFF_save_fm DFF_P372(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1741));
DFF_save_fm DFF_P373(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1751));
DFF_save_fm DFF_P374(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1761));
DFF_save_fm DFF_P375(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1771));
DFF_save_fm DFF_P376(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1781));
DFF_save_fm DFF_P377(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1791));
DFF_save_fm DFF_P378(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17A1));
DFF_save_fm DFF_P379(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17B1));
DFF_save_fm DFF_P380(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17C1));
DFF_save_fm DFF_P381(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17D1));
DFF_save_fm DFF_P382(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17E1));
DFF_save_fm DFF_P383(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17F1));
DFF_save_fm DFF_P384(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1801));
DFF_save_fm DFF_P385(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1811));
DFF_save_fm DFF_P386(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1821));
DFF_save_fm DFF_P387(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1831));
DFF_save_fm DFF_P388(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1841));
DFF_save_fm DFF_P389(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1851));
DFF_save_fm DFF_P390(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1861));
DFF_save_fm DFF_P391(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1871));
DFF_save_fm DFF_P392(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1881));
DFF_save_fm DFF_P393(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1891));
DFF_save_fm DFF_P394(.clk(clk),.rstn(rstn),.reset_value(0),.q(P18A1));
DFF_save_fm DFF_P395(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18B1));
DFF_save_fm DFF_P396(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18C1));
DFF_save_fm DFF_P397(.clk(clk),.rstn(rstn),.reset_value(0),.q(P18D1));
DFF_save_fm DFF_P398(.clk(clk),.rstn(rstn),.reset_value(0),.q(P18E1));
DFF_save_fm DFF_P399(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18F1));
DFF_save_fm DFF_P400(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1901));
DFF_save_fm DFF_P401(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1911));
DFF_save_fm DFF_P402(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1921));
DFF_save_fm DFF_P403(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1931));
DFF_save_fm DFF_P404(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1941));
DFF_save_fm DFF_P405(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1951));
DFF_save_fm DFF_P406(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1961));
DFF_save_fm DFF_P407(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1971));
DFF_save_fm DFF_P408(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1981));
DFF_save_fm DFF_P409(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1991));
DFF_save_fm DFF_P410(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19A1));
DFF_save_fm DFF_P411(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19B1));
DFF_save_fm DFF_P412(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19C1));
DFF_save_fm DFF_P413(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19D1));
DFF_save_fm DFF_P414(.clk(clk),.rstn(rstn),.reset_value(0),.q(P19E1));
DFF_save_fm DFF_P415(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19F1));
DFF_save_fm DFF_P416(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A01));
DFF_save_fm DFF_P417(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A11));
DFF_save_fm DFF_P418(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A21));
DFF_save_fm DFF_P419(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A31));
DFF_save_fm DFF_P420(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A41));
DFF_save_fm DFF_P421(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A51));
DFF_save_fm DFF_P422(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A61));
DFF_save_fm DFF_P423(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A71));
DFF_save_fm DFF_P424(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A81));
DFF_save_fm DFF_P425(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1A91));
DFF_save_fm DFF_P426(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AA1));
DFF_save_fm DFF_P427(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AB1));
DFF_save_fm DFF_P428(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AC1));
DFF_save_fm DFF_P429(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AD1));
DFF_save_fm DFF_P430(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1AE1));
DFF_save_fm DFF_P431(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AF1));
DFF_save_fm DFF_P432(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B01));
DFF_save_fm DFF_P433(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B11));
DFF_save_fm DFF_P434(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B21));
DFF_save_fm DFF_P435(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B31));
DFF_save_fm DFF_P436(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B41));
DFF_save_fm DFF_P437(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B51));
DFF_save_fm DFF_P438(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B61));
DFF_save_fm DFF_P439(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B71));
DFF_save_fm DFF_P440(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1B81));
DFF_save_fm DFF_P441(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B91));
DFF_save_fm DFF_P442(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BA1));
DFF_save_fm DFF_P443(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BB1));
DFF_save_fm DFF_P444(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BC1));
DFF_save_fm DFF_P445(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BD1));
DFF_save_fm DFF_P446(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1BE1));
DFF_save_fm DFF_P447(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BF1));
DFF_save_fm DFF_P448(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C01));
DFF_save_fm DFF_P449(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C11));
DFF_save_fm DFF_P450(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C21));
DFF_save_fm DFF_P451(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C31));
DFF_save_fm DFF_P452(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C41));
DFF_save_fm DFF_P453(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C51));
DFF_save_fm DFF_P454(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C61));
DFF_save_fm DFF_P455(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1C71));
DFF_save_fm DFF_P456(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C81));
DFF_save_fm DFF_P457(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C91));
DFF_save_fm DFF_P458(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CA1));
DFF_save_fm DFF_P459(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CB1));
DFF_save_fm DFF_P460(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CC1));
DFF_save_fm DFF_P461(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CD1));
DFF_save_fm DFF_P462(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CE1));
DFF_save_fm DFF_P463(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CF1));
DFF_save_fm DFF_P464(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D01));
DFF_save_fm DFF_P465(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D11));
DFF_save_fm DFF_P466(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D21));
DFF_save_fm DFF_P467(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D31));
DFF_save_fm DFF_P468(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D41));
DFF_save_fm DFF_P469(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D51));
DFF_save_fm DFF_P470(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D61));
DFF_save_fm DFF_P471(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D71));
DFF_save_fm DFF_P472(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D81));
DFF_save_fm DFF_P473(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D91));
DFF_save_fm DFF_P474(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DA1));
DFF_save_fm DFF_P475(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DB1));
DFF_save_fm DFF_P476(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1DC1));
DFF_save_fm DFF_P477(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1DD1));
DFF_save_fm DFF_P478(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1DE1));
DFF_save_fm DFF_P479(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DF1));
DFF_save_fm DFF_P480(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E01));
DFF_save_fm DFF_P481(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E11));
DFF_save_fm DFF_P482(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E21));
DFF_save_fm DFF_P483(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E31));
DFF_save_fm DFF_P484(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E41));
DFF_save_fm DFF_P485(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E51));
DFF_save_fm DFF_P486(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E61));
DFF_save_fm DFF_P487(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E71));
DFF_save_fm DFF_P488(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E81));
DFF_save_fm DFF_P489(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E91));
DFF_save_fm DFF_P490(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EA1));
DFF_save_fm DFF_P491(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EB1));
DFF_save_fm DFF_P492(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EC1));
DFF_save_fm DFF_P493(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1ED1));
DFF_save_fm DFF_P494(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1EE1));
DFF_save_fm DFF_P495(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EF1));
DFF_save_fm DFF_P496(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F01));
DFF_save_fm DFF_P497(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F11));
DFF_save_fm DFF_P498(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F21));
DFF_save_fm DFF_P499(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F31));
DFF_save_fm DFF_P500(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F41));
DFF_save_fm DFF_P501(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F51));
DFF_save_fm DFF_P502(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F61));
DFF_save_fm DFF_P503(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F71));
DFF_save_fm DFF_P504(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F81));
DFF_save_fm DFF_P505(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F91));
DFF_save_fm DFF_P506(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FA1));
DFF_save_fm DFF_P507(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FB1));
DFF_save_fm DFF_P508(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FC1));
DFF_save_fm DFF_P509(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FD1));
DFF_save_fm DFF_P510(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FE1));
DFF_save_fm DFF_P511(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FF1));
DFF_save_fm DFF_P512(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1002));
DFF_save_fm DFF_P513(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1012));
DFF_save_fm DFF_P514(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1022));
DFF_save_fm DFF_P515(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1032));
DFF_save_fm DFF_P516(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1042));
DFF_save_fm DFF_P517(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1052));
DFF_save_fm DFF_P518(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1062));
DFF_save_fm DFF_P519(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1072));
DFF_save_fm DFF_P520(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1082));
DFF_save_fm DFF_P521(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1092));
DFF_save_fm DFF_P522(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10A2));
DFF_save_fm DFF_P523(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10B2));
DFF_save_fm DFF_P524(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10C2));
DFF_save_fm DFF_P525(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10D2));
DFF_save_fm DFF_P526(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10E2));
DFF_save_fm DFF_P527(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10F2));
DFF_save_fm DFF_P528(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1102));
DFF_save_fm DFF_P529(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1112));
DFF_save_fm DFF_P530(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1122));
DFF_save_fm DFF_P531(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1132));
DFF_save_fm DFF_P532(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1142));
DFF_save_fm DFF_P533(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1152));
DFF_save_fm DFF_P534(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1162));
DFF_save_fm DFF_P535(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1172));
DFF_save_fm DFF_P536(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1182));
DFF_save_fm DFF_P537(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1192));
DFF_save_fm DFF_P538(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11A2));
DFF_save_fm DFF_P539(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11B2));
DFF_save_fm DFF_P540(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11C2));
DFF_save_fm DFF_P541(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11D2));
DFF_save_fm DFF_P542(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11E2));
DFF_save_fm DFF_P543(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11F2));
DFF_save_fm DFF_P544(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1202));
DFF_save_fm DFF_P545(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1212));
DFF_save_fm DFF_P546(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1222));
DFF_save_fm DFF_P547(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1232));
DFF_save_fm DFF_P548(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1242));
DFF_save_fm DFF_P549(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1252));
DFF_save_fm DFF_P550(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1262));
DFF_save_fm DFF_P551(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1272));
DFF_save_fm DFF_P552(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1282));
DFF_save_fm DFF_P553(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1292));
DFF_save_fm DFF_P554(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12A2));
DFF_save_fm DFF_P555(.clk(clk),.rstn(rstn),.reset_value(0),.q(P12B2));
DFF_save_fm DFF_P556(.clk(clk),.rstn(rstn),.reset_value(0),.q(P12C2));
DFF_save_fm DFF_P557(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12D2));
DFF_save_fm DFF_P558(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12E2));
DFF_save_fm DFF_P559(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12F2));
DFF_save_fm DFF_P560(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1302));
DFF_save_fm DFF_P561(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1312));
DFF_save_fm DFF_P562(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1322));
DFF_save_fm DFF_P563(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1332));
DFF_save_fm DFF_P564(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1342));
DFF_save_fm DFF_P565(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1352));
DFF_save_fm DFF_P566(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1362));
DFF_save_fm DFF_P567(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1372));
DFF_save_fm DFF_P568(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1382));
DFF_save_fm DFF_P569(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1392));
DFF_save_fm DFF_P570(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13A2));
DFF_save_fm DFF_P571(.clk(clk),.rstn(rstn),.reset_value(0),.q(P13B2));
DFF_save_fm DFF_P572(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13C2));
DFF_save_fm DFF_P573(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13D2));
DFF_save_fm DFF_P574(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13E2));
DFF_save_fm DFF_P575(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13F2));
DFF_save_fm DFF_P576(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1402));
DFF_save_fm DFF_P577(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1412));
DFF_save_fm DFF_P578(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1422));
DFF_save_fm DFF_P579(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1432));
DFF_save_fm DFF_P580(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1442));
DFF_save_fm DFF_P581(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1452));
DFF_save_fm DFF_P582(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1462));
DFF_save_fm DFF_P583(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1472));
DFF_save_fm DFF_P584(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1482));
DFF_save_fm DFF_P585(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1492));
DFF_save_fm DFF_P586(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14A2));
DFF_save_fm DFF_P587(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14B2));
DFF_save_fm DFF_P588(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14C2));
DFF_save_fm DFF_P589(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14D2));
DFF_save_fm DFF_P590(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14E2));
DFF_save_fm DFF_P591(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14F2));
DFF_save_fm DFF_P592(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1502));
DFF_save_fm DFF_P593(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1512));
DFF_save_fm DFF_P594(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1522));
DFF_save_fm DFF_P595(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1532));
DFF_save_fm DFF_P596(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1542));
DFF_save_fm DFF_P597(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1552));
DFF_save_fm DFF_P598(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1562));
DFF_save_fm DFF_P599(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1572));
DFF_save_fm DFF_P600(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1582));
DFF_save_fm DFF_P601(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1592));
DFF_save_fm DFF_P602(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15A2));
DFF_save_fm DFF_P603(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15B2));
DFF_save_fm DFF_P604(.clk(clk),.rstn(rstn),.reset_value(0),.q(P15C2));
DFF_save_fm DFF_P605(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15D2));
DFF_save_fm DFF_P606(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15E2));
DFF_save_fm DFF_P607(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15F2));
DFF_save_fm DFF_P608(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1602));
DFF_save_fm DFF_P609(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1612));
DFF_save_fm DFF_P610(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1622));
DFF_save_fm DFF_P611(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1632));
DFF_save_fm DFF_P612(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1642));
DFF_save_fm DFF_P613(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1652));
DFF_save_fm DFF_P614(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1662));
DFF_save_fm DFF_P615(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1672));
DFF_save_fm DFF_P616(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1682));
DFF_save_fm DFF_P617(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1692));
DFF_save_fm DFF_P618(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16A2));
DFF_save_fm DFF_P619(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16B2));
DFF_save_fm DFF_P620(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16C2));
DFF_save_fm DFF_P621(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16D2));
DFF_save_fm DFF_P622(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16E2));
DFF_save_fm DFF_P623(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16F2));
DFF_save_fm DFF_P624(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1702));
DFF_save_fm DFF_P625(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1712));
DFF_save_fm DFF_P626(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1722));
DFF_save_fm DFF_P627(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1732));
DFF_save_fm DFF_P628(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1742));
DFF_save_fm DFF_P629(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1752));
DFF_save_fm DFF_P630(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1762));
DFF_save_fm DFF_P631(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1772));
DFF_save_fm DFF_P632(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1782));
DFF_save_fm DFF_P633(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1792));
DFF_save_fm DFF_P634(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17A2));
DFF_save_fm DFF_P635(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17B2));
DFF_save_fm DFF_P636(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17C2));
DFF_save_fm DFF_P637(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17D2));
DFF_save_fm DFF_P638(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17E2));
DFF_save_fm DFF_P639(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17F2));
DFF_save_fm DFF_P640(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1802));
DFF_save_fm DFF_P641(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1812));
DFF_save_fm DFF_P642(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1822));
DFF_save_fm DFF_P643(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1832));
DFF_save_fm DFF_P644(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1842));
DFF_save_fm DFF_P645(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1852));
DFF_save_fm DFF_P646(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1862));
DFF_save_fm DFF_P647(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1872));
DFF_save_fm DFF_P648(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1882));
DFF_save_fm DFF_P649(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1892));
DFF_save_fm DFF_P650(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18A2));
DFF_save_fm DFF_P651(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18B2));
DFF_save_fm DFF_P652(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18C2));
DFF_save_fm DFF_P653(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18D2));
DFF_save_fm DFF_P654(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18E2));
DFF_save_fm DFF_P655(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18F2));
DFF_save_fm DFF_P656(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1902));
DFF_save_fm DFF_P657(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1912));
DFF_save_fm DFF_P658(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1922));
DFF_save_fm DFF_P659(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1932));
DFF_save_fm DFF_P660(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1942));
DFF_save_fm DFF_P661(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1952));
DFF_save_fm DFF_P662(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1962));
DFF_save_fm DFF_P663(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1972));
DFF_save_fm DFF_P664(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1982));
DFF_save_fm DFF_P665(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1992));
DFF_save_fm DFF_P666(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19A2));
DFF_save_fm DFF_P667(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19B2));
DFF_save_fm DFF_P668(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19C2));
DFF_save_fm DFF_P669(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19D2));
DFF_save_fm DFF_P670(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19E2));
DFF_save_fm DFF_P671(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19F2));
DFF_save_fm DFF_P672(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A02));
DFF_save_fm DFF_P673(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A12));
DFF_save_fm DFF_P674(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A22));
DFF_save_fm DFF_P675(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A32));
DFF_save_fm DFF_P676(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A42));
DFF_save_fm DFF_P677(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A52));
DFF_save_fm DFF_P678(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A62));
DFF_save_fm DFF_P679(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A72));
DFF_save_fm DFF_P680(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A82));
DFF_save_fm DFF_P681(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A92));
DFF_save_fm DFF_P682(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AA2));
DFF_save_fm DFF_P683(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AB2));
DFF_save_fm DFF_P684(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AC2));
DFF_save_fm DFF_P685(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AD2));
DFF_save_fm DFF_P686(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AE2));
DFF_save_fm DFF_P687(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AF2));
DFF_save_fm DFF_P688(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B02));
DFF_save_fm DFF_P689(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B12));
DFF_save_fm DFF_P690(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B22));
DFF_save_fm DFF_P691(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B32));
DFF_save_fm DFF_P692(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B42));
DFF_save_fm DFF_P693(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B52));
DFF_save_fm DFF_P694(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B62));
DFF_save_fm DFF_P695(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B72));
DFF_save_fm DFF_P696(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B82));
DFF_save_fm DFF_P697(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B92));
DFF_save_fm DFF_P698(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BA2));
DFF_save_fm DFF_P699(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BB2));
DFF_save_fm DFF_P700(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BC2));
DFF_save_fm DFF_P701(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BD2));
DFF_save_fm DFF_P702(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BE2));
DFF_save_fm DFF_P703(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BF2));
DFF_save_fm DFF_P704(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C02));
DFF_save_fm DFF_P705(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C12));
DFF_save_fm DFF_P706(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C22));
DFF_save_fm DFF_P707(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C32));
DFF_save_fm DFF_P708(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C42));
DFF_save_fm DFF_P709(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C52));
DFF_save_fm DFF_P710(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C62));
DFF_save_fm DFF_P711(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C72));
DFF_save_fm DFF_P712(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C82));
DFF_save_fm DFF_P713(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C92));
DFF_save_fm DFF_P714(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CA2));
DFF_save_fm DFF_P715(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CB2));
DFF_save_fm DFF_P716(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CC2));
DFF_save_fm DFF_P717(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CD2));
DFF_save_fm DFF_P718(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CE2));
DFF_save_fm DFF_P719(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CF2));
DFF_save_fm DFF_P720(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D02));
DFF_save_fm DFF_P721(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D12));
DFF_save_fm DFF_P722(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D22));
DFF_save_fm DFF_P723(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D32));
DFF_save_fm DFF_P724(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D42));
DFF_save_fm DFF_P725(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D52));
DFF_save_fm DFF_P726(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D62));
DFF_save_fm DFF_P727(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D72));
DFF_save_fm DFF_P728(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D82));
DFF_save_fm DFF_P729(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D92));
DFF_save_fm DFF_P730(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DA2));
DFF_save_fm DFF_P731(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DB2));
DFF_save_fm DFF_P732(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DC2));
DFF_save_fm DFF_P733(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DD2));
DFF_save_fm DFF_P734(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DE2));
DFF_save_fm DFF_P735(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DF2));
DFF_save_fm DFF_P736(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E02));
DFF_save_fm DFF_P737(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E12));
DFF_save_fm DFF_P738(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E22));
DFF_save_fm DFF_P739(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E32));
DFF_save_fm DFF_P740(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E42));
DFF_save_fm DFF_P741(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E52));
DFF_save_fm DFF_P742(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E62));
DFF_save_fm DFF_P743(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E72));
DFF_save_fm DFF_P744(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E82));
DFF_save_fm DFF_P745(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E92));
DFF_save_fm DFF_P746(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EA2));
DFF_save_fm DFF_P747(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EB2));
DFF_save_fm DFF_P748(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EC2));
DFF_save_fm DFF_P749(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1ED2));
DFF_save_fm DFF_P750(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EE2));
DFF_save_fm DFF_P751(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EF2));
DFF_save_fm DFF_P752(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F02));
DFF_save_fm DFF_P753(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F12));
DFF_save_fm DFF_P754(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F22));
DFF_save_fm DFF_P755(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F32));
DFF_save_fm DFF_P756(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F42));
DFF_save_fm DFF_P757(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F52));
DFF_save_fm DFF_P758(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F62));
DFF_save_fm DFF_P759(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F72));
DFF_save_fm DFF_P760(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F82));
DFF_save_fm DFF_P761(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F92));
DFF_save_fm DFF_P762(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FA2));
DFF_save_fm DFF_P763(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FB2));
DFF_save_fm DFF_P764(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FC2));
DFF_save_fm DFF_P765(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FD2));
DFF_save_fm DFF_P766(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FE2));
DFF_save_fm DFF_P767(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FF2));
DFF_save_fm DFF_P768(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1003));
DFF_save_fm DFF_P769(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1013));
DFF_save_fm DFF_P770(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1023));
DFF_save_fm DFF_P771(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1033));
DFF_save_fm DFF_P772(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1043));
DFF_save_fm DFF_P773(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1053));
DFF_save_fm DFF_P774(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1063));
DFF_save_fm DFF_P775(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1073));
DFF_save_fm DFF_P776(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1083));
DFF_save_fm DFF_P777(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1093));
DFF_save_fm DFF_P778(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10A3));
DFF_save_fm DFF_P779(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10B3));
DFF_save_fm DFF_P780(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10C3));
DFF_save_fm DFF_P781(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10D3));
DFF_save_fm DFF_P782(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10E3));
DFF_save_fm DFF_P783(.clk(clk),.rstn(rstn),.reset_value(1),.q(P10F3));
DFF_save_fm DFF_P784(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1103));
DFF_save_fm DFF_P785(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1113));
DFF_save_fm DFF_P786(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1123));
DFF_save_fm DFF_P787(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1133));
DFF_save_fm DFF_P788(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1143));
DFF_save_fm DFF_P789(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1153));
DFF_save_fm DFF_P790(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1163));
DFF_save_fm DFF_P791(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1173));
DFF_save_fm DFF_P792(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1183));
DFF_save_fm DFF_P793(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1193));
DFF_save_fm DFF_P794(.clk(clk),.rstn(rstn),.reset_value(0),.q(P11A3));
DFF_save_fm DFF_P795(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11B3));
DFF_save_fm DFF_P796(.clk(clk),.rstn(rstn),.reset_value(0),.q(P11C3));
DFF_save_fm DFF_P797(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11D3));
DFF_save_fm DFF_P798(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11E3));
DFF_save_fm DFF_P799(.clk(clk),.rstn(rstn),.reset_value(1),.q(P11F3));
DFF_save_fm DFF_P800(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1203));
DFF_save_fm DFF_P801(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1213));
DFF_save_fm DFF_P802(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1223));
DFF_save_fm DFF_P803(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1233));
DFF_save_fm DFF_P804(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1243));
DFF_save_fm DFF_P805(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1253));
DFF_save_fm DFF_P806(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1263));
DFF_save_fm DFF_P807(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1273));
DFF_save_fm DFF_P808(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1283));
DFF_save_fm DFF_P809(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1293));
DFF_save_fm DFF_P810(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12A3));
DFF_save_fm DFF_P811(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12B3));
DFF_save_fm DFF_P812(.clk(clk),.rstn(rstn),.reset_value(0),.q(P12C3));
DFF_save_fm DFF_P813(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12D3));
DFF_save_fm DFF_P814(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12E3));
DFF_save_fm DFF_P815(.clk(clk),.rstn(rstn),.reset_value(1),.q(P12F3));
DFF_save_fm DFF_P816(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1303));
DFF_save_fm DFF_P817(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1313));
DFF_save_fm DFF_P818(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1323));
DFF_save_fm DFF_P819(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1333));
DFF_save_fm DFF_P820(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1343));
DFF_save_fm DFF_P821(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1353));
DFF_save_fm DFF_P822(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1363));
DFF_save_fm DFF_P823(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1373));
DFF_save_fm DFF_P824(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1383));
DFF_save_fm DFF_P825(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1393));
DFF_save_fm DFF_P826(.clk(clk),.rstn(rstn),.reset_value(0),.q(P13A3));
DFF_save_fm DFF_P827(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13B3));
DFF_save_fm DFF_P828(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13C3));
DFF_save_fm DFF_P829(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13D3));
DFF_save_fm DFF_P830(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13E3));
DFF_save_fm DFF_P831(.clk(clk),.rstn(rstn),.reset_value(1),.q(P13F3));
DFF_save_fm DFF_P832(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1403));
DFF_save_fm DFF_P833(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1413));
DFF_save_fm DFF_P834(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1423));
DFF_save_fm DFF_P835(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1433));
DFF_save_fm DFF_P836(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1443));
DFF_save_fm DFF_P837(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1453));
DFF_save_fm DFF_P838(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1463));
DFF_save_fm DFF_P839(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1473));
DFF_save_fm DFF_P840(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1483));
DFF_save_fm DFF_P841(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1493));
DFF_save_fm DFF_P842(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14A3));
DFF_save_fm DFF_P843(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14B3));
DFF_save_fm DFF_P844(.clk(clk),.rstn(rstn),.reset_value(0),.q(P14C3));
DFF_save_fm DFF_P845(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14D3));
DFF_save_fm DFF_P846(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14E3));
DFF_save_fm DFF_P847(.clk(clk),.rstn(rstn),.reset_value(1),.q(P14F3));
DFF_save_fm DFF_P848(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1503));
DFF_save_fm DFF_P849(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1513));
DFF_save_fm DFF_P850(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1523));
DFF_save_fm DFF_P851(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1533));
DFF_save_fm DFF_P852(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1543));
DFF_save_fm DFF_P853(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1553));
DFF_save_fm DFF_P854(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1563));
DFF_save_fm DFF_P855(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1573));
DFF_save_fm DFF_P856(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1583));
DFF_save_fm DFF_P857(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1593));
DFF_save_fm DFF_P858(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15A3));
DFF_save_fm DFF_P859(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15B3));
DFF_save_fm DFF_P860(.clk(clk),.rstn(rstn),.reset_value(0),.q(P15C3));
DFF_save_fm DFF_P861(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15D3));
DFF_save_fm DFF_P862(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15E3));
DFF_save_fm DFF_P863(.clk(clk),.rstn(rstn),.reset_value(1),.q(P15F3));
DFF_save_fm DFF_P864(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1603));
DFF_save_fm DFF_P865(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1613));
DFF_save_fm DFF_P866(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1623));
DFF_save_fm DFF_P867(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1633));
DFF_save_fm DFF_P868(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1643));
DFF_save_fm DFF_P869(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1653));
DFF_save_fm DFF_P870(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1663));
DFF_save_fm DFF_P871(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1673));
DFF_save_fm DFF_P872(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1683));
DFF_save_fm DFF_P873(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1693));
DFF_save_fm DFF_P874(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16A3));
DFF_save_fm DFF_P875(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16B3));
DFF_save_fm DFF_P876(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16C3));
DFF_save_fm DFF_P877(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16D3));
DFF_save_fm DFF_P878(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16E3));
DFF_save_fm DFF_P879(.clk(clk),.rstn(rstn),.reset_value(1),.q(P16F3));
DFF_save_fm DFF_P880(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1703));
DFF_save_fm DFF_P881(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1713));
DFF_save_fm DFF_P882(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1723));
DFF_save_fm DFF_P883(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1733));
DFF_save_fm DFF_P884(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1743));
DFF_save_fm DFF_P885(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1753));
DFF_save_fm DFF_P886(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1763));
DFF_save_fm DFF_P887(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1773));
DFF_save_fm DFF_P888(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1783));
DFF_save_fm DFF_P889(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1793));
DFF_save_fm DFF_P890(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17A3));
DFF_save_fm DFF_P891(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17B3));
DFF_save_fm DFF_P892(.clk(clk),.rstn(rstn),.reset_value(0),.q(P17C3));
DFF_save_fm DFF_P893(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17D3));
DFF_save_fm DFF_P894(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17E3));
DFF_save_fm DFF_P895(.clk(clk),.rstn(rstn),.reset_value(1),.q(P17F3));
DFF_save_fm DFF_P896(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1803));
DFF_save_fm DFF_P897(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1813));
DFF_save_fm DFF_P898(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1823));
DFF_save_fm DFF_P899(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1833));
DFF_save_fm DFF_P900(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1843));
DFF_save_fm DFF_P901(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1853));
DFF_save_fm DFF_P902(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1863));
DFF_save_fm DFF_P903(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1873));
DFF_save_fm DFF_P904(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1883));
DFF_save_fm DFF_P905(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1893));
DFF_save_fm DFF_P906(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18A3));
DFF_save_fm DFF_P907(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18B3));
DFF_save_fm DFF_P908(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18C3));
DFF_save_fm DFF_P909(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18D3));
DFF_save_fm DFF_P910(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18E3));
DFF_save_fm DFF_P911(.clk(clk),.rstn(rstn),.reset_value(1),.q(P18F3));
DFF_save_fm DFF_P912(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1903));
DFF_save_fm DFF_P913(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1913));
DFF_save_fm DFF_P914(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1923));
DFF_save_fm DFF_P915(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1933));
DFF_save_fm DFF_P916(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1943));
DFF_save_fm DFF_P917(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1953));
DFF_save_fm DFF_P918(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1963));
DFF_save_fm DFF_P919(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1973));
DFF_save_fm DFF_P920(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1983));
DFF_save_fm DFF_P921(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1993));
DFF_save_fm DFF_P922(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19A3));
DFF_save_fm DFF_P923(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19B3));
DFF_save_fm DFF_P924(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19C3));
DFF_save_fm DFF_P925(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19D3));
DFF_save_fm DFF_P926(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19E3));
DFF_save_fm DFF_P927(.clk(clk),.rstn(rstn),.reset_value(1),.q(P19F3));
DFF_save_fm DFF_P928(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A03));
DFF_save_fm DFF_P929(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A13));
DFF_save_fm DFF_P930(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A23));
DFF_save_fm DFF_P931(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A33));
DFF_save_fm DFF_P932(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A43));
DFF_save_fm DFF_P933(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A53));
DFF_save_fm DFF_P934(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A63));
DFF_save_fm DFF_P935(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A73));
DFF_save_fm DFF_P936(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A83));
DFF_save_fm DFF_P937(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1A93));
DFF_save_fm DFF_P938(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AA3));
DFF_save_fm DFF_P939(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AB3));
DFF_save_fm DFF_P940(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AC3));
DFF_save_fm DFF_P941(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AD3));
DFF_save_fm DFF_P942(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AE3));
DFF_save_fm DFF_P943(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1AF3));
DFF_save_fm DFF_P944(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B03));
DFF_save_fm DFF_P945(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B13));
DFF_save_fm DFF_P946(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B23));
DFF_save_fm DFF_P947(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B33));
DFF_save_fm DFF_P948(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B43));
DFF_save_fm DFF_P949(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B53));
DFF_save_fm DFF_P950(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B63));
DFF_save_fm DFF_P951(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B73));
DFF_save_fm DFF_P952(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B83));
DFF_save_fm DFF_P953(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1B93));
DFF_save_fm DFF_P954(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BA3));
DFF_save_fm DFF_P955(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BB3));
DFF_save_fm DFF_P956(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BC3));
DFF_save_fm DFF_P957(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BD3));
DFF_save_fm DFF_P958(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BE3));
DFF_save_fm DFF_P959(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1BF3));
DFF_save_fm DFF_P960(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C03));
DFF_save_fm DFF_P961(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C13));
DFF_save_fm DFF_P962(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C23));
DFF_save_fm DFF_P963(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C33));
DFF_save_fm DFF_P964(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C43));
DFF_save_fm DFF_P965(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C53));
DFF_save_fm DFF_P966(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C63));
DFF_save_fm DFF_P967(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C73));
DFF_save_fm DFF_P968(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C83));
DFF_save_fm DFF_P969(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1C93));
DFF_save_fm DFF_P970(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1CA3));
DFF_save_fm DFF_P971(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CB3));
DFF_save_fm DFF_P972(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CC3));
DFF_save_fm DFF_P973(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CD3));
DFF_save_fm DFF_P974(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CE3));
DFF_save_fm DFF_P975(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1CF3));
DFF_save_fm DFF_P976(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D03));
DFF_save_fm DFF_P977(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D13));
DFF_save_fm DFF_P978(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D23));
DFF_save_fm DFF_P979(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D33));
DFF_save_fm DFF_P980(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D43));
DFF_save_fm DFF_P981(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D53));
DFF_save_fm DFF_P982(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D63));
DFF_save_fm DFF_P983(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1D73));
DFF_save_fm DFF_P984(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D83));
DFF_save_fm DFF_P985(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1D93));
DFF_save_fm DFF_P986(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DA3));
DFF_save_fm DFF_P987(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DB3));
DFF_save_fm DFF_P988(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DC3));
DFF_save_fm DFF_P989(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DD3));
DFF_save_fm DFF_P990(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DE3));
DFF_save_fm DFF_P991(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1DF3));
DFF_save_fm DFF_P992(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E03));
DFF_save_fm DFF_P993(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E13));
DFF_save_fm DFF_P994(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E23));
DFF_save_fm DFF_P995(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E33));
DFF_save_fm DFF_P996(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E43));
DFF_save_fm DFF_P997(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E53));
DFF_save_fm DFF_P998(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E63));
DFF_save_fm DFF_P999(.clk(clk),.rstn(rstn),.reset_value(0),.q(P1E73));
DFF_save_fm DFF_P1000(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E83));
DFF_save_fm DFF_P1001(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1E93));
DFF_save_fm DFF_P1002(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EA3));
DFF_save_fm DFF_P1003(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EB3));
DFF_save_fm DFF_P1004(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EC3));
DFF_save_fm DFF_P1005(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1ED3));
DFF_save_fm DFF_P1006(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EE3));
DFF_save_fm DFF_P1007(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1EF3));
DFF_save_fm DFF_P1008(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F03));
DFF_save_fm DFF_P1009(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F13));
DFF_save_fm DFF_P1010(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F23));
DFF_save_fm DFF_P1011(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F33));
DFF_save_fm DFF_P1012(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F43));
DFF_save_fm DFF_P1013(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F53));
DFF_save_fm DFF_P1014(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F63));
DFF_save_fm DFF_P1015(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F73));
DFF_save_fm DFF_P1016(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F83));
DFF_save_fm DFF_P1017(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1F93));
DFF_save_fm DFF_P1018(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FA3));
DFF_save_fm DFF_P1019(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FB3));
DFF_save_fm DFF_P1020(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FC3));
DFF_save_fm DFF_P1021(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FD3));
DFF_save_fm DFF_P1022(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FE3));
DFF_save_fm DFF_P1023(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1FF3));
DFF_save_fm DFF_W0(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10000));
DFF_save_fm DFF_W1(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10010));
DFF_save_fm DFF_W2(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10020));
DFF_save_fm DFF_W3(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10100));
DFF_save_fm DFF_W4(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10110));
DFF_save_fm DFF_W5(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10120));
DFF_save_fm DFF_W6(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10200));
DFF_save_fm DFF_W7(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10210));
DFF_save_fm DFF_W8(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10220));
DFF_save_fm DFF_W9(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10001));
DFF_save_fm DFF_W10(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10011));
DFF_save_fm DFF_W11(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10021));
DFF_save_fm DFF_W12(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10101));
DFF_save_fm DFF_W13(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10111));
DFF_save_fm DFF_W14(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10121));
DFF_save_fm DFF_W15(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10201));
DFF_save_fm DFF_W16(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10211));
DFF_save_fm DFF_W17(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10221));
DFF_save_fm DFF_W18(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10002));
DFF_save_fm DFF_W19(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10012));
DFF_save_fm DFF_W20(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10022));
DFF_save_fm DFF_W21(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10102));
DFF_save_fm DFF_W22(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10112));
DFF_save_fm DFF_W23(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10122));
DFF_save_fm DFF_W24(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10202));
DFF_save_fm DFF_W25(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10212));
DFF_save_fm DFF_W26(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10222));
DFF_save_fm DFF_W27(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10003));
DFF_save_fm DFF_W28(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10013));
DFF_save_fm DFF_W29(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10023));
DFF_save_fm DFF_W30(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10103));
DFF_save_fm DFF_W31(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10113));
DFF_save_fm DFF_W32(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10123));
DFF_save_fm DFF_W33(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10203));
DFF_save_fm DFF_W34(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10213));
DFF_save_fm DFF_W35(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10223));
DFF_save_fm DFF_W36(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11000));
DFF_save_fm DFF_W37(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11010));
DFF_save_fm DFF_W38(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11020));
DFF_save_fm DFF_W39(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11100));
DFF_save_fm DFF_W40(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11110));
DFF_save_fm DFF_W41(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11120));
DFF_save_fm DFF_W42(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11200));
DFF_save_fm DFF_W43(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11210));
DFF_save_fm DFF_W44(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11220));
DFF_save_fm DFF_W45(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11001));
DFF_save_fm DFF_W46(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11011));
DFF_save_fm DFF_W47(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11021));
DFF_save_fm DFF_W48(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11101));
DFF_save_fm DFF_W49(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11111));
DFF_save_fm DFF_W50(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11121));
DFF_save_fm DFF_W51(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11201));
DFF_save_fm DFF_W52(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11211));
DFF_save_fm DFF_W53(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11221));
DFF_save_fm DFF_W54(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11002));
DFF_save_fm DFF_W55(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11012));
DFF_save_fm DFF_W56(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11022));
DFF_save_fm DFF_W57(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11102));
DFF_save_fm DFF_W58(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11112));
DFF_save_fm DFF_W59(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11122));
DFF_save_fm DFF_W60(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11202));
DFF_save_fm DFF_W61(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11212));
DFF_save_fm DFF_W62(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11222));
DFF_save_fm DFF_W63(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11003));
DFF_save_fm DFF_W64(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11013));
DFF_save_fm DFF_W65(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11023));
DFF_save_fm DFF_W66(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11103));
DFF_save_fm DFF_W67(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11113));
DFF_save_fm DFF_W68(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11123));
DFF_save_fm DFF_W69(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11203));
DFF_save_fm DFF_W70(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11213));
DFF_save_fm DFF_W71(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11223));
DFF_save_fm DFF_W72(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12000));
DFF_save_fm DFF_W73(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12010));
DFF_save_fm DFF_W74(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12020));
DFF_save_fm DFF_W75(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12100));
DFF_save_fm DFF_W76(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12110));
DFF_save_fm DFF_W77(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12120));
DFF_save_fm DFF_W78(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12200));
DFF_save_fm DFF_W79(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12210));
DFF_save_fm DFF_W80(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12220));
DFF_save_fm DFF_W81(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12001));
DFF_save_fm DFF_W82(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12011));
DFF_save_fm DFF_W83(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12021));
DFF_save_fm DFF_W84(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12101));
DFF_save_fm DFF_W85(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12111));
DFF_save_fm DFF_W86(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12121));
DFF_save_fm DFF_W87(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12201));
DFF_save_fm DFF_W88(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12211));
DFF_save_fm DFF_W89(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12221));
DFF_save_fm DFF_W90(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12002));
DFF_save_fm DFF_W91(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12012));
DFF_save_fm DFF_W92(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12022));
DFF_save_fm DFF_W93(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12102));
DFF_save_fm DFF_W94(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12112));
DFF_save_fm DFF_W95(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12122));
DFF_save_fm DFF_W96(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12202));
DFF_save_fm DFF_W97(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12212));
DFF_save_fm DFF_W98(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12222));
DFF_save_fm DFF_W99(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12003));
DFF_save_fm DFF_W100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12013));
DFF_save_fm DFF_W101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12023));
DFF_save_fm DFF_W102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12103));
DFF_save_fm DFF_W103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12113));
DFF_save_fm DFF_W104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12123));
DFF_save_fm DFF_W105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12203));
DFF_save_fm DFF_W106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12213));
DFF_save_fm DFF_W107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12223));
DFF_save_fm DFF_W108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13000));
DFF_save_fm DFF_W109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13010));
DFF_save_fm DFF_W110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13020));
DFF_save_fm DFF_W111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13100));
DFF_save_fm DFF_W112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13110));
DFF_save_fm DFF_W113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13120));
DFF_save_fm DFF_W114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13200));
DFF_save_fm DFF_W115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13210));
DFF_save_fm DFF_W116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13220));
DFF_save_fm DFF_W117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13001));
DFF_save_fm DFF_W118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13011));
DFF_save_fm DFF_W119(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13021));
DFF_save_fm DFF_W120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13101));
DFF_save_fm DFF_W121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13111));
DFF_save_fm DFF_W122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13121));
DFF_save_fm DFF_W123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13201));
DFF_save_fm DFF_W124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13211));
DFF_save_fm DFF_W125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13221));
DFF_save_fm DFF_W126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13002));
DFF_save_fm DFF_W127(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13012));
DFF_save_fm DFF_W128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13022));
DFF_save_fm DFF_W129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13102));
DFF_save_fm DFF_W130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13112));
DFF_save_fm DFF_W131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13122));
DFF_save_fm DFF_W132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13202));
DFF_save_fm DFF_W133(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13212));
DFF_save_fm DFF_W134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13222));
DFF_save_fm DFF_W135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13003));
DFF_save_fm DFF_W136(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13013));
DFF_save_fm DFF_W137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13023));
DFF_save_fm DFF_W138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13103));
DFF_save_fm DFF_W139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13113));
DFF_save_fm DFF_W140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13123));
DFF_save_fm DFF_W141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13203));
DFF_save_fm DFF_W142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13213));
DFF_save_fm DFF_W143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13223));
DFF_save_fm DFF_W144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14000));
DFF_save_fm DFF_W145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14010));
DFF_save_fm DFF_W146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14020));
DFF_save_fm DFF_W147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14100));
DFF_save_fm DFF_W148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14110));
DFF_save_fm DFF_W149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14120));
DFF_save_fm DFF_W150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14200));
DFF_save_fm DFF_W151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14210));
DFF_save_fm DFF_W152(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14220));
DFF_save_fm DFF_W153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14001));
DFF_save_fm DFF_W154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14011));
DFF_save_fm DFF_W155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14021));
DFF_save_fm DFF_W156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14101));
DFF_save_fm DFF_W157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14111));
DFF_save_fm DFF_W158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14121));
DFF_save_fm DFF_W159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14201));
DFF_save_fm DFF_W160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14211));
DFF_save_fm DFF_W161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14221));
DFF_save_fm DFF_W162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14002));
DFF_save_fm DFF_W163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14012));
DFF_save_fm DFF_W164(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14022));
DFF_save_fm DFF_W165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14102));
DFF_save_fm DFF_W166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14112));
DFF_save_fm DFF_W167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14122));
DFF_save_fm DFF_W168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14202));
DFF_save_fm DFF_W169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14212));
DFF_save_fm DFF_W170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14222));
DFF_save_fm DFF_W171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14003));
DFF_save_fm DFF_W172(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14013));
DFF_save_fm DFF_W173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14023));
DFF_save_fm DFF_W174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14103));
DFF_save_fm DFF_W175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14113));
DFF_save_fm DFF_W176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14123));
DFF_save_fm DFF_W177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14203));
DFF_save_fm DFF_W178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14213));
DFF_save_fm DFF_W179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14223));
DFF_save_fm DFF_W180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15000));
DFF_save_fm DFF_W181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15010));
DFF_save_fm DFF_W182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15020));
DFF_save_fm DFF_W183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15100));
DFF_save_fm DFF_W184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15110));
DFF_save_fm DFF_W185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15120));
DFF_save_fm DFF_W186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15200));
DFF_save_fm DFF_W187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15210));
DFF_save_fm DFF_W188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15220));
DFF_save_fm DFF_W189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15001));
DFF_save_fm DFF_W190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15011));
DFF_save_fm DFF_W191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15021));
DFF_save_fm DFF_W192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15101));
DFF_save_fm DFF_W193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15111));
DFF_save_fm DFF_W194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15121));
DFF_save_fm DFF_W195(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15201));
DFF_save_fm DFF_W196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15211));
DFF_save_fm DFF_W197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15221));
DFF_save_fm DFF_W198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15002));
DFF_save_fm DFF_W199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15012));
DFF_save_fm DFF_W200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15022));
DFF_save_fm DFF_W201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15102));
DFF_save_fm DFF_W202(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15112));
DFF_save_fm DFF_W203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15122));
DFF_save_fm DFF_W204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15202));
DFF_save_fm DFF_W205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15212));
DFF_save_fm DFF_W206(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15222));
DFF_save_fm DFF_W207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15003));
DFF_save_fm DFF_W208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15013));
DFF_save_fm DFF_W209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15023));
DFF_save_fm DFF_W210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15103));
DFF_save_fm DFF_W211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15113));
DFF_save_fm DFF_W212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15123));
DFF_save_fm DFF_W213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15203));
DFF_save_fm DFF_W214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15213));
DFF_save_fm DFF_W215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15223));
DFF_save_fm DFF_W216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16000));
DFF_save_fm DFF_W217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16010));
DFF_save_fm DFF_W218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16020));
DFF_save_fm DFF_W219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16100));
DFF_save_fm DFF_W220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16110));
DFF_save_fm DFF_W221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16120));
DFF_save_fm DFF_W222(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16200));
DFF_save_fm DFF_W223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16210));
DFF_save_fm DFF_W224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16220));
DFF_save_fm DFF_W225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16001));
DFF_save_fm DFF_W226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16011));
DFF_save_fm DFF_W227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16021));
DFF_save_fm DFF_W228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16101));
DFF_save_fm DFF_W229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16111));
DFF_save_fm DFF_W230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16121));
DFF_save_fm DFF_W231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16201));
DFF_save_fm DFF_W232(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16211));
DFF_save_fm DFF_W233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16221));
DFF_save_fm DFF_W234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16002));
DFF_save_fm DFF_W235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16012));
DFF_save_fm DFF_W236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16022));
DFF_save_fm DFF_W237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16102));
DFF_save_fm DFF_W238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16112));
DFF_save_fm DFF_W239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16122));
DFF_save_fm DFF_W240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16202));
DFF_save_fm DFF_W241(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16212));
DFF_save_fm DFF_W242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16222));
DFF_save_fm DFF_W243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16003));
DFF_save_fm DFF_W244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16013));
DFF_save_fm DFF_W245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16023));
DFF_save_fm DFF_W246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16103));
DFF_save_fm DFF_W247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16113));
DFF_save_fm DFF_W248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16123));
DFF_save_fm DFF_W249(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16203));
DFF_save_fm DFF_W250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16213));
DFF_save_fm DFF_W251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16223));
DFF_save_fm DFF_W252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17000));
DFF_save_fm DFF_W253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17010));
DFF_save_fm DFF_W254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17020));
DFF_save_fm DFF_W255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17100));
DFF_save_fm DFF_W256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17110));
DFF_save_fm DFF_W257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17120));
DFF_save_fm DFF_W258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17200));
DFF_save_fm DFF_W259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17210));
DFF_save_fm DFF_W260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17220));
DFF_save_fm DFF_W261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17001));
DFF_save_fm DFF_W262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17011));
DFF_save_fm DFF_W263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17021));
DFF_save_fm DFF_W264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17101));
DFF_save_fm DFF_W265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17111));
DFF_save_fm DFF_W266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17121));
DFF_save_fm DFF_W267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17201));
DFF_save_fm DFF_W268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17211));
DFF_save_fm DFF_W269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17221));
DFF_save_fm DFF_W270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17002));
DFF_save_fm DFF_W271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17012));
DFF_save_fm DFF_W272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17022));
DFF_save_fm DFF_W273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17102));
DFF_save_fm DFF_W274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17112));
DFF_save_fm DFF_W275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17122));
DFF_save_fm DFF_W276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17202));
DFF_save_fm DFF_W277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17212));
DFF_save_fm DFF_W278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17222));
DFF_save_fm DFF_W279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17003));
DFF_save_fm DFF_W280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17013));
DFF_save_fm DFF_W281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17023));
DFF_save_fm DFF_W282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17103));
DFF_save_fm DFF_W283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17113));
DFF_save_fm DFF_W284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17123));
DFF_save_fm DFF_W285(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17203));
DFF_save_fm DFF_W286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17213));
DFF_save_fm DFF_W287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17223));
ninexnine_unit ninexnine_unit_0(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10000)
);

ninexnine_unit ninexnine_unit_1(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11000)
);

ninexnine_unit ninexnine_unit_2(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12000)
);

ninexnine_unit ninexnine_unit_3(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13000)
);

assign C1000=c10000+c11000+c12000+c13000;
assign A1000=(C1000>=0)?1:0;

ninexnine_unit ninexnine_unit_4(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10010)
);

ninexnine_unit ninexnine_unit_5(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11010)
);

ninexnine_unit ninexnine_unit_6(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12010)
);

ninexnine_unit ninexnine_unit_7(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13010)
);

assign C1010=c10010+c11010+c12010+c13010;
assign A1010=(C1010>=0)?1:0;

ninexnine_unit ninexnine_unit_8(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10020)
);

ninexnine_unit ninexnine_unit_9(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11020)
);

ninexnine_unit ninexnine_unit_10(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12020)
);

ninexnine_unit ninexnine_unit_11(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13020)
);

assign C1020=c10020+c11020+c12020+c13020;
assign A1020=(C1020>=0)?1:0;

ninexnine_unit ninexnine_unit_12(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10030)
);

ninexnine_unit ninexnine_unit_13(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11030)
);

ninexnine_unit ninexnine_unit_14(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12030)
);

ninexnine_unit ninexnine_unit_15(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13030)
);

assign C1030=c10030+c11030+c12030+c13030;
assign A1030=(C1030>=0)?1:0;

ninexnine_unit ninexnine_unit_16(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10040)
);

ninexnine_unit ninexnine_unit_17(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11040)
);

ninexnine_unit ninexnine_unit_18(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12040)
);

ninexnine_unit ninexnine_unit_19(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13040)
);

assign C1040=c10040+c11040+c12040+c13040;
assign A1040=(C1040>=0)?1:0;

ninexnine_unit ninexnine_unit_20(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10050)
);

ninexnine_unit ninexnine_unit_21(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11050)
);

ninexnine_unit ninexnine_unit_22(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12050)
);

ninexnine_unit ninexnine_unit_23(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13050)
);

assign C1050=c10050+c11050+c12050+c13050;
assign A1050=(C1050>=0)?1:0;

ninexnine_unit ninexnine_unit_24(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10060)
);

ninexnine_unit ninexnine_unit_25(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11060)
);

ninexnine_unit ninexnine_unit_26(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12060)
);

ninexnine_unit ninexnine_unit_27(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13060)
);

assign C1060=c10060+c11060+c12060+c13060;
assign A1060=(C1060>=0)?1:0;

ninexnine_unit ninexnine_unit_28(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10070)
);

ninexnine_unit ninexnine_unit_29(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11070)
);

ninexnine_unit ninexnine_unit_30(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12070)
);

ninexnine_unit ninexnine_unit_31(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13070)
);

assign C1070=c10070+c11070+c12070+c13070;
assign A1070=(C1070>=0)?1:0;

ninexnine_unit ninexnine_unit_32(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10080)
);

ninexnine_unit ninexnine_unit_33(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11080)
);

ninexnine_unit ninexnine_unit_34(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12080)
);

ninexnine_unit ninexnine_unit_35(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13080)
);

assign C1080=c10080+c11080+c12080+c13080;
assign A1080=(C1080>=0)?1:0;

ninexnine_unit ninexnine_unit_36(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10090)
);

ninexnine_unit ninexnine_unit_37(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11090)
);

ninexnine_unit ninexnine_unit_38(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12090)
);

ninexnine_unit ninexnine_unit_39(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13090)
);

assign C1090=c10090+c11090+c12090+c13090;
assign A1090=(C1090>=0)?1:0;

ninexnine_unit ninexnine_unit_40(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c100A0)
);

ninexnine_unit ninexnine_unit_41(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c110A0)
);

ninexnine_unit ninexnine_unit_42(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c120A0)
);

ninexnine_unit ninexnine_unit_43(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c130A0)
);

assign C10A0=c100A0+c110A0+c120A0+c130A0;
assign A10A0=(C10A0>=0)?1:0;

ninexnine_unit ninexnine_unit_44(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c100B0)
);

ninexnine_unit ninexnine_unit_45(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c110B0)
);

ninexnine_unit ninexnine_unit_46(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c120B0)
);

ninexnine_unit ninexnine_unit_47(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c130B0)
);

assign C10B0=c100B0+c110B0+c120B0+c130B0;
assign A10B0=(C10B0>=0)?1:0;

ninexnine_unit ninexnine_unit_48(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c100C0)
);

ninexnine_unit ninexnine_unit_49(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c110C0)
);

ninexnine_unit ninexnine_unit_50(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c120C0)
);

ninexnine_unit ninexnine_unit_51(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c130C0)
);

assign C10C0=c100C0+c110C0+c120C0+c130C0;
assign A10C0=(C10C0>=0)?1:0;

ninexnine_unit ninexnine_unit_52(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c100D0)
);

ninexnine_unit ninexnine_unit_53(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c110D0)
);

ninexnine_unit ninexnine_unit_54(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c120D0)
);

ninexnine_unit ninexnine_unit_55(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c130D0)
);

assign C10D0=c100D0+c110D0+c120D0+c130D0;
assign A10D0=(C10D0>=0)?1:0;

ninexnine_unit ninexnine_unit_56(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10100)
);

ninexnine_unit ninexnine_unit_57(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11100)
);

ninexnine_unit ninexnine_unit_58(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12100)
);

ninexnine_unit ninexnine_unit_59(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13100)
);

assign C1100=c10100+c11100+c12100+c13100;
assign A1100=(C1100>=0)?1:0;

ninexnine_unit ninexnine_unit_60(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10110)
);

ninexnine_unit ninexnine_unit_61(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11110)
);

ninexnine_unit ninexnine_unit_62(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12110)
);

ninexnine_unit ninexnine_unit_63(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13110)
);

assign C1110=c10110+c11110+c12110+c13110;
assign A1110=(C1110>=0)?1:0;

ninexnine_unit ninexnine_unit_64(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10120)
);

ninexnine_unit ninexnine_unit_65(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11120)
);

ninexnine_unit ninexnine_unit_66(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12120)
);

ninexnine_unit ninexnine_unit_67(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13120)
);

assign C1120=c10120+c11120+c12120+c13120;
assign A1120=(C1120>=0)?1:0;

ninexnine_unit ninexnine_unit_68(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10130)
);

ninexnine_unit ninexnine_unit_69(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11130)
);

ninexnine_unit ninexnine_unit_70(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12130)
);

ninexnine_unit ninexnine_unit_71(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13130)
);

assign C1130=c10130+c11130+c12130+c13130;
assign A1130=(C1130>=0)?1:0;

ninexnine_unit ninexnine_unit_72(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10140)
);

ninexnine_unit ninexnine_unit_73(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11140)
);

ninexnine_unit ninexnine_unit_74(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12140)
);

ninexnine_unit ninexnine_unit_75(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13140)
);

assign C1140=c10140+c11140+c12140+c13140;
assign A1140=(C1140>=0)?1:0;

ninexnine_unit ninexnine_unit_76(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10150)
);

ninexnine_unit ninexnine_unit_77(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11150)
);

ninexnine_unit ninexnine_unit_78(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12150)
);

ninexnine_unit ninexnine_unit_79(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13150)
);

assign C1150=c10150+c11150+c12150+c13150;
assign A1150=(C1150>=0)?1:0;

ninexnine_unit ninexnine_unit_80(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10160)
);

ninexnine_unit ninexnine_unit_81(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11160)
);

ninexnine_unit ninexnine_unit_82(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12160)
);

ninexnine_unit ninexnine_unit_83(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13160)
);

assign C1160=c10160+c11160+c12160+c13160;
assign A1160=(C1160>=0)?1:0;

ninexnine_unit ninexnine_unit_84(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10170)
);

ninexnine_unit ninexnine_unit_85(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11170)
);

ninexnine_unit ninexnine_unit_86(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12170)
);

ninexnine_unit ninexnine_unit_87(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13170)
);

assign C1170=c10170+c11170+c12170+c13170;
assign A1170=(C1170>=0)?1:0;

ninexnine_unit ninexnine_unit_88(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10180)
);

ninexnine_unit ninexnine_unit_89(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11180)
);

ninexnine_unit ninexnine_unit_90(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12180)
);

ninexnine_unit ninexnine_unit_91(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13180)
);

assign C1180=c10180+c11180+c12180+c13180;
assign A1180=(C1180>=0)?1:0;

ninexnine_unit ninexnine_unit_92(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10190)
);

ninexnine_unit ninexnine_unit_93(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11190)
);

ninexnine_unit ninexnine_unit_94(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12190)
);

ninexnine_unit ninexnine_unit_95(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13190)
);

assign C1190=c10190+c11190+c12190+c13190;
assign A1190=(C1190>=0)?1:0;

ninexnine_unit ninexnine_unit_96(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c101A0)
);

ninexnine_unit ninexnine_unit_97(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c111A0)
);

ninexnine_unit ninexnine_unit_98(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c121A0)
);

ninexnine_unit ninexnine_unit_99(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c131A0)
);

assign C11A0=c101A0+c111A0+c121A0+c131A0;
assign A11A0=(C11A0>=0)?1:0;

ninexnine_unit ninexnine_unit_100(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c101B0)
);

ninexnine_unit ninexnine_unit_101(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c111B0)
);

ninexnine_unit ninexnine_unit_102(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c121B0)
);

ninexnine_unit ninexnine_unit_103(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c131B0)
);

assign C11B0=c101B0+c111B0+c121B0+c131B0;
assign A11B0=(C11B0>=0)?1:0;

ninexnine_unit ninexnine_unit_104(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c101C0)
);

ninexnine_unit ninexnine_unit_105(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c111C0)
);

ninexnine_unit ninexnine_unit_106(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c121C0)
);

ninexnine_unit ninexnine_unit_107(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c131C0)
);

assign C11C0=c101C0+c111C0+c121C0+c131C0;
assign A11C0=(C11C0>=0)?1:0;

ninexnine_unit ninexnine_unit_108(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c101D0)
);

ninexnine_unit ninexnine_unit_109(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c111D0)
);

ninexnine_unit ninexnine_unit_110(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c121D0)
);

ninexnine_unit ninexnine_unit_111(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c131D0)
);

assign C11D0=c101D0+c111D0+c121D0+c131D0;
assign A11D0=(C11D0>=0)?1:0;

ninexnine_unit ninexnine_unit_112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10200)
);

ninexnine_unit ninexnine_unit_113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11200)
);

ninexnine_unit ninexnine_unit_114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12200)
);

ninexnine_unit ninexnine_unit_115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13200)
);

assign C1200=c10200+c11200+c12200+c13200;
assign A1200=(C1200>=0)?1:0;

ninexnine_unit ninexnine_unit_116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10210)
);

ninexnine_unit ninexnine_unit_117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11210)
);

ninexnine_unit ninexnine_unit_118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12210)
);

ninexnine_unit ninexnine_unit_119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13210)
);

assign C1210=c10210+c11210+c12210+c13210;
assign A1210=(C1210>=0)?1:0;

ninexnine_unit ninexnine_unit_120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10220)
);

ninexnine_unit ninexnine_unit_121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11220)
);

ninexnine_unit ninexnine_unit_122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12220)
);

ninexnine_unit ninexnine_unit_123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13220)
);

assign C1220=c10220+c11220+c12220+c13220;
assign A1220=(C1220>=0)?1:0;

ninexnine_unit ninexnine_unit_124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10230)
);

ninexnine_unit ninexnine_unit_125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11230)
);

ninexnine_unit ninexnine_unit_126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12230)
);

ninexnine_unit ninexnine_unit_127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13230)
);

assign C1230=c10230+c11230+c12230+c13230;
assign A1230=(C1230>=0)?1:0;

ninexnine_unit ninexnine_unit_128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10240)
);

ninexnine_unit ninexnine_unit_129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11240)
);

ninexnine_unit ninexnine_unit_130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12240)
);

ninexnine_unit ninexnine_unit_131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13240)
);

assign C1240=c10240+c11240+c12240+c13240;
assign A1240=(C1240>=0)?1:0;

ninexnine_unit ninexnine_unit_132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10250)
);

ninexnine_unit ninexnine_unit_133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11250)
);

ninexnine_unit ninexnine_unit_134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12250)
);

ninexnine_unit ninexnine_unit_135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13250)
);

assign C1250=c10250+c11250+c12250+c13250;
assign A1250=(C1250>=0)?1:0;

ninexnine_unit ninexnine_unit_136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10260)
);

ninexnine_unit ninexnine_unit_137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11260)
);

ninexnine_unit ninexnine_unit_138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12260)
);

ninexnine_unit ninexnine_unit_139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13260)
);

assign C1260=c10260+c11260+c12260+c13260;
assign A1260=(C1260>=0)?1:0;

ninexnine_unit ninexnine_unit_140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10270)
);

ninexnine_unit ninexnine_unit_141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11270)
);

ninexnine_unit ninexnine_unit_142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12270)
);

ninexnine_unit ninexnine_unit_143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13270)
);

assign C1270=c10270+c11270+c12270+c13270;
assign A1270=(C1270>=0)?1:0;

ninexnine_unit ninexnine_unit_144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10280)
);

ninexnine_unit ninexnine_unit_145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11280)
);

ninexnine_unit ninexnine_unit_146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12280)
);

ninexnine_unit ninexnine_unit_147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13280)
);

assign C1280=c10280+c11280+c12280+c13280;
assign A1280=(C1280>=0)?1:0;

ninexnine_unit ninexnine_unit_148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10290)
);

ninexnine_unit ninexnine_unit_149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11290)
);

ninexnine_unit ninexnine_unit_150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12290)
);

ninexnine_unit ninexnine_unit_151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13290)
);

assign C1290=c10290+c11290+c12290+c13290;
assign A1290=(C1290>=0)?1:0;

ninexnine_unit ninexnine_unit_152(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c102A0)
);

ninexnine_unit ninexnine_unit_153(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c112A0)
);

ninexnine_unit ninexnine_unit_154(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c122A0)
);

ninexnine_unit ninexnine_unit_155(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c132A0)
);

assign C12A0=c102A0+c112A0+c122A0+c132A0;
assign A12A0=(C12A0>=0)?1:0;

ninexnine_unit ninexnine_unit_156(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c102B0)
);

ninexnine_unit ninexnine_unit_157(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c112B0)
);

ninexnine_unit ninexnine_unit_158(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c122B0)
);

ninexnine_unit ninexnine_unit_159(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c132B0)
);

assign C12B0=c102B0+c112B0+c122B0+c132B0;
assign A12B0=(C12B0>=0)?1:0;

ninexnine_unit ninexnine_unit_160(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c102C0)
);

ninexnine_unit ninexnine_unit_161(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c112C0)
);

ninexnine_unit ninexnine_unit_162(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c122C0)
);

ninexnine_unit ninexnine_unit_163(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c132C0)
);

assign C12C0=c102C0+c112C0+c122C0+c132C0;
assign A12C0=(C12C0>=0)?1:0;

ninexnine_unit ninexnine_unit_164(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c102D0)
);

ninexnine_unit ninexnine_unit_165(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c112D0)
);

ninexnine_unit ninexnine_unit_166(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c122D0)
);

ninexnine_unit ninexnine_unit_167(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c132D0)
);

assign C12D0=c102D0+c112D0+c122D0+c132D0;
assign A12D0=(C12D0>=0)?1:0;

ninexnine_unit ninexnine_unit_168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10300)
);

ninexnine_unit ninexnine_unit_169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11300)
);

ninexnine_unit ninexnine_unit_170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12300)
);

ninexnine_unit ninexnine_unit_171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13300)
);

assign C1300=c10300+c11300+c12300+c13300;
assign A1300=(C1300>=0)?1:0;

ninexnine_unit ninexnine_unit_172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10310)
);

ninexnine_unit ninexnine_unit_173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11310)
);

ninexnine_unit ninexnine_unit_174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12310)
);

ninexnine_unit ninexnine_unit_175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13310)
);

assign C1310=c10310+c11310+c12310+c13310;
assign A1310=(C1310>=0)?1:0;

ninexnine_unit ninexnine_unit_176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10320)
);

ninexnine_unit ninexnine_unit_177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11320)
);

ninexnine_unit ninexnine_unit_178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12320)
);

ninexnine_unit ninexnine_unit_179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13320)
);

assign C1320=c10320+c11320+c12320+c13320;
assign A1320=(C1320>=0)?1:0;

ninexnine_unit ninexnine_unit_180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10330)
);

ninexnine_unit ninexnine_unit_181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11330)
);

ninexnine_unit ninexnine_unit_182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12330)
);

ninexnine_unit ninexnine_unit_183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13330)
);

assign C1330=c10330+c11330+c12330+c13330;
assign A1330=(C1330>=0)?1:0;

ninexnine_unit ninexnine_unit_184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10340)
);

ninexnine_unit ninexnine_unit_185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11340)
);

ninexnine_unit ninexnine_unit_186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12340)
);

ninexnine_unit ninexnine_unit_187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13340)
);

assign C1340=c10340+c11340+c12340+c13340;
assign A1340=(C1340>=0)?1:0;

ninexnine_unit ninexnine_unit_188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10350)
);

ninexnine_unit ninexnine_unit_189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11350)
);

ninexnine_unit ninexnine_unit_190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12350)
);

ninexnine_unit ninexnine_unit_191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13350)
);

assign C1350=c10350+c11350+c12350+c13350;
assign A1350=(C1350>=0)?1:0;

ninexnine_unit ninexnine_unit_192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10360)
);

ninexnine_unit ninexnine_unit_193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11360)
);

ninexnine_unit ninexnine_unit_194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12360)
);

ninexnine_unit ninexnine_unit_195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13360)
);

assign C1360=c10360+c11360+c12360+c13360;
assign A1360=(C1360>=0)?1:0;

ninexnine_unit ninexnine_unit_196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10370)
);

ninexnine_unit ninexnine_unit_197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11370)
);

ninexnine_unit ninexnine_unit_198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12370)
);

ninexnine_unit ninexnine_unit_199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13370)
);

assign C1370=c10370+c11370+c12370+c13370;
assign A1370=(C1370>=0)?1:0;

ninexnine_unit ninexnine_unit_200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10380)
);

ninexnine_unit ninexnine_unit_201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11380)
);

ninexnine_unit ninexnine_unit_202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12380)
);

ninexnine_unit ninexnine_unit_203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13380)
);

assign C1380=c10380+c11380+c12380+c13380;
assign A1380=(C1380>=0)?1:0;

ninexnine_unit ninexnine_unit_204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10390)
);

ninexnine_unit ninexnine_unit_205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11390)
);

ninexnine_unit ninexnine_unit_206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12390)
);

ninexnine_unit ninexnine_unit_207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13390)
);

assign C1390=c10390+c11390+c12390+c13390;
assign A1390=(C1390>=0)?1:0;

ninexnine_unit ninexnine_unit_208(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c103A0)
);

ninexnine_unit ninexnine_unit_209(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c113A0)
);

ninexnine_unit ninexnine_unit_210(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c123A0)
);

ninexnine_unit ninexnine_unit_211(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c133A0)
);

assign C13A0=c103A0+c113A0+c123A0+c133A0;
assign A13A0=(C13A0>=0)?1:0;

ninexnine_unit ninexnine_unit_212(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c103B0)
);

ninexnine_unit ninexnine_unit_213(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c113B0)
);

ninexnine_unit ninexnine_unit_214(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c123B0)
);

ninexnine_unit ninexnine_unit_215(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c133B0)
);

assign C13B0=c103B0+c113B0+c123B0+c133B0;
assign A13B0=(C13B0>=0)?1:0;

ninexnine_unit ninexnine_unit_216(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c103C0)
);

ninexnine_unit ninexnine_unit_217(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c113C0)
);

ninexnine_unit ninexnine_unit_218(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c123C0)
);

ninexnine_unit ninexnine_unit_219(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c133C0)
);

assign C13C0=c103C0+c113C0+c123C0+c133C0;
assign A13C0=(C13C0>=0)?1:0;

ninexnine_unit ninexnine_unit_220(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c103D0)
);

ninexnine_unit ninexnine_unit_221(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c113D0)
);

ninexnine_unit ninexnine_unit_222(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c123D0)
);

ninexnine_unit ninexnine_unit_223(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c133D0)
);

assign C13D0=c103D0+c113D0+c123D0+c133D0;
assign A13D0=(C13D0>=0)?1:0;

ninexnine_unit ninexnine_unit_224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10400)
);

ninexnine_unit ninexnine_unit_225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11400)
);

ninexnine_unit ninexnine_unit_226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12400)
);

ninexnine_unit ninexnine_unit_227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13400)
);

assign C1400=c10400+c11400+c12400+c13400;
assign A1400=(C1400>=0)?1:0;

ninexnine_unit ninexnine_unit_228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10410)
);

ninexnine_unit ninexnine_unit_229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11410)
);

ninexnine_unit ninexnine_unit_230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12410)
);

ninexnine_unit ninexnine_unit_231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13410)
);

assign C1410=c10410+c11410+c12410+c13410;
assign A1410=(C1410>=0)?1:0;

ninexnine_unit ninexnine_unit_232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10420)
);

ninexnine_unit ninexnine_unit_233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11420)
);

ninexnine_unit ninexnine_unit_234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12420)
);

ninexnine_unit ninexnine_unit_235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13420)
);

assign C1420=c10420+c11420+c12420+c13420;
assign A1420=(C1420>=0)?1:0;

ninexnine_unit ninexnine_unit_236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10430)
);

ninexnine_unit ninexnine_unit_237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11430)
);

ninexnine_unit ninexnine_unit_238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12430)
);

ninexnine_unit ninexnine_unit_239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13430)
);

assign C1430=c10430+c11430+c12430+c13430;
assign A1430=(C1430>=0)?1:0;

ninexnine_unit ninexnine_unit_240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10440)
);

ninexnine_unit ninexnine_unit_241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11440)
);

ninexnine_unit ninexnine_unit_242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12440)
);

ninexnine_unit ninexnine_unit_243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13440)
);

assign C1440=c10440+c11440+c12440+c13440;
assign A1440=(C1440>=0)?1:0;

ninexnine_unit ninexnine_unit_244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10450)
);

ninexnine_unit ninexnine_unit_245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11450)
);

ninexnine_unit ninexnine_unit_246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12450)
);

ninexnine_unit ninexnine_unit_247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13450)
);

assign C1450=c10450+c11450+c12450+c13450;
assign A1450=(C1450>=0)?1:0;

ninexnine_unit ninexnine_unit_248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10460)
);

ninexnine_unit ninexnine_unit_249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11460)
);

ninexnine_unit ninexnine_unit_250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12460)
);

ninexnine_unit ninexnine_unit_251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13460)
);

assign C1460=c10460+c11460+c12460+c13460;
assign A1460=(C1460>=0)?1:0;

ninexnine_unit ninexnine_unit_252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10470)
);

ninexnine_unit ninexnine_unit_253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11470)
);

ninexnine_unit ninexnine_unit_254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12470)
);

ninexnine_unit ninexnine_unit_255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13470)
);

assign C1470=c10470+c11470+c12470+c13470;
assign A1470=(C1470>=0)?1:0;

ninexnine_unit ninexnine_unit_256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10480)
);

ninexnine_unit ninexnine_unit_257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11480)
);

ninexnine_unit ninexnine_unit_258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12480)
);

ninexnine_unit ninexnine_unit_259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13480)
);

assign C1480=c10480+c11480+c12480+c13480;
assign A1480=(C1480>=0)?1:0;

ninexnine_unit ninexnine_unit_260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10490)
);

ninexnine_unit ninexnine_unit_261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11490)
);

ninexnine_unit ninexnine_unit_262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12490)
);

ninexnine_unit ninexnine_unit_263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13490)
);

assign C1490=c10490+c11490+c12490+c13490;
assign A1490=(C1490>=0)?1:0;

ninexnine_unit ninexnine_unit_264(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c104A0)
);

ninexnine_unit ninexnine_unit_265(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c114A0)
);

ninexnine_unit ninexnine_unit_266(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c124A0)
);

ninexnine_unit ninexnine_unit_267(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c134A0)
);

assign C14A0=c104A0+c114A0+c124A0+c134A0;
assign A14A0=(C14A0>=0)?1:0;

ninexnine_unit ninexnine_unit_268(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c104B0)
);

ninexnine_unit ninexnine_unit_269(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c114B0)
);

ninexnine_unit ninexnine_unit_270(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c124B0)
);

ninexnine_unit ninexnine_unit_271(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c134B0)
);

assign C14B0=c104B0+c114B0+c124B0+c134B0;
assign A14B0=(C14B0>=0)?1:0;

ninexnine_unit ninexnine_unit_272(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c104C0)
);

ninexnine_unit ninexnine_unit_273(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c114C0)
);

ninexnine_unit ninexnine_unit_274(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c124C0)
);

ninexnine_unit ninexnine_unit_275(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c134C0)
);

assign C14C0=c104C0+c114C0+c124C0+c134C0;
assign A14C0=(C14C0>=0)?1:0;

ninexnine_unit ninexnine_unit_276(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c104D0)
);

ninexnine_unit ninexnine_unit_277(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c114D0)
);

ninexnine_unit ninexnine_unit_278(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c124D0)
);

ninexnine_unit ninexnine_unit_279(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c134D0)
);

assign C14D0=c104D0+c114D0+c124D0+c134D0;
assign A14D0=(C14D0>=0)?1:0;

ninexnine_unit ninexnine_unit_280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10500)
);

ninexnine_unit ninexnine_unit_281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11500)
);

ninexnine_unit ninexnine_unit_282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12500)
);

ninexnine_unit ninexnine_unit_283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13500)
);

assign C1500=c10500+c11500+c12500+c13500;
assign A1500=(C1500>=0)?1:0;

ninexnine_unit ninexnine_unit_284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10510)
);

ninexnine_unit ninexnine_unit_285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11510)
);

ninexnine_unit ninexnine_unit_286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12510)
);

ninexnine_unit ninexnine_unit_287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13510)
);

assign C1510=c10510+c11510+c12510+c13510;
assign A1510=(C1510>=0)?1:0;

ninexnine_unit ninexnine_unit_288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10520)
);

ninexnine_unit ninexnine_unit_289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11520)
);

ninexnine_unit ninexnine_unit_290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12520)
);

ninexnine_unit ninexnine_unit_291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13520)
);

assign C1520=c10520+c11520+c12520+c13520;
assign A1520=(C1520>=0)?1:0;

ninexnine_unit ninexnine_unit_292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10530)
);

ninexnine_unit ninexnine_unit_293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11530)
);

ninexnine_unit ninexnine_unit_294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12530)
);

ninexnine_unit ninexnine_unit_295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13530)
);

assign C1530=c10530+c11530+c12530+c13530;
assign A1530=(C1530>=0)?1:0;

ninexnine_unit ninexnine_unit_296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10540)
);

ninexnine_unit ninexnine_unit_297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11540)
);

ninexnine_unit ninexnine_unit_298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12540)
);

ninexnine_unit ninexnine_unit_299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13540)
);

assign C1540=c10540+c11540+c12540+c13540;
assign A1540=(C1540>=0)?1:0;

ninexnine_unit ninexnine_unit_300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10550)
);

ninexnine_unit ninexnine_unit_301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11550)
);

ninexnine_unit ninexnine_unit_302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12550)
);

ninexnine_unit ninexnine_unit_303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13550)
);

assign C1550=c10550+c11550+c12550+c13550;
assign A1550=(C1550>=0)?1:0;

ninexnine_unit ninexnine_unit_304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10560)
);

ninexnine_unit ninexnine_unit_305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11560)
);

ninexnine_unit ninexnine_unit_306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12560)
);

ninexnine_unit ninexnine_unit_307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13560)
);

assign C1560=c10560+c11560+c12560+c13560;
assign A1560=(C1560>=0)?1:0;

ninexnine_unit ninexnine_unit_308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10570)
);

ninexnine_unit ninexnine_unit_309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11570)
);

ninexnine_unit ninexnine_unit_310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12570)
);

ninexnine_unit ninexnine_unit_311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13570)
);

assign C1570=c10570+c11570+c12570+c13570;
assign A1570=(C1570>=0)?1:0;

ninexnine_unit ninexnine_unit_312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10580)
);

ninexnine_unit ninexnine_unit_313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11580)
);

ninexnine_unit ninexnine_unit_314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12580)
);

ninexnine_unit ninexnine_unit_315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13580)
);

assign C1580=c10580+c11580+c12580+c13580;
assign A1580=(C1580>=0)?1:0;

ninexnine_unit ninexnine_unit_316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10590)
);

ninexnine_unit ninexnine_unit_317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11590)
);

ninexnine_unit ninexnine_unit_318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12590)
);

ninexnine_unit ninexnine_unit_319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13590)
);

assign C1590=c10590+c11590+c12590+c13590;
assign A1590=(C1590>=0)?1:0;

ninexnine_unit ninexnine_unit_320(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c105A0)
);

ninexnine_unit ninexnine_unit_321(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c115A0)
);

ninexnine_unit ninexnine_unit_322(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c125A0)
);

ninexnine_unit ninexnine_unit_323(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c135A0)
);

assign C15A0=c105A0+c115A0+c125A0+c135A0;
assign A15A0=(C15A0>=0)?1:0;

ninexnine_unit ninexnine_unit_324(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c105B0)
);

ninexnine_unit ninexnine_unit_325(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c115B0)
);

ninexnine_unit ninexnine_unit_326(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c125B0)
);

ninexnine_unit ninexnine_unit_327(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c135B0)
);

assign C15B0=c105B0+c115B0+c125B0+c135B0;
assign A15B0=(C15B0>=0)?1:0;

ninexnine_unit ninexnine_unit_328(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c105C0)
);

ninexnine_unit ninexnine_unit_329(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c115C0)
);

ninexnine_unit ninexnine_unit_330(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c125C0)
);

ninexnine_unit ninexnine_unit_331(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c135C0)
);

assign C15C0=c105C0+c115C0+c125C0+c135C0;
assign A15C0=(C15C0>=0)?1:0;

ninexnine_unit ninexnine_unit_332(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c105D0)
);

ninexnine_unit ninexnine_unit_333(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c115D0)
);

ninexnine_unit ninexnine_unit_334(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c125D0)
);

ninexnine_unit ninexnine_unit_335(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c135D0)
);

assign C15D0=c105D0+c115D0+c125D0+c135D0;
assign A15D0=(C15D0>=0)?1:0;

ninexnine_unit ninexnine_unit_336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10600)
);

ninexnine_unit ninexnine_unit_337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11600)
);

ninexnine_unit ninexnine_unit_338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12600)
);

ninexnine_unit ninexnine_unit_339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13600)
);

assign C1600=c10600+c11600+c12600+c13600;
assign A1600=(C1600>=0)?1:0;

ninexnine_unit ninexnine_unit_340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10610)
);

ninexnine_unit ninexnine_unit_341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11610)
);

ninexnine_unit ninexnine_unit_342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12610)
);

ninexnine_unit ninexnine_unit_343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13610)
);

assign C1610=c10610+c11610+c12610+c13610;
assign A1610=(C1610>=0)?1:0;

ninexnine_unit ninexnine_unit_344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10620)
);

ninexnine_unit ninexnine_unit_345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11620)
);

ninexnine_unit ninexnine_unit_346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12620)
);

ninexnine_unit ninexnine_unit_347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13620)
);

assign C1620=c10620+c11620+c12620+c13620;
assign A1620=(C1620>=0)?1:0;

ninexnine_unit ninexnine_unit_348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10630)
);

ninexnine_unit ninexnine_unit_349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11630)
);

ninexnine_unit ninexnine_unit_350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12630)
);

ninexnine_unit ninexnine_unit_351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13630)
);

assign C1630=c10630+c11630+c12630+c13630;
assign A1630=(C1630>=0)?1:0;

ninexnine_unit ninexnine_unit_352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10640)
);

ninexnine_unit ninexnine_unit_353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11640)
);

ninexnine_unit ninexnine_unit_354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12640)
);

ninexnine_unit ninexnine_unit_355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13640)
);

assign C1640=c10640+c11640+c12640+c13640;
assign A1640=(C1640>=0)?1:0;

ninexnine_unit ninexnine_unit_356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10650)
);

ninexnine_unit ninexnine_unit_357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11650)
);

ninexnine_unit ninexnine_unit_358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12650)
);

ninexnine_unit ninexnine_unit_359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13650)
);

assign C1650=c10650+c11650+c12650+c13650;
assign A1650=(C1650>=0)?1:0;

ninexnine_unit ninexnine_unit_360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10660)
);

ninexnine_unit ninexnine_unit_361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11660)
);

ninexnine_unit ninexnine_unit_362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12660)
);

ninexnine_unit ninexnine_unit_363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13660)
);

assign C1660=c10660+c11660+c12660+c13660;
assign A1660=(C1660>=0)?1:0;

ninexnine_unit ninexnine_unit_364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10670)
);

ninexnine_unit ninexnine_unit_365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11670)
);

ninexnine_unit ninexnine_unit_366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12670)
);

ninexnine_unit ninexnine_unit_367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13670)
);

assign C1670=c10670+c11670+c12670+c13670;
assign A1670=(C1670>=0)?1:0;

ninexnine_unit ninexnine_unit_368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10680)
);

ninexnine_unit ninexnine_unit_369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11680)
);

ninexnine_unit ninexnine_unit_370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12680)
);

ninexnine_unit ninexnine_unit_371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13680)
);

assign C1680=c10680+c11680+c12680+c13680;
assign A1680=(C1680>=0)?1:0;

ninexnine_unit ninexnine_unit_372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10690)
);

ninexnine_unit ninexnine_unit_373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11690)
);

ninexnine_unit ninexnine_unit_374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12690)
);

ninexnine_unit ninexnine_unit_375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13690)
);

assign C1690=c10690+c11690+c12690+c13690;
assign A1690=(C1690>=0)?1:0;

ninexnine_unit ninexnine_unit_376(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c106A0)
);

ninexnine_unit ninexnine_unit_377(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c116A0)
);

ninexnine_unit ninexnine_unit_378(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c126A0)
);

ninexnine_unit ninexnine_unit_379(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c136A0)
);

assign C16A0=c106A0+c116A0+c126A0+c136A0;
assign A16A0=(C16A0>=0)?1:0;

ninexnine_unit ninexnine_unit_380(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c106B0)
);

ninexnine_unit ninexnine_unit_381(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c116B0)
);

ninexnine_unit ninexnine_unit_382(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c126B0)
);

ninexnine_unit ninexnine_unit_383(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c136B0)
);

assign C16B0=c106B0+c116B0+c126B0+c136B0;
assign A16B0=(C16B0>=0)?1:0;

ninexnine_unit ninexnine_unit_384(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c106C0)
);

ninexnine_unit ninexnine_unit_385(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c116C0)
);

ninexnine_unit ninexnine_unit_386(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c126C0)
);

ninexnine_unit ninexnine_unit_387(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c136C0)
);

assign C16C0=c106C0+c116C0+c126C0+c136C0;
assign A16C0=(C16C0>=0)?1:0;

ninexnine_unit ninexnine_unit_388(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c106D0)
);

ninexnine_unit ninexnine_unit_389(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c116D0)
);

ninexnine_unit ninexnine_unit_390(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c126D0)
);

ninexnine_unit ninexnine_unit_391(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c136D0)
);

assign C16D0=c106D0+c116D0+c126D0+c136D0;
assign A16D0=(C16D0>=0)?1:0;

ninexnine_unit ninexnine_unit_392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10700)
);

ninexnine_unit ninexnine_unit_393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11700)
);

ninexnine_unit ninexnine_unit_394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12700)
);

ninexnine_unit ninexnine_unit_395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13700)
);

assign C1700=c10700+c11700+c12700+c13700;
assign A1700=(C1700>=0)?1:0;

ninexnine_unit ninexnine_unit_396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10710)
);

ninexnine_unit ninexnine_unit_397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11710)
);

ninexnine_unit ninexnine_unit_398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12710)
);

ninexnine_unit ninexnine_unit_399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13710)
);

assign C1710=c10710+c11710+c12710+c13710;
assign A1710=(C1710>=0)?1:0;

ninexnine_unit ninexnine_unit_400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10720)
);

ninexnine_unit ninexnine_unit_401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11720)
);

ninexnine_unit ninexnine_unit_402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12720)
);

ninexnine_unit ninexnine_unit_403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13720)
);

assign C1720=c10720+c11720+c12720+c13720;
assign A1720=(C1720>=0)?1:0;

ninexnine_unit ninexnine_unit_404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10730)
);

ninexnine_unit ninexnine_unit_405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11730)
);

ninexnine_unit ninexnine_unit_406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12730)
);

ninexnine_unit ninexnine_unit_407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13730)
);

assign C1730=c10730+c11730+c12730+c13730;
assign A1730=(C1730>=0)?1:0;

ninexnine_unit ninexnine_unit_408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10740)
);

ninexnine_unit ninexnine_unit_409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11740)
);

ninexnine_unit ninexnine_unit_410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12740)
);

ninexnine_unit ninexnine_unit_411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13740)
);

assign C1740=c10740+c11740+c12740+c13740;
assign A1740=(C1740>=0)?1:0;

ninexnine_unit ninexnine_unit_412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10750)
);

ninexnine_unit ninexnine_unit_413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11750)
);

ninexnine_unit ninexnine_unit_414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12750)
);

ninexnine_unit ninexnine_unit_415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13750)
);

assign C1750=c10750+c11750+c12750+c13750;
assign A1750=(C1750>=0)?1:0;

ninexnine_unit ninexnine_unit_416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10760)
);

ninexnine_unit ninexnine_unit_417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11760)
);

ninexnine_unit ninexnine_unit_418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12760)
);

ninexnine_unit ninexnine_unit_419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13760)
);

assign C1760=c10760+c11760+c12760+c13760;
assign A1760=(C1760>=0)?1:0;

ninexnine_unit ninexnine_unit_420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10770)
);

ninexnine_unit ninexnine_unit_421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11770)
);

ninexnine_unit ninexnine_unit_422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12770)
);

ninexnine_unit ninexnine_unit_423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13770)
);

assign C1770=c10770+c11770+c12770+c13770;
assign A1770=(C1770>=0)?1:0;

ninexnine_unit ninexnine_unit_424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10780)
);

ninexnine_unit ninexnine_unit_425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11780)
);

ninexnine_unit ninexnine_unit_426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12780)
);

ninexnine_unit ninexnine_unit_427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13780)
);

assign C1780=c10780+c11780+c12780+c13780;
assign A1780=(C1780>=0)?1:0;

ninexnine_unit ninexnine_unit_428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10790)
);

ninexnine_unit ninexnine_unit_429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11790)
);

ninexnine_unit ninexnine_unit_430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12790)
);

ninexnine_unit ninexnine_unit_431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13790)
);

assign C1790=c10790+c11790+c12790+c13790;
assign A1790=(C1790>=0)?1:0;

ninexnine_unit ninexnine_unit_432(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c107A0)
);

ninexnine_unit ninexnine_unit_433(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c117A0)
);

ninexnine_unit ninexnine_unit_434(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c127A0)
);

ninexnine_unit ninexnine_unit_435(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c137A0)
);

assign C17A0=c107A0+c117A0+c127A0+c137A0;
assign A17A0=(C17A0>=0)?1:0;

ninexnine_unit ninexnine_unit_436(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c107B0)
);

ninexnine_unit ninexnine_unit_437(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c117B0)
);

ninexnine_unit ninexnine_unit_438(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c127B0)
);

ninexnine_unit ninexnine_unit_439(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c137B0)
);

assign C17B0=c107B0+c117B0+c127B0+c137B0;
assign A17B0=(C17B0>=0)?1:0;

ninexnine_unit ninexnine_unit_440(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c107C0)
);

ninexnine_unit ninexnine_unit_441(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c117C0)
);

ninexnine_unit ninexnine_unit_442(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c127C0)
);

ninexnine_unit ninexnine_unit_443(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c137C0)
);

assign C17C0=c107C0+c117C0+c127C0+c137C0;
assign A17C0=(C17C0>=0)?1:0;

ninexnine_unit ninexnine_unit_444(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c107D0)
);

ninexnine_unit ninexnine_unit_445(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c117D0)
);

ninexnine_unit ninexnine_unit_446(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c127D0)
);

ninexnine_unit ninexnine_unit_447(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c137D0)
);

assign C17D0=c107D0+c117D0+c127D0+c137D0;
assign A17D0=(C17D0>=0)?1:0;

ninexnine_unit ninexnine_unit_448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10800)
);

ninexnine_unit ninexnine_unit_449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11800)
);

ninexnine_unit ninexnine_unit_450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12800)
);

ninexnine_unit ninexnine_unit_451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13800)
);

assign C1800=c10800+c11800+c12800+c13800;
assign A1800=(C1800>=0)?1:0;

ninexnine_unit ninexnine_unit_452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10810)
);

ninexnine_unit ninexnine_unit_453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11810)
);

ninexnine_unit ninexnine_unit_454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12810)
);

ninexnine_unit ninexnine_unit_455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13810)
);

assign C1810=c10810+c11810+c12810+c13810;
assign A1810=(C1810>=0)?1:0;

ninexnine_unit ninexnine_unit_456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10820)
);

ninexnine_unit ninexnine_unit_457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11820)
);

ninexnine_unit ninexnine_unit_458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12820)
);

ninexnine_unit ninexnine_unit_459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13820)
);

assign C1820=c10820+c11820+c12820+c13820;
assign A1820=(C1820>=0)?1:0;

ninexnine_unit ninexnine_unit_460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10830)
);

ninexnine_unit ninexnine_unit_461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11830)
);

ninexnine_unit ninexnine_unit_462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12830)
);

ninexnine_unit ninexnine_unit_463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13830)
);

assign C1830=c10830+c11830+c12830+c13830;
assign A1830=(C1830>=0)?1:0;

ninexnine_unit ninexnine_unit_464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10840)
);

ninexnine_unit ninexnine_unit_465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11840)
);

ninexnine_unit ninexnine_unit_466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12840)
);

ninexnine_unit ninexnine_unit_467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13840)
);

assign C1840=c10840+c11840+c12840+c13840;
assign A1840=(C1840>=0)?1:0;

ninexnine_unit ninexnine_unit_468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10850)
);

ninexnine_unit ninexnine_unit_469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11850)
);

ninexnine_unit ninexnine_unit_470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12850)
);

ninexnine_unit ninexnine_unit_471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13850)
);

assign C1850=c10850+c11850+c12850+c13850;
assign A1850=(C1850>=0)?1:0;

ninexnine_unit ninexnine_unit_472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10860)
);

ninexnine_unit ninexnine_unit_473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11860)
);

ninexnine_unit ninexnine_unit_474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12860)
);

ninexnine_unit ninexnine_unit_475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13860)
);

assign C1860=c10860+c11860+c12860+c13860;
assign A1860=(C1860>=0)?1:0;

ninexnine_unit ninexnine_unit_476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10870)
);

ninexnine_unit ninexnine_unit_477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11870)
);

ninexnine_unit ninexnine_unit_478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12870)
);

ninexnine_unit ninexnine_unit_479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13870)
);

assign C1870=c10870+c11870+c12870+c13870;
assign A1870=(C1870>=0)?1:0;

ninexnine_unit ninexnine_unit_480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10880)
);

ninexnine_unit ninexnine_unit_481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11880)
);

ninexnine_unit ninexnine_unit_482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12880)
);

ninexnine_unit ninexnine_unit_483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13880)
);

assign C1880=c10880+c11880+c12880+c13880;
assign A1880=(C1880>=0)?1:0;

ninexnine_unit ninexnine_unit_484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10890)
);

ninexnine_unit ninexnine_unit_485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11890)
);

ninexnine_unit ninexnine_unit_486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12890)
);

ninexnine_unit ninexnine_unit_487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13890)
);

assign C1890=c10890+c11890+c12890+c13890;
assign A1890=(C1890>=0)?1:0;

ninexnine_unit ninexnine_unit_488(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c108A0)
);

ninexnine_unit ninexnine_unit_489(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c118A0)
);

ninexnine_unit ninexnine_unit_490(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c128A0)
);

ninexnine_unit ninexnine_unit_491(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c138A0)
);

assign C18A0=c108A0+c118A0+c128A0+c138A0;
assign A18A0=(C18A0>=0)?1:0;

ninexnine_unit ninexnine_unit_492(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c108B0)
);

ninexnine_unit ninexnine_unit_493(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c118B0)
);

ninexnine_unit ninexnine_unit_494(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c128B0)
);

ninexnine_unit ninexnine_unit_495(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c138B0)
);

assign C18B0=c108B0+c118B0+c128B0+c138B0;
assign A18B0=(C18B0>=0)?1:0;

ninexnine_unit ninexnine_unit_496(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c108C0)
);

ninexnine_unit ninexnine_unit_497(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c118C0)
);

ninexnine_unit ninexnine_unit_498(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c128C0)
);

ninexnine_unit ninexnine_unit_499(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c138C0)
);

assign C18C0=c108C0+c118C0+c128C0+c138C0;
assign A18C0=(C18C0>=0)?1:0;

ninexnine_unit ninexnine_unit_500(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c108D0)
);

ninexnine_unit ninexnine_unit_501(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c118D0)
);

ninexnine_unit ninexnine_unit_502(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c128D0)
);

ninexnine_unit ninexnine_unit_503(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c138D0)
);

assign C18D0=c108D0+c118D0+c128D0+c138D0;
assign A18D0=(C18D0>=0)?1:0;

ninexnine_unit ninexnine_unit_504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10900)
);

ninexnine_unit ninexnine_unit_505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11900)
);

ninexnine_unit ninexnine_unit_506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12900)
);

ninexnine_unit ninexnine_unit_507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13900)
);

assign C1900=c10900+c11900+c12900+c13900;
assign A1900=(C1900>=0)?1:0;

ninexnine_unit ninexnine_unit_508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10910)
);

ninexnine_unit ninexnine_unit_509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11910)
);

ninexnine_unit ninexnine_unit_510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12910)
);

ninexnine_unit ninexnine_unit_511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13910)
);

assign C1910=c10910+c11910+c12910+c13910;
assign A1910=(C1910>=0)?1:0;

ninexnine_unit ninexnine_unit_512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10920)
);

ninexnine_unit ninexnine_unit_513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11920)
);

ninexnine_unit ninexnine_unit_514(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12920)
);

ninexnine_unit ninexnine_unit_515(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13920)
);

assign C1920=c10920+c11920+c12920+c13920;
assign A1920=(C1920>=0)?1:0;

ninexnine_unit ninexnine_unit_516(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10930)
);

ninexnine_unit ninexnine_unit_517(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11930)
);

ninexnine_unit ninexnine_unit_518(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12930)
);

ninexnine_unit ninexnine_unit_519(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13930)
);

assign C1930=c10930+c11930+c12930+c13930;
assign A1930=(C1930>=0)?1:0;

ninexnine_unit ninexnine_unit_520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10940)
);

ninexnine_unit ninexnine_unit_521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11940)
);

ninexnine_unit ninexnine_unit_522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12940)
);

ninexnine_unit ninexnine_unit_523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13940)
);

assign C1940=c10940+c11940+c12940+c13940;
assign A1940=(C1940>=0)?1:0;

ninexnine_unit ninexnine_unit_524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10950)
);

ninexnine_unit ninexnine_unit_525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11950)
);

ninexnine_unit ninexnine_unit_526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12950)
);

ninexnine_unit ninexnine_unit_527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13950)
);

assign C1950=c10950+c11950+c12950+c13950;
assign A1950=(C1950>=0)?1:0;

ninexnine_unit ninexnine_unit_528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10960)
);

ninexnine_unit ninexnine_unit_529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11960)
);

ninexnine_unit ninexnine_unit_530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12960)
);

ninexnine_unit ninexnine_unit_531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13960)
);

assign C1960=c10960+c11960+c12960+c13960;
assign A1960=(C1960>=0)?1:0;

ninexnine_unit ninexnine_unit_532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10970)
);

ninexnine_unit ninexnine_unit_533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11970)
);

ninexnine_unit ninexnine_unit_534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12970)
);

ninexnine_unit ninexnine_unit_535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13970)
);

assign C1970=c10970+c11970+c12970+c13970;
assign A1970=(C1970>=0)?1:0;

ninexnine_unit ninexnine_unit_536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10980)
);

ninexnine_unit ninexnine_unit_537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11980)
);

ninexnine_unit ninexnine_unit_538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12980)
);

ninexnine_unit ninexnine_unit_539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13980)
);

assign C1980=c10980+c11980+c12980+c13980;
assign A1980=(C1980>=0)?1:0;

ninexnine_unit ninexnine_unit_540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10990)
);

ninexnine_unit ninexnine_unit_541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11990)
);

ninexnine_unit ninexnine_unit_542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12990)
);

ninexnine_unit ninexnine_unit_543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13990)
);

assign C1990=c10990+c11990+c12990+c13990;
assign A1990=(C1990>=0)?1:0;

ninexnine_unit ninexnine_unit_544(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c109A0)
);

ninexnine_unit ninexnine_unit_545(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c119A0)
);

ninexnine_unit ninexnine_unit_546(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c129A0)
);

ninexnine_unit ninexnine_unit_547(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c139A0)
);

assign C19A0=c109A0+c119A0+c129A0+c139A0;
assign A19A0=(C19A0>=0)?1:0;

ninexnine_unit ninexnine_unit_548(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c109B0)
);

ninexnine_unit ninexnine_unit_549(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c119B0)
);

ninexnine_unit ninexnine_unit_550(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c129B0)
);

ninexnine_unit ninexnine_unit_551(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c139B0)
);

assign C19B0=c109B0+c119B0+c129B0+c139B0;
assign A19B0=(C19B0>=0)?1:0;

ninexnine_unit ninexnine_unit_552(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c109C0)
);

ninexnine_unit ninexnine_unit_553(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c119C0)
);

ninexnine_unit ninexnine_unit_554(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c129C0)
);

ninexnine_unit ninexnine_unit_555(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c139C0)
);

assign C19C0=c109C0+c119C0+c129C0+c139C0;
assign A19C0=(C19C0>=0)?1:0;

ninexnine_unit ninexnine_unit_556(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c109D0)
);

ninexnine_unit ninexnine_unit_557(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c119D0)
);

ninexnine_unit ninexnine_unit_558(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c129D0)
);

ninexnine_unit ninexnine_unit_559(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c139D0)
);

assign C19D0=c109D0+c119D0+c129D0+c139D0;
assign A19D0=(C19D0>=0)?1:0;

ninexnine_unit ninexnine_unit_560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A00)
);

ninexnine_unit ninexnine_unit_561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A00)
);

ninexnine_unit ninexnine_unit_562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A00)
);

ninexnine_unit ninexnine_unit_563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A00)
);

assign C1A00=c10A00+c11A00+c12A00+c13A00;
assign A1A00=(C1A00>=0)?1:0;

ninexnine_unit ninexnine_unit_564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A10)
);

ninexnine_unit ninexnine_unit_565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A10)
);

ninexnine_unit ninexnine_unit_566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A10)
);

ninexnine_unit ninexnine_unit_567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A10)
);

assign C1A10=c10A10+c11A10+c12A10+c13A10;
assign A1A10=(C1A10>=0)?1:0;

ninexnine_unit ninexnine_unit_568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A20)
);

ninexnine_unit ninexnine_unit_569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A20)
);

ninexnine_unit ninexnine_unit_570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A20)
);

ninexnine_unit ninexnine_unit_571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A20)
);

assign C1A20=c10A20+c11A20+c12A20+c13A20;
assign A1A20=(C1A20>=0)?1:0;

ninexnine_unit ninexnine_unit_572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A30)
);

ninexnine_unit ninexnine_unit_573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A30)
);

ninexnine_unit ninexnine_unit_574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A30)
);

ninexnine_unit ninexnine_unit_575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A30)
);

assign C1A30=c10A30+c11A30+c12A30+c13A30;
assign A1A30=(C1A30>=0)?1:0;

ninexnine_unit ninexnine_unit_576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A40)
);

ninexnine_unit ninexnine_unit_577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A40)
);

ninexnine_unit ninexnine_unit_578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A40)
);

ninexnine_unit ninexnine_unit_579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A40)
);

assign C1A40=c10A40+c11A40+c12A40+c13A40;
assign A1A40=(C1A40>=0)?1:0;

ninexnine_unit ninexnine_unit_580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A50)
);

ninexnine_unit ninexnine_unit_581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A50)
);

ninexnine_unit ninexnine_unit_582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A50)
);

ninexnine_unit ninexnine_unit_583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A50)
);

assign C1A50=c10A50+c11A50+c12A50+c13A50;
assign A1A50=(C1A50>=0)?1:0;

ninexnine_unit ninexnine_unit_584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A60)
);

ninexnine_unit ninexnine_unit_585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A60)
);

ninexnine_unit ninexnine_unit_586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A60)
);

ninexnine_unit ninexnine_unit_587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A60)
);

assign C1A60=c10A60+c11A60+c12A60+c13A60;
assign A1A60=(C1A60>=0)?1:0;

ninexnine_unit ninexnine_unit_588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A70)
);

ninexnine_unit ninexnine_unit_589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A70)
);

ninexnine_unit ninexnine_unit_590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A70)
);

ninexnine_unit ninexnine_unit_591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A70)
);

assign C1A70=c10A70+c11A70+c12A70+c13A70;
assign A1A70=(C1A70>=0)?1:0;

ninexnine_unit ninexnine_unit_592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A80)
);

ninexnine_unit ninexnine_unit_593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A80)
);

ninexnine_unit ninexnine_unit_594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A80)
);

ninexnine_unit ninexnine_unit_595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A80)
);

assign C1A80=c10A80+c11A80+c12A80+c13A80;
assign A1A80=(C1A80>=0)?1:0;

ninexnine_unit ninexnine_unit_596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10A90)
);

ninexnine_unit ninexnine_unit_597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11A90)
);

ninexnine_unit ninexnine_unit_598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12A90)
);

ninexnine_unit ninexnine_unit_599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13A90)
);

assign C1A90=c10A90+c11A90+c12A90+c13A90;
assign A1A90=(C1A90>=0)?1:0;

ninexnine_unit ninexnine_unit_600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10AA0)
);

ninexnine_unit ninexnine_unit_601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11AA0)
);

ninexnine_unit ninexnine_unit_602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12AA0)
);

ninexnine_unit ninexnine_unit_603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13AA0)
);

assign C1AA0=c10AA0+c11AA0+c12AA0+c13AA0;
assign A1AA0=(C1AA0>=0)?1:0;

ninexnine_unit ninexnine_unit_604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10AB0)
);

ninexnine_unit ninexnine_unit_605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11AB0)
);

ninexnine_unit ninexnine_unit_606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12AB0)
);

ninexnine_unit ninexnine_unit_607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13AB0)
);

assign C1AB0=c10AB0+c11AB0+c12AB0+c13AB0;
assign A1AB0=(C1AB0>=0)?1:0;

ninexnine_unit ninexnine_unit_608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10AC0)
);

ninexnine_unit ninexnine_unit_609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11AC0)
);

ninexnine_unit ninexnine_unit_610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12AC0)
);

ninexnine_unit ninexnine_unit_611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13AC0)
);

assign C1AC0=c10AC0+c11AC0+c12AC0+c13AC0;
assign A1AC0=(C1AC0>=0)?1:0;

ninexnine_unit ninexnine_unit_612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10AD0)
);

ninexnine_unit ninexnine_unit_613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11AD0)
);

ninexnine_unit ninexnine_unit_614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12AD0)
);

ninexnine_unit ninexnine_unit_615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13AD0)
);

assign C1AD0=c10AD0+c11AD0+c12AD0+c13AD0;
assign A1AD0=(C1AD0>=0)?1:0;

ninexnine_unit ninexnine_unit_616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B00)
);

ninexnine_unit ninexnine_unit_617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B00)
);

ninexnine_unit ninexnine_unit_618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B00)
);

ninexnine_unit ninexnine_unit_619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B00)
);

assign C1B00=c10B00+c11B00+c12B00+c13B00;
assign A1B00=(C1B00>=0)?1:0;

ninexnine_unit ninexnine_unit_620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B10)
);

ninexnine_unit ninexnine_unit_621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B10)
);

ninexnine_unit ninexnine_unit_622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B10)
);

ninexnine_unit ninexnine_unit_623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B10)
);

assign C1B10=c10B10+c11B10+c12B10+c13B10;
assign A1B10=(C1B10>=0)?1:0;

ninexnine_unit ninexnine_unit_624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B20)
);

ninexnine_unit ninexnine_unit_625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B20)
);

ninexnine_unit ninexnine_unit_626(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B20)
);

ninexnine_unit ninexnine_unit_627(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B20)
);

assign C1B20=c10B20+c11B20+c12B20+c13B20;
assign A1B20=(C1B20>=0)?1:0;

ninexnine_unit ninexnine_unit_628(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B30)
);

ninexnine_unit ninexnine_unit_629(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B30)
);

ninexnine_unit ninexnine_unit_630(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B30)
);

ninexnine_unit ninexnine_unit_631(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B30)
);

assign C1B30=c10B30+c11B30+c12B30+c13B30;
assign A1B30=(C1B30>=0)?1:0;

ninexnine_unit ninexnine_unit_632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B40)
);

ninexnine_unit ninexnine_unit_633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B40)
);

ninexnine_unit ninexnine_unit_634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B40)
);

ninexnine_unit ninexnine_unit_635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B40)
);

assign C1B40=c10B40+c11B40+c12B40+c13B40;
assign A1B40=(C1B40>=0)?1:0;

ninexnine_unit ninexnine_unit_636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B50)
);

ninexnine_unit ninexnine_unit_637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B50)
);

ninexnine_unit ninexnine_unit_638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B50)
);

ninexnine_unit ninexnine_unit_639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B50)
);

assign C1B50=c10B50+c11B50+c12B50+c13B50;
assign A1B50=(C1B50>=0)?1:0;

ninexnine_unit ninexnine_unit_640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B60)
);

ninexnine_unit ninexnine_unit_641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B60)
);

ninexnine_unit ninexnine_unit_642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B60)
);

ninexnine_unit ninexnine_unit_643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B60)
);

assign C1B60=c10B60+c11B60+c12B60+c13B60;
assign A1B60=(C1B60>=0)?1:0;

ninexnine_unit ninexnine_unit_644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B70)
);

ninexnine_unit ninexnine_unit_645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B70)
);

ninexnine_unit ninexnine_unit_646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B70)
);

ninexnine_unit ninexnine_unit_647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B70)
);

assign C1B70=c10B70+c11B70+c12B70+c13B70;
assign A1B70=(C1B70>=0)?1:0;

ninexnine_unit ninexnine_unit_648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B80)
);

ninexnine_unit ninexnine_unit_649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B80)
);

ninexnine_unit ninexnine_unit_650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B80)
);

ninexnine_unit ninexnine_unit_651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B80)
);

assign C1B80=c10B80+c11B80+c12B80+c13B80;
assign A1B80=(C1B80>=0)?1:0;

ninexnine_unit ninexnine_unit_652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10B90)
);

ninexnine_unit ninexnine_unit_653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11B90)
);

ninexnine_unit ninexnine_unit_654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12B90)
);

ninexnine_unit ninexnine_unit_655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13B90)
);

assign C1B90=c10B90+c11B90+c12B90+c13B90;
assign A1B90=(C1B90>=0)?1:0;

ninexnine_unit ninexnine_unit_656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10BA0)
);

ninexnine_unit ninexnine_unit_657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11BA0)
);

ninexnine_unit ninexnine_unit_658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12BA0)
);

ninexnine_unit ninexnine_unit_659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13BA0)
);

assign C1BA0=c10BA0+c11BA0+c12BA0+c13BA0;
assign A1BA0=(C1BA0>=0)?1:0;

ninexnine_unit ninexnine_unit_660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10BB0)
);

ninexnine_unit ninexnine_unit_661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11BB0)
);

ninexnine_unit ninexnine_unit_662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12BB0)
);

ninexnine_unit ninexnine_unit_663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13BB0)
);

assign C1BB0=c10BB0+c11BB0+c12BB0+c13BB0;
assign A1BB0=(C1BB0>=0)?1:0;

ninexnine_unit ninexnine_unit_664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10BC0)
);

ninexnine_unit ninexnine_unit_665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11BC0)
);

ninexnine_unit ninexnine_unit_666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12BC0)
);

ninexnine_unit ninexnine_unit_667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13BC0)
);

assign C1BC0=c10BC0+c11BC0+c12BC0+c13BC0;
assign A1BC0=(C1BC0>=0)?1:0;

ninexnine_unit ninexnine_unit_668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10BD0)
);

ninexnine_unit ninexnine_unit_669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11BD0)
);

ninexnine_unit ninexnine_unit_670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12BD0)
);

ninexnine_unit ninexnine_unit_671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13BD0)
);

assign C1BD0=c10BD0+c11BD0+c12BD0+c13BD0;
assign A1BD0=(C1BD0>=0)?1:0;

ninexnine_unit ninexnine_unit_672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C00)
);

ninexnine_unit ninexnine_unit_673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C00)
);

ninexnine_unit ninexnine_unit_674(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C00)
);

ninexnine_unit ninexnine_unit_675(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C00)
);

assign C1C00=c10C00+c11C00+c12C00+c13C00;
assign A1C00=(C1C00>=0)?1:0;

ninexnine_unit ninexnine_unit_676(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C10)
);

ninexnine_unit ninexnine_unit_677(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C10)
);

ninexnine_unit ninexnine_unit_678(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C10)
);

ninexnine_unit ninexnine_unit_679(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C10)
);

assign C1C10=c10C10+c11C10+c12C10+c13C10;
assign A1C10=(C1C10>=0)?1:0;

ninexnine_unit ninexnine_unit_680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C20)
);

ninexnine_unit ninexnine_unit_681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C20)
);

ninexnine_unit ninexnine_unit_682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C20)
);

ninexnine_unit ninexnine_unit_683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C20)
);

assign C1C20=c10C20+c11C20+c12C20+c13C20;
assign A1C20=(C1C20>=0)?1:0;

ninexnine_unit ninexnine_unit_684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C30)
);

ninexnine_unit ninexnine_unit_685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C30)
);

ninexnine_unit ninexnine_unit_686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C30)
);

ninexnine_unit ninexnine_unit_687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C30)
);

assign C1C30=c10C30+c11C30+c12C30+c13C30;
assign A1C30=(C1C30>=0)?1:0;

ninexnine_unit ninexnine_unit_688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C40)
);

ninexnine_unit ninexnine_unit_689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C40)
);

ninexnine_unit ninexnine_unit_690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C40)
);

ninexnine_unit ninexnine_unit_691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C40)
);

assign C1C40=c10C40+c11C40+c12C40+c13C40;
assign A1C40=(C1C40>=0)?1:0;

ninexnine_unit ninexnine_unit_692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C50)
);

ninexnine_unit ninexnine_unit_693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C50)
);

ninexnine_unit ninexnine_unit_694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C50)
);

ninexnine_unit ninexnine_unit_695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C50)
);

assign C1C50=c10C50+c11C50+c12C50+c13C50;
assign A1C50=(C1C50>=0)?1:0;

ninexnine_unit ninexnine_unit_696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C60)
);

ninexnine_unit ninexnine_unit_697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C60)
);

ninexnine_unit ninexnine_unit_698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C60)
);

ninexnine_unit ninexnine_unit_699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C60)
);

assign C1C60=c10C60+c11C60+c12C60+c13C60;
assign A1C60=(C1C60>=0)?1:0;

ninexnine_unit ninexnine_unit_700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C70)
);

ninexnine_unit ninexnine_unit_701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C70)
);

ninexnine_unit ninexnine_unit_702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C70)
);

ninexnine_unit ninexnine_unit_703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C70)
);

assign C1C70=c10C70+c11C70+c12C70+c13C70;
assign A1C70=(C1C70>=0)?1:0;

ninexnine_unit ninexnine_unit_704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C80)
);

ninexnine_unit ninexnine_unit_705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C80)
);

ninexnine_unit ninexnine_unit_706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C80)
);

ninexnine_unit ninexnine_unit_707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C80)
);

assign C1C80=c10C80+c11C80+c12C80+c13C80;
assign A1C80=(C1C80>=0)?1:0;

ninexnine_unit ninexnine_unit_708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10C90)
);

ninexnine_unit ninexnine_unit_709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11C90)
);

ninexnine_unit ninexnine_unit_710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12C90)
);

ninexnine_unit ninexnine_unit_711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13C90)
);

assign C1C90=c10C90+c11C90+c12C90+c13C90;
assign A1C90=(C1C90>=0)?1:0;

ninexnine_unit ninexnine_unit_712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10CA0)
);

ninexnine_unit ninexnine_unit_713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11CA0)
);

ninexnine_unit ninexnine_unit_714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12CA0)
);

ninexnine_unit ninexnine_unit_715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13CA0)
);

assign C1CA0=c10CA0+c11CA0+c12CA0+c13CA0;
assign A1CA0=(C1CA0>=0)?1:0;

ninexnine_unit ninexnine_unit_716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10CB0)
);

ninexnine_unit ninexnine_unit_717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11CB0)
);

ninexnine_unit ninexnine_unit_718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12CB0)
);

ninexnine_unit ninexnine_unit_719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13CB0)
);

assign C1CB0=c10CB0+c11CB0+c12CB0+c13CB0;
assign A1CB0=(C1CB0>=0)?1:0;

ninexnine_unit ninexnine_unit_720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10CC0)
);

ninexnine_unit ninexnine_unit_721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11CC0)
);

ninexnine_unit ninexnine_unit_722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12CC0)
);

ninexnine_unit ninexnine_unit_723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13CC0)
);

assign C1CC0=c10CC0+c11CC0+c12CC0+c13CC0;
assign A1CC0=(C1CC0>=0)?1:0;

ninexnine_unit ninexnine_unit_724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10CD0)
);

ninexnine_unit ninexnine_unit_725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11CD0)
);

ninexnine_unit ninexnine_unit_726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12CD0)
);

ninexnine_unit ninexnine_unit_727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13CD0)
);

assign C1CD0=c10CD0+c11CD0+c12CD0+c13CD0;
assign A1CD0=(C1CD0>=0)?1:0;

ninexnine_unit ninexnine_unit_728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D00)
);

ninexnine_unit ninexnine_unit_729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D00)
);

ninexnine_unit ninexnine_unit_730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D00)
);

ninexnine_unit ninexnine_unit_731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D00)
);

assign C1D00=c10D00+c11D00+c12D00+c13D00;
assign A1D00=(C1D00>=0)?1:0;

ninexnine_unit ninexnine_unit_732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D10)
);

ninexnine_unit ninexnine_unit_733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D10)
);

ninexnine_unit ninexnine_unit_734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D10)
);

ninexnine_unit ninexnine_unit_735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D10)
);

assign C1D10=c10D10+c11D10+c12D10+c13D10;
assign A1D10=(C1D10>=0)?1:0;

ninexnine_unit ninexnine_unit_736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D20)
);

ninexnine_unit ninexnine_unit_737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D20)
);

ninexnine_unit ninexnine_unit_738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D20)
);

ninexnine_unit ninexnine_unit_739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D20)
);

assign C1D20=c10D20+c11D20+c12D20+c13D20;
assign A1D20=(C1D20>=0)?1:0;

ninexnine_unit ninexnine_unit_740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D30)
);

ninexnine_unit ninexnine_unit_741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D30)
);

ninexnine_unit ninexnine_unit_742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D30)
);

ninexnine_unit ninexnine_unit_743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D30)
);

assign C1D30=c10D30+c11D30+c12D30+c13D30;
assign A1D30=(C1D30>=0)?1:0;

ninexnine_unit ninexnine_unit_744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D40)
);

ninexnine_unit ninexnine_unit_745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D40)
);

ninexnine_unit ninexnine_unit_746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D40)
);

ninexnine_unit ninexnine_unit_747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D40)
);

assign C1D40=c10D40+c11D40+c12D40+c13D40;
assign A1D40=(C1D40>=0)?1:0;

ninexnine_unit ninexnine_unit_748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D50)
);

ninexnine_unit ninexnine_unit_749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D50)
);

ninexnine_unit ninexnine_unit_750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D50)
);

ninexnine_unit ninexnine_unit_751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D50)
);

assign C1D50=c10D50+c11D50+c12D50+c13D50;
assign A1D50=(C1D50>=0)?1:0;

ninexnine_unit ninexnine_unit_752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D60)
);

ninexnine_unit ninexnine_unit_753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D60)
);

ninexnine_unit ninexnine_unit_754(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D60)
);

ninexnine_unit ninexnine_unit_755(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D60)
);

assign C1D60=c10D60+c11D60+c12D60+c13D60;
assign A1D60=(C1D60>=0)?1:0;

ninexnine_unit ninexnine_unit_756(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D70)
);

ninexnine_unit ninexnine_unit_757(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D70)
);

ninexnine_unit ninexnine_unit_758(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D70)
);

ninexnine_unit ninexnine_unit_759(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D70)
);

assign C1D70=c10D70+c11D70+c12D70+c13D70;
assign A1D70=(C1D70>=0)?1:0;

ninexnine_unit ninexnine_unit_760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D80)
);

ninexnine_unit ninexnine_unit_761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D80)
);

ninexnine_unit ninexnine_unit_762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D80)
);

ninexnine_unit ninexnine_unit_763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D80)
);

assign C1D80=c10D80+c11D80+c12D80+c13D80;
assign A1D80=(C1D80>=0)?1:0;

ninexnine_unit ninexnine_unit_764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10D90)
);

ninexnine_unit ninexnine_unit_765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11D90)
);

ninexnine_unit ninexnine_unit_766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12D90)
);

ninexnine_unit ninexnine_unit_767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13D90)
);

assign C1D90=c10D90+c11D90+c12D90+c13D90;
assign A1D90=(C1D90>=0)?1:0;

ninexnine_unit ninexnine_unit_768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10DA0)
);

ninexnine_unit ninexnine_unit_769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11DA0)
);

ninexnine_unit ninexnine_unit_770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12DA0)
);

ninexnine_unit ninexnine_unit_771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13DA0)
);

assign C1DA0=c10DA0+c11DA0+c12DA0+c13DA0;
assign A1DA0=(C1DA0>=0)?1:0;

ninexnine_unit ninexnine_unit_772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10DB0)
);

ninexnine_unit ninexnine_unit_773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11DB0)
);

ninexnine_unit ninexnine_unit_774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12DB0)
);

ninexnine_unit ninexnine_unit_775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13DB0)
);

assign C1DB0=c10DB0+c11DB0+c12DB0+c13DB0;
assign A1DB0=(C1DB0>=0)?1:0;

ninexnine_unit ninexnine_unit_776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10DC0)
);

ninexnine_unit ninexnine_unit_777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11DC0)
);

ninexnine_unit ninexnine_unit_778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12DC0)
);

ninexnine_unit ninexnine_unit_779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13DC0)
);

assign C1DC0=c10DC0+c11DC0+c12DC0+c13DC0;
assign A1DC0=(C1DC0>=0)?1:0;

ninexnine_unit ninexnine_unit_780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10DD0)
);

ninexnine_unit ninexnine_unit_781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11DD0)
);

ninexnine_unit ninexnine_unit_782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12DD0)
);

ninexnine_unit ninexnine_unit_783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13DD0)
);

assign C1DD0=c10DD0+c11DD0+c12DD0+c13DD0;
assign A1DD0=(C1DD0>=0)?1:0;

ninexnine_unit ninexnine_unit_784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10001)
);

ninexnine_unit ninexnine_unit_785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11001)
);

ninexnine_unit ninexnine_unit_786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12001)
);

ninexnine_unit ninexnine_unit_787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13001)
);

assign C1001=c10001+c11001+c12001+c13001;
assign A1001=(C1001>=0)?1:0;

ninexnine_unit ninexnine_unit_788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10011)
);

ninexnine_unit ninexnine_unit_789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11011)
);

ninexnine_unit ninexnine_unit_790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12011)
);

ninexnine_unit ninexnine_unit_791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13011)
);

assign C1011=c10011+c11011+c12011+c13011;
assign A1011=(C1011>=0)?1:0;

ninexnine_unit ninexnine_unit_792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10021)
);

ninexnine_unit ninexnine_unit_793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11021)
);

ninexnine_unit ninexnine_unit_794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12021)
);

ninexnine_unit ninexnine_unit_795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13021)
);

assign C1021=c10021+c11021+c12021+c13021;
assign A1021=(C1021>=0)?1:0;

ninexnine_unit ninexnine_unit_796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10031)
);

ninexnine_unit ninexnine_unit_797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11031)
);

ninexnine_unit ninexnine_unit_798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12031)
);

ninexnine_unit ninexnine_unit_799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13031)
);

assign C1031=c10031+c11031+c12031+c13031;
assign A1031=(C1031>=0)?1:0;

ninexnine_unit ninexnine_unit_800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10041)
);

ninexnine_unit ninexnine_unit_801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11041)
);

ninexnine_unit ninexnine_unit_802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12041)
);

ninexnine_unit ninexnine_unit_803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13041)
);

assign C1041=c10041+c11041+c12041+c13041;
assign A1041=(C1041>=0)?1:0;

ninexnine_unit ninexnine_unit_804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10051)
);

ninexnine_unit ninexnine_unit_805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11051)
);

ninexnine_unit ninexnine_unit_806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12051)
);

ninexnine_unit ninexnine_unit_807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13051)
);

assign C1051=c10051+c11051+c12051+c13051;
assign A1051=(C1051>=0)?1:0;

ninexnine_unit ninexnine_unit_808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10061)
);

ninexnine_unit ninexnine_unit_809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11061)
);

ninexnine_unit ninexnine_unit_810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12061)
);

ninexnine_unit ninexnine_unit_811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13061)
);

assign C1061=c10061+c11061+c12061+c13061;
assign A1061=(C1061>=0)?1:0;

ninexnine_unit ninexnine_unit_812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10071)
);

ninexnine_unit ninexnine_unit_813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11071)
);

ninexnine_unit ninexnine_unit_814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12071)
);

ninexnine_unit ninexnine_unit_815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13071)
);

assign C1071=c10071+c11071+c12071+c13071;
assign A1071=(C1071>=0)?1:0;

ninexnine_unit ninexnine_unit_816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10081)
);

ninexnine_unit ninexnine_unit_817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11081)
);

ninexnine_unit ninexnine_unit_818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12081)
);

ninexnine_unit ninexnine_unit_819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13081)
);

assign C1081=c10081+c11081+c12081+c13081;
assign A1081=(C1081>=0)?1:0;

ninexnine_unit ninexnine_unit_820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10091)
);

ninexnine_unit ninexnine_unit_821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11091)
);

ninexnine_unit ninexnine_unit_822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12091)
);

ninexnine_unit ninexnine_unit_823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13091)
);

assign C1091=c10091+c11091+c12091+c13091;
assign A1091=(C1091>=0)?1:0;

ninexnine_unit ninexnine_unit_824(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c100A1)
);

ninexnine_unit ninexnine_unit_825(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c110A1)
);

ninexnine_unit ninexnine_unit_826(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c120A1)
);

ninexnine_unit ninexnine_unit_827(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c130A1)
);

assign C10A1=c100A1+c110A1+c120A1+c130A1;
assign A10A1=(C10A1>=0)?1:0;

ninexnine_unit ninexnine_unit_828(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c100B1)
);

ninexnine_unit ninexnine_unit_829(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c110B1)
);

ninexnine_unit ninexnine_unit_830(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c120B1)
);

ninexnine_unit ninexnine_unit_831(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c130B1)
);

assign C10B1=c100B1+c110B1+c120B1+c130B1;
assign A10B1=(C10B1>=0)?1:0;

ninexnine_unit ninexnine_unit_832(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c100C1)
);

ninexnine_unit ninexnine_unit_833(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c110C1)
);

ninexnine_unit ninexnine_unit_834(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c120C1)
);

ninexnine_unit ninexnine_unit_835(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c130C1)
);

assign C10C1=c100C1+c110C1+c120C1+c130C1;
assign A10C1=(C10C1>=0)?1:0;

ninexnine_unit ninexnine_unit_836(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c100D1)
);

ninexnine_unit ninexnine_unit_837(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c110D1)
);

ninexnine_unit ninexnine_unit_838(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c120D1)
);

ninexnine_unit ninexnine_unit_839(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c130D1)
);

assign C10D1=c100D1+c110D1+c120D1+c130D1;
assign A10D1=(C10D1>=0)?1:0;

ninexnine_unit ninexnine_unit_840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10101)
);

ninexnine_unit ninexnine_unit_841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11101)
);

ninexnine_unit ninexnine_unit_842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12101)
);

ninexnine_unit ninexnine_unit_843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13101)
);

assign C1101=c10101+c11101+c12101+c13101;
assign A1101=(C1101>=0)?1:0;

ninexnine_unit ninexnine_unit_844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10111)
);

ninexnine_unit ninexnine_unit_845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11111)
);

ninexnine_unit ninexnine_unit_846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12111)
);

ninexnine_unit ninexnine_unit_847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13111)
);

assign C1111=c10111+c11111+c12111+c13111;
assign A1111=(C1111>=0)?1:0;

ninexnine_unit ninexnine_unit_848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10121)
);

ninexnine_unit ninexnine_unit_849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11121)
);

ninexnine_unit ninexnine_unit_850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12121)
);

ninexnine_unit ninexnine_unit_851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13121)
);

assign C1121=c10121+c11121+c12121+c13121;
assign A1121=(C1121>=0)?1:0;

ninexnine_unit ninexnine_unit_852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10131)
);

ninexnine_unit ninexnine_unit_853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11131)
);

ninexnine_unit ninexnine_unit_854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12131)
);

ninexnine_unit ninexnine_unit_855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13131)
);

assign C1131=c10131+c11131+c12131+c13131;
assign A1131=(C1131>=0)?1:0;

ninexnine_unit ninexnine_unit_856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10141)
);

ninexnine_unit ninexnine_unit_857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11141)
);

ninexnine_unit ninexnine_unit_858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12141)
);

ninexnine_unit ninexnine_unit_859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13141)
);

assign C1141=c10141+c11141+c12141+c13141;
assign A1141=(C1141>=0)?1:0;

ninexnine_unit ninexnine_unit_860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10151)
);

ninexnine_unit ninexnine_unit_861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11151)
);

ninexnine_unit ninexnine_unit_862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12151)
);

ninexnine_unit ninexnine_unit_863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13151)
);

assign C1151=c10151+c11151+c12151+c13151;
assign A1151=(C1151>=0)?1:0;

ninexnine_unit ninexnine_unit_864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10161)
);

ninexnine_unit ninexnine_unit_865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11161)
);

ninexnine_unit ninexnine_unit_866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12161)
);

ninexnine_unit ninexnine_unit_867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13161)
);

assign C1161=c10161+c11161+c12161+c13161;
assign A1161=(C1161>=0)?1:0;

ninexnine_unit ninexnine_unit_868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10171)
);

ninexnine_unit ninexnine_unit_869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11171)
);

ninexnine_unit ninexnine_unit_870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12171)
);

ninexnine_unit ninexnine_unit_871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13171)
);

assign C1171=c10171+c11171+c12171+c13171;
assign A1171=(C1171>=0)?1:0;

ninexnine_unit ninexnine_unit_872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10181)
);

ninexnine_unit ninexnine_unit_873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11181)
);

ninexnine_unit ninexnine_unit_874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12181)
);

ninexnine_unit ninexnine_unit_875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13181)
);

assign C1181=c10181+c11181+c12181+c13181;
assign A1181=(C1181>=0)?1:0;

ninexnine_unit ninexnine_unit_876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10191)
);

ninexnine_unit ninexnine_unit_877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11191)
);

ninexnine_unit ninexnine_unit_878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12191)
);

ninexnine_unit ninexnine_unit_879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13191)
);

assign C1191=c10191+c11191+c12191+c13191;
assign A1191=(C1191>=0)?1:0;

ninexnine_unit ninexnine_unit_880(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c101A1)
);

ninexnine_unit ninexnine_unit_881(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c111A1)
);

ninexnine_unit ninexnine_unit_882(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c121A1)
);

ninexnine_unit ninexnine_unit_883(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c131A1)
);

assign C11A1=c101A1+c111A1+c121A1+c131A1;
assign A11A1=(C11A1>=0)?1:0;

ninexnine_unit ninexnine_unit_884(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c101B1)
);

ninexnine_unit ninexnine_unit_885(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c111B1)
);

ninexnine_unit ninexnine_unit_886(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c121B1)
);

ninexnine_unit ninexnine_unit_887(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c131B1)
);

assign C11B1=c101B1+c111B1+c121B1+c131B1;
assign A11B1=(C11B1>=0)?1:0;

ninexnine_unit ninexnine_unit_888(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c101C1)
);

ninexnine_unit ninexnine_unit_889(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c111C1)
);

ninexnine_unit ninexnine_unit_890(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c121C1)
);

ninexnine_unit ninexnine_unit_891(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c131C1)
);

assign C11C1=c101C1+c111C1+c121C1+c131C1;
assign A11C1=(C11C1>=0)?1:0;

ninexnine_unit ninexnine_unit_892(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c101D1)
);

ninexnine_unit ninexnine_unit_893(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c111D1)
);

ninexnine_unit ninexnine_unit_894(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c121D1)
);

ninexnine_unit ninexnine_unit_895(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c131D1)
);

assign C11D1=c101D1+c111D1+c121D1+c131D1;
assign A11D1=(C11D1>=0)?1:0;

ninexnine_unit ninexnine_unit_896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10201)
);

ninexnine_unit ninexnine_unit_897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11201)
);

ninexnine_unit ninexnine_unit_898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12201)
);

ninexnine_unit ninexnine_unit_899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13201)
);

assign C1201=c10201+c11201+c12201+c13201;
assign A1201=(C1201>=0)?1:0;

ninexnine_unit ninexnine_unit_900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10211)
);

ninexnine_unit ninexnine_unit_901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11211)
);

ninexnine_unit ninexnine_unit_902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12211)
);

ninexnine_unit ninexnine_unit_903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13211)
);

assign C1211=c10211+c11211+c12211+c13211;
assign A1211=(C1211>=0)?1:0;

ninexnine_unit ninexnine_unit_904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10221)
);

ninexnine_unit ninexnine_unit_905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11221)
);

ninexnine_unit ninexnine_unit_906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12221)
);

ninexnine_unit ninexnine_unit_907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13221)
);

assign C1221=c10221+c11221+c12221+c13221;
assign A1221=(C1221>=0)?1:0;

ninexnine_unit ninexnine_unit_908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10231)
);

ninexnine_unit ninexnine_unit_909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11231)
);

ninexnine_unit ninexnine_unit_910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12231)
);

ninexnine_unit ninexnine_unit_911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13231)
);

assign C1231=c10231+c11231+c12231+c13231;
assign A1231=(C1231>=0)?1:0;

ninexnine_unit ninexnine_unit_912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10241)
);

ninexnine_unit ninexnine_unit_913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11241)
);

ninexnine_unit ninexnine_unit_914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12241)
);

ninexnine_unit ninexnine_unit_915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13241)
);

assign C1241=c10241+c11241+c12241+c13241;
assign A1241=(C1241>=0)?1:0;

ninexnine_unit ninexnine_unit_916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10251)
);

ninexnine_unit ninexnine_unit_917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11251)
);

ninexnine_unit ninexnine_unit_918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12251)
);

ninexnine_unit ninexnine_unit_919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13251)
);

assign C1251=c10251+c11251+c12251+c13251;
assign A1251=(C1251>=0)?1:0;

ninexnine_unit ninexnine_unit_920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10261)
);

ninexnine_unit ninexnine_unit_921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11261)
);

ninexnine_unit ninexnine_unit_922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12261)
);

ninexnine_unit ninexnine_unit_923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13261)
);

assign C1261=c10261+c11261+c12261+c13261;
assign A1261=(C1261>=0)?1:0;

ninexnine_unit ninexnine_unit_924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10271)
);

ninexnine_unit ninexnine_unit_925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11271)
);

ninexnine_unit ninexnine_unit_926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12271)
);

ninexnine_unit ninexnine_unit_927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13271)
);

assign C1271=c10271+c11271+c12271+c13271;
assign A1271=(C1271>=0)?1:0;

ninexnine_unit ninexnine_unit_928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10281)
);

ninexnine_unit ninexnine_unit_929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11281)
);

ninexnine_unit ninexnine_unit_930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12281)
);

ninexnine_unit ninexnine_unit_931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13281)
);

assign C1281=c10281+c11281+c12281+c13281;
assign A1281=(C1281>=0)?1:0;

ninexnine_unit ninexnine_unit_932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10291)
);

ninexnine_unit ninexnine_unit_933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11291)
);

ninexnine_unit ninexnine_unit_934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12291)
);

ninexnine_unit ninexnine_unit_935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13291)
);

assign C1291=c10291+c11291+c12291+c13291;
assign A1291=(C1291>=0)?1:0;

ninexnine_unit ninexnine_unit_936(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c102A1)
);

ninexnine_unit ninexnine_unit_937(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c112A1)
);

ninexnine_unit ninexnine_unit_938(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c122A1)
);

ninexnine_unit ninexnine_unit_939(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c132A1)
);

assign C12A1=c102A1+c112A1+c122A1+c132A1;
assign A12A1=(C12A1>=0)?1:0;

ninexnine_unit ninexnine_unit_940(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c102B1)
);

ninexnine_unit ninexnine_unit_941(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c112B1)
);

ninexnine_unit ninexnine_unit_942(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c122B1)
);

ninexnine_unit ninexnine_unit_943(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c132B1)
);

assign C12B1=c102B1+c112B1+c122B1+c132B1;
assign A12B1=(C12B1>=0)?1:0;

ninexnine_unit ninexnine_unit_944(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c102C1)
);

ninexnine_unit ninexnine_unit_945(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c112C1)
);

ninexnine_unit ninexnine_unit_946(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c122C1)
);

ninexnine_unit ninexnine_unit_947(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c132C1)
);

assign C12C1=c102C1+c112C1+c122C1+c132C1;
assign A12C1=(C12C1>=0)?1:0;

ninexnine_unit ninexnine_unit_948(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c102D1)
);

ninexnine_unit ninexnine_unit_949(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c112D1)
);

ninexnine_unit ninexnine_unit_950(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c122D1)
);

ninexnine_unit ninexnine_unit_951(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c132D1)
);

assign C12D1=c102D1+c112D1+c122D1+c132D1;
assign A12D1=(C12D1>=0)?1:0;

ninexnine_unit ninexnine_unit_952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10301)
);

ninexnine_unit ninexnine_unit_953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11301)
);

ninexnine_unit ninexnine_unit_954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12301)
);

ninexnine_unit ninexnine_unit_955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13301)
);

assign C1301=c10301+c11301+c12301+c13301;
assign A1301=(C1301>=0)?1:0;

ninexnine_unit ninexnine_unit_956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10311)
);

ninexnine_unit ninexnine_unit_957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11311)
);

ninexnine_unit ninexnine_unit_958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12311)
);

ninexnine_unit ninexnine_unit_959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13311)
);

assign C1311=c10311+c11311+c12311+c13311;
assign A1311=(C1311>=0)?1:0;

ninexnine_unit ninexnine_unit_960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10321)
);

ninexnine_unit ninexnine_unit_961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11321)
);

ninexnine_unit ninexnine_unit_962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12321)
);

ninexnine_unit ninexnine_unit_963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13321)
);

assign C1321=c10321+c11321+c12321+c13321;
assign A1321=(C1321>=0)?1:0;

ninexnine_unit ninexnine_unit_964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10331)
);

ninexnine_unit ninexnine_unit_965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11331)
);

ninexnine_unit ninexnine_unit_966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12331)
);

ninexnine_unit ninexnine_unit_967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13331)
);

assign C1331=c10331+c11331+c12331+c13331;
assign A1331=(C1331>=0)?1:0;

ninexnine_unit ninexnine_unit_968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10341)
);

ninexnine_unit ninexnine_unit_969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11341)
);

ninexnine_unit ninexnine_unit_970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12341)
);

ninexnine_unit ninexnine_unit_971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13341)
);

assign C1341=c10341+c11341+c12341+c13341;
assign A1341=(C1341>=0)?1:0;

ninexnine_unit ninexnine_unit_972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10351)
);

ninexnine_unit ninexnine_unit_973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11351)
);

ninexnine_unit ninexnine_unit_974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12351)
);

ninexnine_unit ninexnine_unit_975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13351)
);

assign C1351=c10351+c11351+c12351+c13351;
assign A1351=(C1351>=0)?1:0;

ninexnine_unit ninexnine_unit_976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10361)
);

ninexnine_unit ninexnine_unit_977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11361)
);

ninexnine_unit ninexnine_unit_978(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12361)
);

ninexnine_unit ninexnine_unit_979(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13361)
);

assign C1361=c10361+c11361+c12361+c13361;
assign A1361=(C1361>=0)?1:0;

ninexnine_unit ninexnine_unit_980(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10371)
);

ninexnine_unit ninexnine_unit_981(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11371)
);

ninexnine_unit ninexnine_unit_982(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12371)
);

ninexnine_unit ninexnine_unit_983(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13371)
);

assign C1371=c10371+c11371+c12371+c13371;
assign A1371=(C1371>=0)?1:0;

ninexnine_unit ninexnine_unit_984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10381)
);

ninexnine_unit ninexnine_unit_985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11381)
);

ninexnine_unit ninexnine_unit_986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12381)
);

ninexnine_unit ninexnine_unit_987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13381)
);

assign C1381=c10381+c11381+c12381+c13381;
assign A1381=(C1381>=0)?1:0;

ninexnine_unit ninexnine_unit_988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10391)
);

ninexnine_unit ninexnine_unit_989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11391)
);

ninexnine_unit ninexnine_unit_990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12391)
);

ninexnine_unit ninexnine_unit_991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13391)
);

assign C1391=c10391+c11391+c12391+c13391;
assign A1391=(C1391>=0)?1:0;

ninexnine_unit ninexnine_unit_992(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c103A1)
);

ninexnine_unit ninexnine_unit_993(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c113A1)
);

ninexnine_unit ninexnine_unit_994(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c123A1)
);

ninexnine_unit ninexnine_unit_995(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c133A1)
);

assign C13A1=c103A1+c113A1+c123A1+c133A1;
assign A13A1=(C13A1>=0)?1:0;

ninexnine_unit ninexnine_unit_996(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c103B1)
);

ninexnine_unit ninexnine_unit_997(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c113B1)
);

ninexnine_unit ninexnine_unit_998(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c123B1)
);

ninexnine_unit ninexnine_unit_999(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c133B1)
);

assign C13B1=c103B1+c113B1+c123B1+c133B1;
assign A13B1=(C13B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1000(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c103C1)
);

ninexnine_unit ninexnine_unit_1001(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c113C1)
);

ninexnine_unit ninexnine_unit_1002(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c123C1)
);

ninexnine_unit ninexnine_unit_1003(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c133C1)
);

assign C13C1=c103C1+c113C1+c123C1+c133C1;
assign A13C1=(C13C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1004(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c103D1)
);

ninexnine_unit ninexnine_unit_1005(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c113D1)
);

ninexnine_unit ninexnine_unit_1006(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c123D1)
);

ninexnine_unit ninexnine_unit_1007(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c133D1)
);

assign C13D1=c103D1+c113D1+c123D1+c133D1;
assign A13D1=(C13D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10401)
);

ninexnine_unit ninexnine_unit_1009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11401)
);

ninexnine_unit ninexnine_unit_1010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12401)
);

ninexnine_unit ninexnine_unit_1011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13401)
);

assign C1401=c10401+c11401+c12401+c13401;
assign A1401=(C1401>=0)?1:0;

ninexnine_unit ninexnine_unit_1012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10411)
);

ninexnine_unit ninexnine_unit_1013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11411)
);

ninexnine_unit ninexnine_unit_1014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12411)
);

ninexnine_unit ninexnine_unit_1015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13411)
);

assign C1411=c10411+c11411+c12411+c13411;
assign A1411=(C1411>=0)?1:0;

ninexnine_unit ninexnine_unit_1016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10421)
);

ninexnine_unit ninexnine_unit_1017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11421)
);

ninexnine_unit ninexnine_unit_1018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12421)
);

ninexnine_unit ninexnine_unit_1019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13421)
);

assign C1421=c10421+c11421+c12421+c13421;
assign A1421=(C1421>=0)?1:0;

ninexnine_unit ninexnine_unit_1020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10431)
);

ninexnine_unit ninexnine_unit_1021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11431)
);

ninexnine_unit ninexnine_unit_1022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12431)
);

ninexnine_unit ninexnine_unit_1023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13431)
);

assign C1431=c10431+c11431+c12431+c13431;
assign A1431=(C1431>=0)?1:0;

ninexnine_unit ninexnine_unit_1024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10441)
);

ninexnine_unit ninexnine_unit_1025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11441)
);

ninexnine_unit ninexnine_unit_1026(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12441)
);

ninexnine_unit ninexnine_unit_1027(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13441)
);

assign C1441=c10441+c11441+c12441+c13441;
assign A1441=(C1441>=0)?1:0;

ninexnine_unit ninexnine_unit_1028(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10451)
);

ninexnine_unit ninexnine_unit_1029(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11451)
);

ninexnine_unit ninexnine_unit_1030(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12451)
);

ninexnine_unit ninexnine_unit_1031(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13451)
);

assign C1451=c10451+c11451+c12451+c13451;
assign A1451=(C1451>=0)?1:0;

ninexnine_unit ninexnine_unit_1032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10461)
);

ninexnine_unit ninexnine_unit_1033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11461)
);

ninexnine_unit ninexnine_unit_1034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12461)
);

ninexnine_unit ninexnine_unit_1035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13461)
);

assign C1461=c10461+c11461+c12461+c13461;
assign A1461=(C1461>=0)?1:0;

ninexnine_unit ninexnine_unit_1036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10471)
);

ninexnine_unit ninexnine_unit_1037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11471)
);

ninexnine_unit ninexnine_unit_1038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12471)
);

ninexnine_unit ninexnine_unit_1039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13471)
);

assign C1471=c10471+c11471+c12471+c13471;
assign A1471=(C1471>=0)?1:0;

ninexnine_unit ninexnine_unit_1040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10481)
);

ninexnine_unit ninexnine_unit_1041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11481)
);

ninexnine_unit ninexnine_unit_1042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12481)
);

ninexnine_unit ninexnine_unit_1043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13481)
);

assign C1481=c10481+c11481+c12481+c13481;
assign A1481=(C1481>=0)?1:0;

ninexnine_unit ninexnine_unit_1044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10491)
);

ninexnine_unit ninexnine_unit_1045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11491)
);

ninexnine_unit ninexnine_unit_1046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12491)
);

ninexnine_unit ninexnine_unit_1047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13491)
);

assign C1491=c10491+c11491+c12491+c13491;
assign A1491=(C1491>=0)?1:0;

ninexnine_unit ninexnine_unit_1048(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c104A1)
);

ninexnine_unit ninexnine_unit_1049(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c114A1)
);

ninexnine_unit ninexnine_unit_1050(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c124A1)
);

ninexnine_unit ninexnine_unit_1051(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c134A1)
);

assign C14A1=c104A1+c114A1+c124A1+c134A1;
assign A14A1=(C14A1>=0)?1:0;

ninexnine_unit ninexnine_unit_1052(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c104B1)
);

ninexnine_unit ninexnine_unit_1053(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c114B1)
);

ninexnine_unit ninexnine_unit_1054(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c124B1)
);

ninexnine_unit ninexnine_unit_1055(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c134B1)
);

assign C14B1=c104B1+c114B1+c124B1+c134B1;
assign A14B1=(C14B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1056(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c104C1)
);

ninexnine_unit ninexnine_unit_1057(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c114C1)
);

ninexnine_unit ninexnine_unit_1058(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c124C1)
);

ninexnine_unit ninexnine_unit_1059(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c134C1)
);

assign C14C1=c104C1+c114C1+c124C1+c134C1;
assign A14C1=(C14C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1060(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c104D1)
);

ninexnine_unit ninexnine_unit_1061(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c114D1)
);

ninexnine_unit ninexnine_unit_1062(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c124D1)
);

ninexnine_unit ninexnine_unit_1063(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c134D1)
);

assign C14D1=c104D1+c114D1+c124D1+c134D1;
assign A14D1=(C14D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10501)
);

ninexnine_unit ninexnine_unit_1065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11501)
);

ninexnine_unit ninexnine_unit_1066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12501)
);

ninexnine_unit ninexnine_unit_1067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13501)
);

assign C1501=c10501+c11501+c12501+c13501;
assign A1501=(C1501>=0)?1:0;

ninexnine_unit ninexnine_unit_1068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10511)
);

ninexnine_unit ninexnine_unit_1069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11511)
);

ninexnine_unit ninexnine_unit_1070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12511)
);

ninexnine_unit ninexnine_unit_1071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13511)
);

assign C1511=c10511+c11511+c12511+c13511;
assign A1511=(C1511>=0)?1:0;

ninexnine_unit ninexnine_unit_1072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10521)
);

ninexnine_unit ninexnine_unit_1073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11521)
);

ninexnine_unit ninexnine_unit_1074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12521)
);

ninexnine_unit ninexnine_unit_1075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13521)
);

assign C1521=c10521+c11521+c12521+c13521;
assign A1521=(C1521>=0)?1:0;

ninexnine_unit ninexnine_unit_1076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10531)
);

ninexnine_unit ninexnine_unit_1077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11531)
);

ninexnine_unit ninexnine_unit_1078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12531)
);

ninexnine_unit ninexnine_unit_1079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13531)
);

assign C1531=c10531+c11531+c12531+c13531;
assign A1531=(C1531>=0)?1:0;

ninexnine_unit ninexnine_unit_1080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10541)
);

ninexnine_unit ninexnine_unit_1081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11541)
);

ninexnine_unit ninexnine_unit_1082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12541)
);

ninexnine_unit ninexnine_unit_1083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13541)
);

assign C1541=c10541+c11541+c12541+c13541;
assign A1541=(C1541>=0)?1:0;

ninexnine_unit ninexnine_unit_1084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10551)
);

ninexnine_unit ninexnine_unit_1085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11551)
);

ninexnine_unit ninexnine_unit_1086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12551)
);

ninexnine_unit ninexnine_unit_1087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13551)
);

assign C1551=c10551+c11551+c12551+c13551;
assign A1551=(C1551>=0)?1:0;

ninexnine_unit ninexnine_unit_1088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10561)
);

ninexnine_unit ninexnine_unit_1089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11561)
);

ninexnine_unit ninexnine_unit_1090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12561)
);

ninexnine_unit ninexnine_unit_1091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13561)
);

assign C1561=c10561+c11561+c12561+c13561;
assign A1561=(C1561>=0)?1:0;

ninexnine_unit ninexnine_unit_1092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10571)
);

ninexnine_unit ninexnine_unit_1093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11571)
);

ninexnine_unit ninexnine_unit_1094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12571)
);

ninexnine_unit ninexnine_unit_1095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13571)
);

assign C1571=c10571+c11571+c12571+c13571;
assign A1571=(C1571>=0)?1:0;

ninexnine_unit ninexnine_unit_1096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10581)
);

ninexnine_unit ninexnine_unit_1097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11581)
);

ninexnine_unit ninexnine_unit_1098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12581)
);

ninexnine_unit ninexnine_unit_1099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13581)
);

assign C1581=c10581+c11581+c12581+c13581;
assign A1581=(C1581>=0)?1:0;

ninexnine_unit ninexnine_unit_1100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10591)
);

ninexnine_unit ninexnine_unit_1101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11591)
);

ninexnine_unit ninexnine_unit_1102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12591)
);

ninexnine_unit ninexnine_unit_1103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13591)
);

assign C1591=c10591+c11591+c12591+c13591;
assign A1591=(C1591>=0)?1:0;

ninexnine_unit ninexnine_unit_1104(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c105A1)
);

ninexnine_unit ninexnine_unit_1105(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c115A1)
);

ninexnine_unit ninexnine_unit_1106(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c125A1)
);

ninexnine_unit ninexnine_unit_1107(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c135A1)
);

assign C15A1=c105A1+c115A1+c125A1+c135A1;
assign A15A1=(C15A1>=0)?1:0;

ninexnine_unit ninexnine_unit_1108(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c105B1)
);

ninexnine_unit ninexnine_unit_1109(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c115B1)
);

ninexnine_unit ninexnine_unit_1110(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c125B1)
);

ninexnine_unit ninexnine_unit_1111(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c135B1)
);

assign C15B1=c105B1+c115B1+c125B1+c135B1;
assign A15B1=(C15B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1112(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c105C1)
);

ninexnine_unit ninexnine_unit_1113(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c115C1)
);

ninexnine_unit ninexnine_unit_1114(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c125C1)
);

ninexnine_unit ninexnine_unit_1115(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c135C1)
);

assign C15C1=c105C1+c115C1+c125C1+c135C1;
assign A15C1=(C15C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1116(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c105D1)
);

ninexnine_unit ninexnine_unit_1117(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c115D1)
);

ninexnine_unit ninexnine_unit_1118(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c125D1)
);

ninexnine_unit ninexnine_unit_1119(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c135D1)
);

assign C15D1=c105D1+c115D1+c125D1+c135D1;
assign A15D1=(C15D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10601)
);

ninexnine_unit ninexnine_unit_1121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11601)
);

ninexnine_unit ninexnine_unit_1122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12601)
);

ninexnine_unit ninexnine_unit_1123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13601)
);

assign C1601=c10601+c11601+c12601+c13601;
assign A1601=(C1601>=0)?1:0;

ninexnine_unit ninexnine_unit_1124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10611)
);

ninexnine_unit ninexnine_unit_1125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11611)
);

ninexnine_unit ninexnine_unit_1126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12611)
);

ninexnine_unit ninexnine_unit_1127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13611)
);

assign C1611=c10611+c11611+c12611+c13611;
assign A1611=(C1611>=0)?1:0;

ninexnine_unit ninexnine_unit_1128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10621)
);

ninexnine_unit ninexnine_unit_1129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11621)
);

ninexnine_unit ninexnine_unit_1130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12621)
);

ninexnine_unit ninexnine_unit_1131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13621)
);

assign C1621=c10621+c11621+c12621+c13621;
assign A1621=(C1621>=0)?1:0;

ninexnine_unit ninexnine_unit_1132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10631)
);

ninexnine_unit ninexnine_unit_1133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11631)
);

ninexnine_unit ninexnine_unit_1134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12631)
);

ninexnine_unit ninexnine_unit_1135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13631)
);

assign C1631=c10631+c11631+c12631+c13631;
assign A1631=(C1631>=0)?1:0;

ninexnine_unit ninexnine_unit_1136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10641)
);

ninexnine_unit ninexnine_unit_1137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11641)
);

ninexnine_unit ninexnine_unit_1138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12641)
);

ninexnine_unit ninexnine_unit_1139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13641)
);

assign C1641=c10641+c11641+c12641+c13641;
assign A1641=(C1641>=0)?1:0;

ninexnine_unit ninexnine_unit_1140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10651)
);

ninexnine_unit ninexnine_unit_1141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11651)
);

ninexnine_unit ninexnine_unit_1142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12651)
);

ninexnine_unit ninexnine_unit_1143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13651)
);

assign C1651=c10651+c11651+c12651+c13651;
assign A1651=(C1651>=0)?1:0;

ninexnine_unit ninexnine_unit_1144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10661)
);

ninexnine_unit ninexnine_unit_1145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11661)
);

ninexnine_unit ninexnine_unit_1146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12661)
);

ninexnine_unit ninexnine_unit_1147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13661)
);

assign C1661=c10661+c11661+c12661+c13661;
assign A1661=(C1661>=0)?1:0;

ninexnine_unit ninexnine_unit_1148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10671)
);

ninexnine_unit ninexnine_unit_1149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11671)
);

ninexnine_unit ninexnine_unit_1150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12671)
);

ninexnine_unit ninexnine_unit_1151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13671)
);

assign C1671=c10671+c11671+c12671+c13671;
assign A1671=(C1671>=0)?1:0;

ninexnine_unit ninexnine_unit_1152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10681)
);

ninexnine_unit ninexnine_unit_1153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11681)
);

ninexnine_unit ninexnine_unit_1154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12681)
);

ninexnine_unit ninexnine_unit_1155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13681)
);

assign C1681=c10681+c11681+c12681+c13681;
assign A1681=(C1681>=0)?1:0;

ninexnine_unit ninexnine_unit_1156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10691)
);

ninexnine_unit ninexnine_unit_1157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11691)
);

ninexnine_unit ninexnine_unit_1158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12691)
);

ninexnine_unit ninexnine_unit_1159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13691)
);

assign C1691=c10691+c11691+c12691+c13691;
assign A1691=(C1691>=0)?1:0;

ninexnine_unit ninexnine_unit_1160(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c106A1)
);

ninexnine_unit ninexnine_unit_1161(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c116A1)
);

ninexnine_unit ninexnine_unit_1162(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c126A1)
);

ninexnine_unit ninexnine_unit_1163(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c136A1)
);

assign C16A1=c106A1+c116A1+c126A1+c136A1;
assign A16A1=(C16A1>=0)?1:0;

ninexnine_unit ninexnine_unit_1164(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c106B1)
);

ninexnine_unit ninexnine_unit_1165(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c116B1)
);

ninexnine_unit ninexnine_unit_1166(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c126B1)
);

ninexnine_unit ninexnine_unit_1167(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c136B1)
);

assign C16B1=c106B1+c116B1+c126B1+c136B1;
assign A16B1=(C16B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1168(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c106C1)
);

ninexnine_unit ninexnine_unit_1169(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c116C1)
);

ninexnine_unit ninexnine_unit_1170(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c126C1)
);

ninexnine_unit ninexnine_unit_1171(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c136C1)
);

assign C16C1=c106C1+c116C1+c126C1+c136C1;
assign A16C1=(C16C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1172(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c106D1)
);

ninexnine_unit ninexnine_unit_1173(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c116D1)
);

ninexnine_unit ninexnine_unit_1174(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c126D1)
);

ninexnine_unit ninexnine_unit_1175(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c136D1)
);

assign C16D1=c106D1+c116D1+c126D1+c136D1;
assign A16D1=(C16D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10701)
);

ninexnine_unit ninexnine_unit_1177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11701)
);

ninexnine_unit ninexnine_unit_1178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12701)
);

ninexnine_unit ninexnine_unit_1179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13701)
);

assign C1701=c10701+c11701+c12701+c13701;
assign A1701=(C1701>=0)?1:0;

ninexnine_unit ninexnine_unit_1180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10711)
);

ninexnine_unit ninexnine_unit_1181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11711)
);

ninexnine_unit ninexnine_unit_1182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12711)
);

ninexnine_unit ninexnine_unit_1183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13711)
);

assign C1711=c10711+c11711+c12711+c13711;
assign A1711=(C1711>=0)?1:0;

ninexnine_unit ninexnine_unit_1184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10721)
);

ninexnine_unit ninexnine_unit_1185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11721)
);

ninexnine_unit ninexnine_unit_1186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12721)
);

ninexnine_unit ninexnine_unit_1187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13721)
);

assign C1721=c10721+c11721+c12721+c13721;
assign A1721=(C1721>=0)?1:0;

ninexnine_unit ninexnine_unit_1188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10731)
);

ninexnine_unit ninexnine_unit_1189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11731)
);

ninexnine_unit ninexnine_unit_1190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12731)
);

ninexnine_unit ninexnine_unit_1191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13731)
);

assign C1731=c10731+c11731+c12731+c13731;
assign A1731=(C1731>=0)?1:0;

ninexnine_unit ninexnine_unit_1192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10741)
);

ninexnine_unit ninexnine_unit_1193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11741)
);

ninexnine_unit ninexnine_unit_1194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12741)
);

ninexnine_unit ninexnine_unit_1195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13741)
);

assign C1741=c10741+c11741+c12741+c13741;
assign A1741=(C1741>=0)?1:0;

ninexnine_unit ninexnine_unit_1196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10751)
);

ninexnine_unit ninexnine_unit_1197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11751)
);

ninexnine_unit ninexnine_unit_1198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12751)
);

ninexnine_unit ninexnine_unit_1199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13751)
);

assign C1751=c10751+c11751+c12751+c13751;
assign A1751=(C1751>=0)?1:0;

ninexnine_unit ninexnine_unit_1200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10761)
);

ninexnine_unit ninexnine_unit_1201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11761)
);

ninexnine_unit ninexnine_unit_1202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12761)
);

ninexnine_unit ninexnine_unit_1203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13761)
);

assign C1761=c10761+c11761+c12761+c13761;
assign A1761=(C1761>=0)?1:0;

ninexnine_unit ninexnine_unit_1204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10771)
);

ninexnine_unit ninexnine_unit_1205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11771)
);

ninexnine_unit ninexnine_unit_1206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12771)
);

ninexnine_unit ninexnine_unit_1207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13771)
);

assign C1771=c10771+c11771+c12771+c13771;
assign A1771=(C1771>=0)?1:0;

ninexnine_unit ninexnine_unit_1208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10781)
);

ninexnine_unit ninexnine_unit_1209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11781)
);

ninexnine_unit ninexnine_unit_1210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12781)
);

ninexnine_unit ninexnine_unit_1211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13781)
);

assign C1781=c10781+c11781+c12781+c13781;
assign A1781=(C1781>=0)?1:0;

ninexnine_unit ninexnine_unit_1212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10791)
);

ninexnine_unit ninexnine_unit_1213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11791)
);

ninexnine_unit ninexnine_unit_1214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12791)
);

ninexnine_unit ninexnine_unit_1215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13791)
);

assign C1791=c10791+c11791+c12791+c13791;
assign A1791=(C1791>=0)?1:0;

ninexnine_unit ninexnine_unit_1216(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c107A1)
);

ninexnine_unit ninexnine_unit_1217(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c117A1)
);

ninexnine_unit ninexnine_unit_1218(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c127A1)
);

ninexnine_unit ninexnine_unit_1219(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c137A1)
);

assign C17A1=c107A1+c117A1+c127A1+c137A1;
assign A17A1=(C17A1>=0)?1:0;

ninexnine_unit ninexnine_unit_1220(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c107B1)
);

ninexnine_unit ninexnine_unit_1221(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c117B1)
);

ninexnine_unit ninexnine_unit_1222(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c127B1)
);

ninexnine_unit ninexnine_unit_1223(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c137B1)
);

assign C17B1=c107B1+c117B1+c127B1+c137B1;
assign A17B1=(C17B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1224(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c107C1)
);

ninexnine_unit ninexnine_unit_1225(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c117C1)
);

ninexnine_unit ninexnine_unit_1226(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c127C1)
);

ninexnine_unit ninexnine_unit_1227(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c137C1)
);

assign C17C1=c107C1+c117C1+c127C1+c137C1;
assign A17C1=(C17C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1228(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c107D1)
);

ninexnine_unit ninexnine_unit_1229(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c117D1)
);

ninexnine_unit ninexnine_unit_1230(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c127D1)
);

ninexnine_unit ninexnine_unit_1231(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c137D1)
);

assign C17D1=c107D1+c117D1+c127D1+c137D1;
assign A17D1=(C17D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10801)
);

ninexnine_unit ninexnine_unit_1233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11801)
);

ninexnine_unit ninexnine_unit_1234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12801)
);

ninexnine_unit ninexnine_unit_1235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13801)
);

assign C1801=c10801+c11801+c12801+c13801;
assign A1801=(C1801>=0)?1:0;

ninexnine_unit ninexnine_unit_1236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10811)
);

ninexnine_unit ninexnine_unit_1237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11811)
);

ninexnine_unit ninexnine_unit_1238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12811)
);

ninexnine_unit ninexnine_unit_1239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13811)
);

assign C1811=c10811+c11811+c12811+c13811;
assign A1811=(C1811>=0)?1:0;

ninexnine_unit ninexnine_unit_1240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10821)
);

ninexnine_unit ninexnine_unit_1241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11821)
);

ninexnine_unit ninexnine_unit_1242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12821)
);

ninexnine_unit ninexnine_unit_1243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13821)
);

assign C1821=c10821+c11821+c12821+c13821;
assign A1821=(C1821>=0)?1:0;

ninexnine_unit ninexnine_unit_1244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10831)
);

ninexnine_unit ninexnine_unit_1245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11831)
);

ninexnine_unit ninexnine_unit_1246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12831)
);

ninexnine_unit ninexnine_unit_1247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13831)
);

assign C1831=c10831+c11831+c12831+c13831;
assign A1831=(C1831>=0)?1:0;

ninexnine_unit ninexnine_unit_1248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10841)
);

ninexnine_unit ninexnine_unit_1249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11841)
);

ninexnine_unit ninexnine_unit_1250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12841)
);

ninexnine_unit ninexnine_unit_1251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13841)
);

assign C1841=c10841+c11841+c12841+c13841;
assign A1841=(C1841>=0)?1:0;

ninexnine_unit ninexnine_unit_1252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10851)
);

ninexnine_unit ninexnine_unit_1253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11851)
);

ninexnine_unit ninexnine_unit_1254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12851)
);

ninexnine_unit ninexnine_unit_1255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13851)
);

assign C1851=c10851+c11851+c12851+c13851;
assign A1851=(C1851>=0)?1:0;

ninexnine_unit ninexnine_unit_1256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10861)
);

ninexnine_unit ninexnine_unit_1257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11861)
);

ninexnine_unit ninexnine_unit_1258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12861)
);

ninexnine_unit ninexnine_unit_1259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13861)
);

assign C1861=c10861+c11861+c12861+c13861;
assign A1861=(C1861>=0)?1:0;

ninexnine_unit ninexnine_unit_1260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10871)
);

ninexnine_unit ninexnine_unit_1261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11871)
);

ninexnine_unit ninexnine_unit_1262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12871)
);

ninexnine_unit ninexnine_unit_1263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13871)
);

assign C1871=c10871+c11871+c12871+c13871;
assign A1871=(C1871>=0)?1:0;

ninexnine_unit ninexnine_unit_1264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10881)
);

ninexnine_unit ninexnine_unit_1265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11881)
);

ninexnine_unit ninexnine_unit_1266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12881)
);

ninexnine_unit ninexnine_unit_1267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13881)
);

assign C1881=c10881+c11881+c12881+c13881;
assign A1881=(C1881>=0)?1:0;

ninexnine_unit ninexnine_unit_1268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10891)
);

ninexnine_unit ninexnine_unit_1269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11891)
);

ninexnine_unit ninexnine_unit_1270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12891)
);

ninexnine_unit ninexnine_unit_1271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13891)
);

assign C1891=c10891+c11891+c12891+c13891;
assign A1891=(C1891>=0)?1:0;

ninexnine_unit ninexnine_unit_1272(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c108A1)
);

ninexnine_unit ninexnine_unit_1273(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c118A1)
);

ninexnine_unit ninexnine_unit_1274(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c128A1)
);

ninexnine_unit ninexnine_unit_1275(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c138A1)
);

assign C18A1=c108A1+c118A1+c128A1+c138A1;
assign A18A1=(C18A1>=0)?1:0;

ninexnine_unit ninexnine_unit_1276(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c108B1)
);

ninexnine_unit ninexnine_unit_1277(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c118B1)
);

ninexnine_unit ninexnine_unit_1278(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c128B1)
);

ninexnine_unit ninexnine_unit_1279(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c138B1)
);

assign C18B1=c108B1+c118B1+c128B1+c138B1;
assign A18B1=(C18B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1280(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c108C1)
);

ninexnine_unit ninexnine_unit_1281(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c118C1)
);

ninexnine_unit ninexnine_unit_1282(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c128C1)
);

ninexnine_unit ninexnine_unit_1283(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c138C1)
);

assign C18C1=c108C1+c118C1+c128C1+c138C1;
assign A18C1=(C18C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1284(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c108D1)
);

ninexnine_unit ninexnine_unit_1285(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c118D1)
);

ninexnine_unit ninexnine_unit_1286(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c128D1)
);

ninexnine_unit ninexnine_unit_1287(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c138D1)
);

assign C18D1=c108D1+c118D1+c128D1+c138D1;
assign A18D1=(C18D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10901)
);

ninexnine_unit ninexnine_unit_1289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11901)
);

ninexnine_unit ninexnine_unit_1290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12901)
);

ninexnine_unit ninexnine_unit_1291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13901)
);

assign C1901=c10901+c11901+c12901+c13901;
assign A1901=(C1901>=0)?1:0;

ninexnine_unit ninexnine_unit_1292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10911)
);

ninexnine_unit ninexnine_unit_1293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11911)
);

ninexnine_unit ninexnine_unit_1294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12911)
);

ninexnine_unit ninexnine_unit_1295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13911)
);

assign C1911=c10911+c11911+c12911+c13911;
assign A1911=(C1911>=0)?1:0;

ninexnine_unit ninexnine_unit_1296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10921)
);

ninexnine_unit ninexnine_unit_1297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11921)
);

ninexnine_unit ninexnine_unit_1298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12921)
);

ninexnine_unit ninexnine_unit_1299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13921)
);

assign C1921=c10921+c11921+c12921+c13921;
assign A1921=(C1921>=0)?1:0;

ninexnine_unit ninexnine_unit_1300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10931)
);

ninexnine_unit ninexnine_unit_1301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11931)
);

ninexnine_unit ninexnine_unit_1302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12931)
);

ninexnine_unit ninexnine_unit_1303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13931)
);

assign C1931=c10931+c11931+c12931+c13931;
assign A1931=(C1931>=0)?1:0;

ninexnine_unit ninexnine_unit_1304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10941)
);

ninexnine_unit ninexnine_unit_1305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11941)
);

ninexnine_unit ninexnine_unit_1306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12941)
);

ninexnine_unit ninexnine_unit_1307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13941)
);

assign C1941=c10941+c11941+c12941+c13941;
assign A1941=(C1941>=0)?1:0;

ninexnine_unit ninexnine_unit_1308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10951)
);

ninexnine_unit ninexnine_unit_1309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11951)
);

ninexnine_unit ninexnine_unit_1310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12951)
);

ninexnine_unit ninexnine_unit_1311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13951)
);

assign C1951=c10951+c11951+c12951+c13951;
assign A1951=(C1951>=0)?1:0;

ninexnine_unit ninexnine_unit_1312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10961)
);

ninexnine_unit ninexnine_unit_1313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11961)
);

ninexnine_unit ninexnine_unit_1314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12961)
);

ninexnine_unit ninexnine_unit_1315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13961)
);

assign C1961=c10961+c11961+c12961+c13961;
assign A1961=(C1961>=0)?1:0;

ninexnine_unit ninexnine_unit_1316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10971)
);

ninexnine_unit ninexnine_unit_1317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11971)
);

ninexnine_unit ninexnine_unit_1318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12971)
);

ninexnine_unit ninexnine_unit_1319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13971)
);

assign C1971=c10971+c11971+c12971+c13971;
assign A1971=(C1971>=0)?1:0;

ninexnine_unit ninexnine_unit_1320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10981)
);

ninexnine_unit ninexnine_unit_1321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11981)
);

ninexnine_unit ninexnine_unit_1322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12981)
);

ninexnine_unit ninexnine_unit_1323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13981)
);

assign C1981=c10981+c11981+c12981+c13981;
assign A1981=(C1981>=0)?1:0;

ninexnine_unit ninexnine_unit_1324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10991)
);

ninexnine_unit ninexnine_unit_1325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11991)
);

ninexnine_unit ninexnine_unit_1326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12991)
);

ninexnine_unit ninexnine_unit_1327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13991)
);

assign C1991=c10991+c11991+c12991+c13991;
assign A1991=(C1991>=0)?1:0;

ninexnine_unit ninexnine_unit_1328(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c109A1)
);

ninexnine_unit ninexnine_unit_1329(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c119A1)
);

ninexnine_unit ninexnine_unit_1330(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c129A1)
);

ninexnine_unit ninexnine_unit_1331(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c139A1)
);

assign C19A1=c109A1+c119A1+c129A1+c139A1;
assign A19A1=(C19A1>=0)?1:0;

ninexnine_unit ninexnine_unit_1332(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c109B1)
);

ninexnine_unit ninexnine_unit_1333(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c119B1)
);

ninexnine_unit ninexnine_unit_1334(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c129B1)
);

ninexnine_unit ninexnine_unit_1335(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c139B1)
);

assign C19B1=c109B1+c119B1+c129B1+c139B1;
assign A19B1=(C19B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1336(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c109C1)
);

ninexnine_unit ninexnine_unit_1337(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c119C1)
);

ninexnine_unit ninexnine_unit_1338(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c129C1)
);

ninexnine_unit ninexnine_unit_1339(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c139C1)
);

assign C19C1=c109C1+c119C1+c129C1+c139C1;
assign A19C1=(C19C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1340(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c109D1)
);

ninexnine_unit ninexnine_unit_1341(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c119D1)
);

ninexnine_unit ninexnine_unit_1342(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c129D1)
);

ninexnine_unit ninexnine_unit_1343(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c139D1)
);

assign C19D1=c109D1+c119D1+c129D1+c139D1;
assign A19D1=(C19D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A01)
);

ninexnine_unit ninexnine_unit_1345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A01)
);

ninexnine_unit ninexnine_unit_1346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A01)
);

ninexnine_unit ninexnine_unit_1347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A01)
);

assign C1A01=c10A01+c11A01+c12A01+c13A01;
assign A1A01=(C1A01>=0)?1:0;

ninexnine_unit ninexnine_unit_1348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A11)
);

ninexnine_unit ninexnine_unit_1349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A11)
);

ninexnine_unit ninexnine_unit_1350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A11)
);

ninexnine_unit ninexnine_unit_1351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A11)
);

assign C1A11=c10A11+c11A11+c12A11+c13A11;
assign A1A11=(C1A11>=0)?1:0;

ninexnine_unit ninexnine_unit_1352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A21)
);

ninexnine_unit ninexnine_unit_1353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A21)
);

ninexnine_unit ninexnine_unit_1354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A21)
);

ninexnine_unit ninexnine_unit_1355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A21)
);

assign C1A21=c10A21+c11A21+c12A21+c13A21;
assign A1A21=(C1A21>=0)?1:0;

ninexnine_unit ninexnine_unit_1356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A31)
);

ninexnine_unit ninexnine_unit_1357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A31)
);

ninexnine_unit ninexnine_unit_1358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A31)
);

ninexnine_unit ninexnine_unit_1359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A31)
);

assign C1A31=c10A31+c11A31+c12A31+c13A31;
assign A1A31=(C1A31>=0)?1:0;

ninexnine_unit ninexnine_unit_1360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A41)
);

ninexnine_unit ninexnine_unit_1361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A41)
);

ninexnine_unit ninexnine_unit_1362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A41)
);

ninexnine_unit ninexnine_unit_1363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A41)
);

assign C1A41=c10A41+c11A41+c12A41+c13A41;
assign A1A41=(C1A41>=0)?1:0;

ninexnine_unit ninexnine_unit_1364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A51)
);

ninexnine_unit ninexnine_unit_1365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A51)
);

ninexnine_unit ninexnine_unit_1366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A51)
);

ninexnine_unit ninexnine_unit_1367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A51)
);

assign C1A51=c10A51+c11A51+c12A51+c13A51;
assign A1A51=(C1A51>=0)?1:0;

ninexnine_unit ninexnine_unit_1368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A61)
);

ninexnine_unit ninexnine_unit_1369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A61)
);

ninexnine_unit ninexnine_unit_1370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A61)
);

ninexnine_unit ninexnine_unit_1371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A61)
);

assign C1A61=c10A61+c11A61+c12A61+c13A61;
assign A1A61=(C1A61>=0)?1:0;

ninexnine_unit ninexnine_unit_1372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A71)
);

ninexnine_unit ninexnine_unit_1373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A71)
);

ninexnine_unit ninexnine_unit_1374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A71)
);

ninexnine_unit ninexnine_unit_1375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A71)
);

assign C1A71=c10A71+c11A71+c12A71+c13A71;
assign A1A71=(C1A71>=0)?1:0;

ninexnine_unit ninexnine_unit_1376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A81)
);

ninexnine_unit ninexnine_unit_1377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A81)
);

ninexnine_unit ninexnine_unit_1378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A81)
);

ninexnine_unit ninexnine_unit_1379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A81)
);

assign C1A81=c10A81+c11A81+c12A81+c13A81;
assign A1A81=(C1A81>=0)?1:0;

ninexnine_unit ninexnine_unit_1380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10A91)
);

ninexnine_unit ninexnine_unit_1381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11A91)
);

ninexnine_unit ninexnine_unit_1382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12A91)
);

ninexnine_unit ninexnine_unit_1383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13A91)
);

assign C1A91=c10A91+c11A91+c12A91+c13A91;
assign A1A91=(C1A91>=0)?1:0;

ninexnine_unit ninexnine_unit_1384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10AA1)
);

ninexnine_unit ninexnine_unit_1385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11AA1)
);

ninexnine_unit ninexnine_unit_1386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12AA1)
);

ninexnine_unit ninexnine_unit_1387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13AA1)
);

assign C1AA1=c10AA1+c11AA1+c12AA1+c13AA1;
assign A1AA1=(C1AA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10AB1)
);

ninexnine_unit ninexnine_unit_1389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11AB1)
);

ninexnine_unit ninexnine_unit_1390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12AB1)
);

ninexnine_unit ninexnine_unit_1391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13AB1)
);

assign C1AB1=c10AB1+c11AB1+c12AB1+c13AB1;
assign A1AB1=(C1AB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10AC1)
);

ninexnine_unit ninexnine_unit_1393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11AC1)
);

ninexnine_unit ninexnine_unit_1394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12AC1)
);

ninexnine_unit ninexnine_unit_1395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13AC1)
);

assign C1AC1=c10AC1+c11AC1+c12AC1+c13AC1;
assign A1AC1=(C1AC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10AD1)
);

ninexnine_unit ninexnine_unit_1397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11AD1)
);

ninexnine_unit ninexnine_unit_1398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12AD1)
);

ninexnine_unit ninexnine_unit_1399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13AD1)
);

assign C1AD1=c10AD1+c11AD1+c12AD1+c13AD1;
assign A1AD1=(C1AD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B01)
);

ninexnine_unit ninexnine_unit_1401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B01)
);

ninexnine_unit ninexnine_unit_1402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B01)
);

ninexnine_unit ninexnine_unit_1403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B01)
);

assign C1B01=c10B01+c11B01+c12B01+c13B01;
assign A1B01=(C1B01>=0)?1:0;

ninexnine_unit ninexnine_unit_1404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B11)
);

ninexnine_unit ninexnine_unit_1405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B11)
);

ninexnine_unit ninexnine_unit_1406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B11)
);

ninexnine_unit ninexnine_unit_1407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B11)
);

assign C1B11=c10B11+c11B11+c12B11+c13B11;
assign A1B11=(C1B11>=0)?1:0;

ninexnine_unit ninexnine_unit_1408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B21)
);

ninexnine_unit ninexnine_unit_1409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B21)
);

ninexnine_unit ninexnine_unit_1410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B21)
);

ninexnine_unit ninexnine_unit_1411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B21)
);

assign C1B21=c10B21+c11B21+c12B21+c13B21;
assign A1B21=(C1B21>=0)?1:0;

ninexnine_unit ninexnine_unit_1412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B31)
);

ninexnine_unit ninexnine_unit_1413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B31)
);

ninexnine_unit ninexnine_unit_1414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B31)
);

ninexnine_unit ninexnine_unit_1415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B31)
);

assign C1B31=c10B31+c11B31+c12B31+c13B31;
assign A1B31=(C1B31>=0)?1:0;

ninexnine_unit ninexnine_unit_1416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B41)
);

ninexnine_unit ninexnine_unit_1417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B41)
);

ninexnine_unit ninexnine_unit_1418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B41)
);

ninexnine_unit ninexnine_unit_1419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B41)
);

assign C1B41=c10B41+c11B41+c12B41+c13B41;
assign A1B41=(C1B41>=0)?1:0;

ninexnine_unit ninexnine_unit_1420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B51)
);

ninexnine_unit ninexnine_unit_1421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B51)
);

ninexnine_unit ninexnine_unit_1422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B51)
);

ninexnine_unit ninexnine_unit_1423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B51)
);

assign C1B51=c10B51+c11B51+c12B51+c13B51;
assign A1B51=(C1B51>=0)?1:0;

ninexnine_unit ninexnine_unit_1424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B61)
);

ninexnine_unit ninexnine_unit_1425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B61)
);

ninexnine_unit ninexnine_unit_1426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B61)
);

ninexnine_unit ninexnine_unit_1427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B61)
);

assign C1B61=c10B61+c11B61+c12B61+c13B61;
assign A1B61=(C1B61>=0)?1:0;

ninexnine_unit ninexnine_unit_1428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B71)
);

ninexnine_unit ninexnine_unit_1429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B71)
);

ninexnine_unit ninexnine_unit_1430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B71)
);

ninexnine_unit ninexnine_unit_1431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B71)
);

assign C1B71=c10B71+c11B71+c12B71+c13B71;
assign A1B71=(C1B71>=0)?1:0;

ninexnine_unit ninexnine_unit_1432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B81)
);

ninexnine_unit ninexnine_unit_1433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B81)
);

ninexnine_unit ninexnine_unit_1434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B81)
);

ninexnine_unit ninexnine_unit_1435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B81)
);

assign C1B81=c10B81+c11B81+c12B81+c13B81;
assign A1B81=(C1B81>=0)?1:0;

ninexnine_unit ninexnine_unit_1436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10B91)
);

ninexnine_unit ninexnine_unit_1437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11B91)
);

ninexnine_unit ninexnine_unit_1438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12B91)
);

ninexnine_unit ninexnine_unit_1439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13B91)
);

assign C1B91=c10B91+c11B91+c12B91+c13B91;
assign A1B91=(C1B91>=0)?1:0;

ninexnine_unit ninexnine_unit_1440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10BA1)
);

ninexnine_unit ninexnine_unit_1441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11BA1)
);

ninexnine_unit ninexnine_unit_1442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12BA1)
);

ninexnine_unit ninexnine_unit_1443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13BA1)
);

assign C1BA1=c10BA1+c11BA1+c12BA1+c13BA1;
assign A1BA1=(C1BA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10BB1)
);

ninexnine_unit ninexnine_unit_1445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11BB1)
);

ninexnine_unit ninexnine_unit_1446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12BB1)
);

ninexnine_unit ninexnine_unit_1447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13BB1)
);

assign C1BB1=c10BB1+c11BB1+c12BB1+c13BB1;
assign A1BB1=(C1BB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10BC1)
);

ninexnine_unit ninexnine_unit_1449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11BC1)
);

ninexnine_unit ninexnine_unit_1450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12BC1)
);

ninexnine_unit ninexnine_unit_1451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13BC1)
);

assign C1BC1=c10BC1+c11BC1+c12BC1+c13BC1;
assign A1BC1=(C1BC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10BD1)
);

ninexnine_unit ninexnine_unit_1453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11BD1)
);

ninexnine_unit ninexnine_unit_1454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12BD1)
);

ninexnine_unit ninexnine_unit_1455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13BD1)
);

assign C1BD1=c10BD1+c11BD1+c12BD1+c13BD1;
assign A1BD1=(C1BD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C01)
);

ninexnine_unit ninexnine_unit_1457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C01)
);

ninexnine_unit ninexnine_unit_1458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C01)
);

ninexnine_unit ninexnine_unit_1459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C01)
);

assign C1C01=c10C01+c11C01+c12C01+c13C01;
assign A1C01=(C1C01>=0)?1:0;

ninexnine_unit ninexnine_unit_1460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C11)
);

ninexnine_unit ninexnine_unit_1461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C11)
);

ninexnine_unit ninexnine_unit_1462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C11)
);

ninexnine_unit ninexnine_unit_1463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C11)
);

assign C1C11=c10C11+c11C11+c12C11+c13C11;
assign A1C11=(C1C11>=0)?1:0;

ninexnine_unit ninexnine_unit_1464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C21)
);

ninexnine_unit ninexnine_unit_1465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C21)
);

ninexnine_unit ninexnine_unit_1466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C21)
);

ninexnine_unit ninexnine_unit_1467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C21)
);

assign C1C21=c10C21+c11C21+c12C21+c13C21;
assign A1C21=(C1C21>=0)?1:0;

ninexnine_unit ninexnine_unit_1468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C31)
);

ninexnine_unit ninexnine_unit_1469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C31)
);

ninexnine_unit ninexnine_unit_1470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C31)
);

ninexnine_unit ninexnine_unit_1471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C31)
);

assign C1C31=c10C31+c11C31+c12C31+c13C31;
assign A1C31=(C1C31>=0)?1:0;

ninexnine_unit ninexnine_unit_1472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C41)
);

ninexnine_unit ninexnine_unit_1473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C41)
);

ninexnine_unit ninexnine_unit_1474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C41)
);

ninexnine_unit ninexnine_unit_1475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C41)
);

assign C1C41=c10C41+c11C41+c12C41+c13C41;
assign A1C41=(C1C41>=0)?1:0;

ninexnine_unit ninexnine_unit_1476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C51)
);

ninexnine_unit ninexnine_unit_1477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C51)
);

ninexnine_unit ninexnine_unit_1478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C51)
);

ninexnine_unit ninexnine_unit_1479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C51)
);

assign C1C51=c10C51+c11C51+c12C51+c13C51;
assign A1C51=(C1C51>=0)?1:0;

ninexnine_unit ninexnine_unit_1480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C61)
);

ninexnine_unit ninexnine_unit_1481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C61)
);

ninexnine_unit ninexnine_unit_1482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C61)
);

ninexnine_unit ninexnine_unit_1483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C61)
);

assign C1C61=c10C61+c11C61+c12C61+c13C61;
assign A1C61=(C1C61>=0)?1:0;

ninexnine_unit ninexnine_unit_1484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C71)
);

ninexnine_unit ninexnine_unit_1485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C71)
);

ninexnine_unit ninexnine_unit_1486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C71)
);

ninexnine_unit ninexnine_unit_1487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C71)
);

assign C1C71=c10C71+c11C71+c12C71+c13C71;
assign A1C71=(C1C71>=0)?1:0;

ninexnine_unit ninexnine_unit_1488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C81)
);

ninexnine_unit ninexnine_unit_1489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C81)
);

ninexnine_unit ninexnine_unit_1490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C81)
);

ninexnine_unit ninexnine_unit_1491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C81)
);

assign C1C81=c10C81+c11C81+c12C81+c13C81;
assign A1C81=(C1C81>=0)?1:0;

ninexnine_unit ninexnine_unit_1492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10C91)
);

ninexnine_unit ninexnine_unit_1493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11C91)
);

ninexnine_unit ninexnine_unit_1494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12C91)
);

ninexnine_unit ninexnine_unit_1495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13C91)
);

assign C1C91=c10C91+c11C91+c12C91+c13C91;
assign A1C91=(C1C91>=0)?1:0;

ninexnine_unit ninexnine_unit_1496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10CA1)
);

ninexnine_unit ninexnine_unit_1497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11CA1)
);

ninexnine_unit ninexnine_unit_1498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12CA1)
);

ninexnine_unit ninexnine_unit_1499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13CA1)
);

assign C1CA1=c10CA1+c11CA1+c12CA1+c13CA1;
assign A1CA1=(C1CA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10CB1)
);

ninexnine_unit ninexnine_unit_1501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11CB1)
);

ninexnine_unit ninexnine_unit_1502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12CB1)
);

ninexnine_unit ninexnine_unit_1503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13CB1)
);

assign C1CB1=c10CB1+c11CB1+c12CB1+c13CB1;
assign A1CB1=(C1CB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10CC1)
);

ninexnine_unit ninexnine_unit_1505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11CC1)
);

ninexnine_unit ninexnine_unit_1506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12CC1)
);

ninexnine_unit ninexnine_unit_1507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13CC1)
);

assign C1CC1=c10CC1+c11CC1+c12CC1+c13CC1;
assign A1CC1=(C1CC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10CD1)
);

ninexnine_unit ninexnine_unit_1509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11CD1)
);

ninexnine_unit ninexnine_unit_1510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12CD1)
);

ninexnine_unit ninexnine_unit_1511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13CD1)
);

assign C1CD1=c10CD1+c11CD1+c12CD1+c13CD1;
assign A1CD1=(C1CD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D01)
);

ninexnine_unit ninexnine_unit_1513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D01)
);

ninexnine_unit ninexnine_unit_1514(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D01)
);

ninexnine_unit ninexnine_unit_1515(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D01)
);

assign C1D01=c10D01+c11D01+c12D01+c13D01;
assign A1D01=(C1D01>=0)?1:0;

ninexnine_unit ninexnine_unit_1516(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D11)
);

ninexnine_unit ninexnine_unit_1517(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D11)
);

ninexnine_unit ninexnine_unit_1518(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D11)
);

ninexnine_unit ninexnine_unit_1519(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D11)
);

assign C1D11=c10D11+c11D11+c12D11+c13D11;
assign A1D11=(C1D11>=0)?1:0;

ninexnine_unit ninexnine_unit_1520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D21)
);

ninexnine_unit ninexnine_unit_1521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D21)
);

ninexnine_unit ninexnine_unit_1522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D21)
);

ninexnine_unit ninexnine_unit_1523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D21)
);

assign C1D21=c10D21+c11D21+c12D21+c13D21;
assign A1D21=(C1D21>=0)?1:0;

ninexnine_unit ninexnine_unit_1524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D31)
);

ninexnine_unit ninexnine_unit_1525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D31)
);

ninexnine_unit ninexnine_unit_1526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D31)
);

ninexnine_unit ninexnine_unit_1527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D31)
);

assign C1D31=c10D31+c11D31+c12D31+c13D31;
assign A1D31=(C1D31>=0)?1:0;

ninexnine_unit ninexnine_unit_1528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D41)
);

ninexnine_unit ninexnine_unit_1529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D41)
);

ninexnine_unit ninexnine_unit_1530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D41)
);

ninexnine_unit ninexnine_unit_1531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D41)
);

assign C1D41=c10D41+c11D41+c12D41+c13D41;
assign A1D41=(C1D41>=0)?1:0;

ninexnine_unit ninexnine_unit_1532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D51)
);

ninexnine_unit ninexnine_unit_1533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D51)
);

ninexnine_unit ninexnine_unit_1534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D51)
);

ninexnine_unit ninexnine_unit_1535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D51)
);

assign C1D51=c10D51+c11D51+c12D51+c13D51;
assign A1D51=(C1D51>=0)?1:0;

ninexnine_unit ninexnine_unit_1536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D61)
);

ninexnine_unit ninexnine_unit_1537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D61)
);

ninexnine_unit ninexnine_unit_1538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D61)
);

ninexnine_unit ninexnine_unit_1539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D61)
);

assign C1D61=c10D61+c11D61+c12D61+c13D61;
assign A1D61=(C1D61>=0)?1:0;

ninexnine_unit ninexnine_unit_1540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D71)
);

ninexnine_unit ninexnine_unit_1541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D71)
);

ninexnine_unit ninexnine_unit_1542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D71)
);

ninexnine_unit ninexnine_unit_1543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D71)
);

assign C1D71=c10D71+c11D71+c12D71+c13D71;
assign A1D71=(C1D71>=0)?1:0;

ninexnine_unit ninexnine_unit_1544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D81)
);

ninexnine_unit ninexnine_unit_1545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D81)
);

ninexnine_unit ninexnine_unit_1546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D81)
);

ninexnine_unit ninexnine_unit_1547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D81)
);

assign C1D81=c10D81+c11D81+c12D81+c13D81;
assign A1D81=(C1D81>=0)?1:0;

ninexnine_unit ninexnine_unit_1548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10D91)
);

ninexnine_unit ninexnine_unit_1549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11D91)
);

ninexnine_unit ninexnine_unit_1550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12D91)
);

ninexnine_unit ninexnine_unit_1551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13D91)
);

assign C1D91=c10D91+c11D91+c12D91+c13D91;
assign A1D91=(C1D91>=0)?1:0;

ninexnine_unit ninexnine_unit_1552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10DA1)
);

ninexnine_unit ninexnine_unit_1553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11DA1)
);

ninexnine_unit ninexnine_unit_1554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12DA1)
);

ninexnine_unit ninexnine_unit_1555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13DA1)
);

assign C1DA1=c10DA1+c11DA1+c12DA1+c13DA1;
assign A1DA1=(C1DA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10DB1)
);

ninexnine_unit ninexnine_unit_1557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11DB1)
);

ninexnine_unit ninexnine_unit_1558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12DB1)
);

ninexnine_unit ninexnine_unit_1559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13DB1)
);

assign C1DB1=c10DB1+c11DB1+c12DB1+c13DB1;
assign A1DB1=(C1DB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10DC1)
);

ninexnine_unit ninexnine_unit_1561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11DC1)
);

ninexnine_unit ninexnine_unit_1562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12DC1)
);

ninexnine_unit ninexnine_unit_1563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13DC1)
);

assign C1DC1=c10DC1+c11DC1+c12DC1+c13DC1;
assign A1DC1=(C1DC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10DD1)
);

ninexnine_unit ninexnine_unit_1565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11DD1)
);

ninexnine_unit ninexnine_unit_1566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12DD1)
);

ninexnine_unit ninexnine_unit_1567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13DD1)
);

assign C1DD1=c10DD1+c11DD1+c12DD1+c13DD1;
assign A1DD1=(C1DD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10002)
);

ninexnine_unit ninexnine_unit_1569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11002)
);

ninexnine_unit ninexnine_unit_1570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12002)
);

ninexnine_unit ninexnine_unit_1571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13002)
);

assign C1002=c10002+c11002+c12002+c13002;
assign A1002=(C1002>=0)?1:0;

ninexnine_unit ninexnine_unit_1572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10012)
);

ninexnine_unit ninexnine_unit_1573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11012)
);

ninexnine_unit ninexnine_unit_1574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12012)
);

ninexnine_unit ninexnine_unit_1575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13012)
);

assign C1012=c10012+c11012+c12012+c13012;
assign A1012=(C1012>=0)?1:0;

ninexnine_unit ninexnine_unit_1576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10022)
);

ninexnine_unit ninexnine_unit_1577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11022)
);

ninexnine_unit ninexnine_unit_1578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12022)
);

ninexnine_unit ninexnine_unit_1579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13022)
);

assign C1022=c10022+c11022+c12022+c13022;
assign A1022=(C1022>=0)?1:0;

ninexnine_unit ninexnine_unit_1580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10032)
);

ninexnine_unit ninexnine_unit_1581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11032)
);

ninexnine_unit ninexnine_unit_1582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12032)
);

ninexnine_unit ninexnine_unit_1583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13032)
);

assign C1032=c10032+c11032+c12032+c13032;
assign A1032=(C1032>=0)?1:0;

ninexnine_unit ninexnine_unit_1584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10042)
);

ninexnine_unit ninexnine_unit_1585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11042)
);

ninexnine_unit ninexnine_unit_1586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12042)
);

ninexnine_unit ninexnine_unit_1587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13042)
);

assign C1042=c10042+c11042+c12042+c13042;
assign A1042=(C1042>=0)?1:0;

ninexnine_unit ninexnine_unit_1588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10052)
);

ninexnine_unit ninexnine_unit_1589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11052)
);

ninexnine_unit ninexnine_unit_1590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12052)
);

ninexnine_unit ninexnine_unit_1591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13052)
);

assign C1052=c10052+c11052+c12052+c13052;
assign A1052=(C1052>=0)?1:0;

ninexnine_unit ninexnine_unit_1592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10062)
);

ninexnine_unit ninexnine_unit_1593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11062)
);

ninexnine_unit ninexnine_unit_1594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12062)
);

ninexnine_unit ninexnine_unit_1595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13062)
);

assign C1062=c10062+c11062+c12062+c13062;
assign A1062=(C1062>=0)?1:0;

ninexnine_unit ninexnine_unit_1596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10072)
);

ninexnine_unit ninexnine_unit_1597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11072)
);

ninexnine_unit ninexnine_unit_1598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12072)
);

ninexnine_unit ninexnine_unit_1599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13072)
);

assign C1072=c10072+c11072+c12072+c13072;
assign A1072=(C1072>=0)?1:0;

ninexnine_unit ninexnine_unit_1600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10082)
);

ninexnine_unit ninexnine_unit_1601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11082)
);

ninexnine_unit ninexnine_unit_1602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12082)
);

ninexnine_unit ninexnine_unit_1603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13082)
);

assign C1082=c10082+c11082+c12082+c13082;
assign A1082=(C1082>=0)?1:0;

ninexnine_unit ninexnine_unit_1604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10092)
);

ninexnine_unit ninexnine_unit_1605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11092)
);

ninexnine_unit ninexnine_unit_1606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12092)
);

ninexnine_unit ninexnine_unit_1607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13092)
);

assign C1092=c10092+c11092+c12092+c13092;
assign A1092=(C1092>=0)?1:0;

ninexnine_unit ninexnine_unit_1608(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c100A2)
);

ninexnine_unit ninexnine_unit_1609(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c110A2)
);

ninexnine_unit ninexnine_unit_1610(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c120A2)
);

ninexnine_unit ninexnine_unit_1611(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c130A2)
);

assign C10A2=c100A2+c110A2+c120A2+c130A2;
assign A10A2=(C10A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1612(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c100B2)
);

ninexnine_unit ninexnine_unit_1613(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c110B2)
);

ninexnine_unit ninexnine_unit_1614(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c120B2)
);

ninexnine_unit ninexnine_unit_1615(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c130B2)
);

assign C10B2=c100B2+c110B2+c120B2+c130B2;
assign A10B2=(C10B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1616(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c100C2)
);

ninexnine_unit ninexnine_unit_1617(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c110C2)
);

ninexnine_unit ninexnine_unit_1618(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c120C2)
);

ninexnine_unit ninexnine_unit_1619(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c130C2)
);

assign C10C2=c100C2+c110C2+c120C2+c130C2;
assign A10C2=(C10C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1620(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c100D2)
);

ninexnine_unit ninexnine_unit_1621(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c110D2)
);

ninexnine_unit ninexnine_unit_1622(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c120D2)
);

ninexnine_unit ninexnine_unit_1623(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c130D2)
);

assign C10D2=c100D2+c110D2+c120D2+c130D2;
assign A10D2=(C10D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10102)
);

ninexnine_unit ninexnine_unit_1625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11102)
);

ninexnine_unit ninexnine_unit_1626(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12102)
);

ninexnine_unit ninexnine_unit_1627(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13102)
);

assign C1102=c10102+c11102+c12102+c13102;
assign A1102=(C1102>=0)?1:0;

ninexnine_unit ninexnine_unit_1628(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10112)
);

ninexnine_unit ninexnine_unit_1629(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11112)
);

ninexnine_unit ninexnine_unit_1630(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12112)
);

ninexnine_unit ninexnine_unit_1631(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13112)
);

assign C1112=c10112+c11112+c12112+c13112;
assign A1112=(C1112>=0)?1:0;

ninexnine_unit ninexnine_unit_1632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10122)
);

ninexnine_unit ninexnine_unit_1633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11122)
);

ninexnine_unit ninexnine_unit_1634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12122)
);

ninexnine_unit ninexnine_unit_1635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13122)
);

assign C1122=c10122+c11122+c12122+c13122;
assign A1122=(C1122>=0)?1:0;

ninexnine_unit ninexnine_unit_1636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10132)
);

ninexnine_unit ninexnine_unit_1637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11132)
);

ninexnine_unit ninexnine_unit_1638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12132)
);

ninexnine_unit ninexnine_unit_1639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13132)
);

assign C1132=c10132+c11132+c12132+c13132;
assign A1132=(C1132>=0)?1:0;

ninexnine_unit ninexnine_unit_1640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10142)
);

ninexnine_unit ninexnine_unit_1641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11142)
);

ninexnine_unit ninexnine_unit_1642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12142)
);

ninexnine_unit ninexnine_unit_1643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13142)
);

assign C1142=c10142+c11142+c12142+c13142;
assign A1142=(C1142>=0)?1:0;

ninexnine_unit ninexnine_unit_1644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10152)
);

ninexnine_unit ninexnine_unit_1645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11152)
);

ninexnine_unit ninexnine_unit_1646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12152)
);

ninexnine_unit ninexnine_unit_1647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13152)
);

assign C1152=c10152+c11152+c12152+c13152;
assign A1152=(C1152>=0)?1:0;

ninexnine_unit ninexnine_unit_1648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10162)
);

ninexnine_unit ninexnine_unit_1649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11162)
);

ninexnine_unit ninexnine_unit_1650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12162)
);

ninexnine_unit ninexnine_unit_1651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13162)
);

assign C1162=c10162+c11162+c12162+c13162;
assign A1162=(C1162>=0)?1:0;

ninexnine_unit ninexnine_unit_1652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10172)
);

ninexnine_unit ninexnine_unit_1653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11172)
);

ninexnine_unit ninexnine_unit_1654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12172)
);

ninexnine_unit ninexnine_unit_1655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13172)
);

assign C1172=c10172+c11172+c12172+c13172;
assign A1172=(C1172>=0)?1:0;

ninexnine_unit ninexnine_unit_1656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10182)
);

ninexnine_unit ninexnine_unit_1657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11182)
);

ninexnine_unit ninexnine_unit_1658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12182)
);

ninexnine_unit ninexnine_unit_1659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13182)
);

assign C1182=c10182+c11182+c12182+c13182;
assign A1182=(C1182>=0)?1:0;

ninexnine_unit ninexnine_unit_1660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10192)
);

ninexnine_unit ninexnine_unit_1661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11192)
);

ninexnine_unit ninexnine_unit_1662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12192)
);

ninexnine_unit ninexnine_unit_1663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13192)
);

assign C1192=c10192+c11192+c12192+c13192;
assign A1192=(C1192>=0)?1:0;

ninexnine_unit ninexnine_unit_1664(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c101A2)
);

ninexnine_unit ninexnine_unit_1665(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c111A2)
);

ninexnine_unit ninexnine_unit_1666(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c121A2)
);

ninexnine_unit ninexnine_unit_1667(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c131A2)
);

assign C11A2=c101A2+c111A2+c121A2+c131A2;
assign A11A2=(C11A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1668(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c101B2)
);

ninexnine_unit ninexnine_unit_1669(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c111B2)
);

ninexnine_unit ninexnine_unit_1670(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c121B2)
);

ninexnine_unit ninexnine_unit_1671(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c131B2)
);

assign C11B2=c101B2+c111B2+c121B2+c131B2;
assign A11B2=(C11B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1672(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c101C2)
);

ninexnine_unit ninexnine_unit_1673(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c111C2)
);

ninexnine_unit ninexnine_unit_1674(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c121C2)
);

ninexnine_unit ninexnine_unit_1675(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c131C2)
);

assign C11C2=c101C2+c111C2+c121C2+c131C2;
assign A11C2=(C11C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1676(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c101D2)
);

ninexnine_unit ninexnine_unit_1677(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c111D2)
);

ninexnine_unit ninexnine_unit_1678(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c121D2)
);

ninexnine_unit ninexnine_unit_1679(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c131D2)
);

assign C11D2=c101D2+c111D2+c121D2+c131D2;
assign A11D2=(C11D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10202)
);

ninexnine_unit ninexnine_unit_1681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11202)
);

ninexnine_unit ninexnine_unit_1682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12202)
);

ninexnine_unit ninexnine_unit_1683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13202)
);

assign C1202=c10202+c11202+c12202+c13202;
assign A1202=(C1202>=0)?1:0;

ninexnine_unit ninexnine_unit_1684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10212)
);

ninexnine_unit ninexnine_unit_1685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11212)
);

ninexnine_unit ninexnine_unit_1686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12212)
);

ninexnine_unit ninexnine_unit_1687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13212)
);

assign C1212=c10212+c11212+c12212+c13212;
assign A1212=(C1212>=0)?1:0;

ninexnine_unit ninexnine_unit_1688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10222)
);

ninexnine_unit ninexnine_unit_1689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11222)
);

ninexnine_unit ninexnine_unit_1690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12222)
);

ninexnine_unit ninexnine_unit_1691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13222)
);

assign C1222=c10222+c11222+c12222+c13222;
assign A1222=(C1222>=0)?1:0;

ninexnine_unit ninexnine_unit_1692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10232)
);

ninexnine_unit ninexnine_unit_1693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11232)
);

ninexnine_unit ninexnine_unit_1694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12232)
);

ninexnine_unit ninexnine_unit_1695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13232)
);

assign C1232=c10232+c11232+c12232+c13232;
assign A1232=(C1232>=0)?1:0;

ninexnine_unit ninexnine_unit_1696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10242)
);

ninexnine_unit ninexnine_unit_1697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11242)
);

ninexnine_unit ninexnine_unit_1698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12242)
);

ninexnine_unit ninexnine_unit_1699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13242)
);

assign C1242=c10242+c11242+c12242+c13242;
assign A1242=(C1242>=0)?1:0;

ninexnine_unit ninexnine_unit_1700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10252)
);

ninexnine_unit ninexnine_unit_1701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11252)
);

ninexnine_unit ninexnine_unit_1702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12252)
);

ninexnine_unit ninexnine_unit_1703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13252)
);

assign C1252=c10252+c11252+c12252+c13252;
assign A1252=(C1252>=0)?1:0;

ninexnine_unit ninexnine_unit_1704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10262)
);

ninexnine_unit ninexnine_unit_1705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11262)
);

ninexnine_unit ninexnine_unit_1706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12262)
);

ninexnine_unit ninexnine_unit_1707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13262)
);

assign C1262=c10262+c11262+c12262+c13262;
assign A1262=(C1262>=0)?1:0;

ninexnine_unit ninexnine_unit_1708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10272)
);

ninexnine_unit ninexnine_unit_1709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11272)
);

ninexnine_unit ninexnine_unit_1710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12272)
);

ninexnine_unit ninexnine_unit_1711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13272)
);

assign C1272=c10272+c11272+c12272+c13272;
assign A1272=(C1272>=0)?1:0;

ninexnine_unit ninexnine_unit_1712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10282)
);

ninexnine_unit ninexnine_unit_1713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11282)
);

ninexnine_unit ninexnine_unit_1714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12282)
);

ninexnine_unit ninexnine_unit_1715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13282)
);

assign C1282=c10282+c11282+c12282+c13282;
assign A1282=(C1282>=0)?1:0;

ninexnine_unit ninexnine_unit_1716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10292)
);

ninexnine_unit ninexnine_unit_1717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11292)
);

ninexnine_unit ninexnine_unit_1718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12292)
);

ninexnine_unit ninexnine_unit_1719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13292)
);

assign C1292=c10292+c11292+c12292+c13292;
assign A1292=(C1292>=0)?1:0;

ninexnine_unit ninexnine_unit_1720(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c102A2)
);

ninexnine_unit ninexnine_unit_1721(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c112A2)
);

ninexnine_unit ninexnine_unit_1722(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c122A2)
);

ninexnine_unit ninexnine_unit_1723(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c132A2)
);

assign C12A2=c102A2+c112A2+c122A2+c132A2;
assign A12A2=(C12A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1724(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c102B2)
);

ninexnine_unit ninexnine_unit_1725(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c112B2)
);

ninexnine_unit ninexnine_unit_1726(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c122B2)
);

ninexnine_unit ninexnine_unit_1727(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c132B2)
);

assign C12B2=c102B2+c112B2+c122B2+c132B2;
assign A12B2=(C12B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1728(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c102C2)
);

ninexnine_unit ninexnine_unit_1729(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c112C2)
);

ninexnine_unit ninexnine_unit_1730(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c122C2)
);

ninexnine_unit ninexnine_unit_1731(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c132C2)
);

assign C12C2=c102C2+c112C2+c122C2+c132C2;
assign A12C2=(C12C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1732(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c102D2)
);

ninexnine_unit ninexnine_unit_1733(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c112D2)
);

ninexnine_unit ninexnine_unit_1734(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c122D2)
);

ninexnine_unit ninexnine_unit_1735(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c132D2)
);

assign C12D2=c102D2+c112D2+c122D2+c132D2;
assign A12D2=(C12D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10302)
);

ninexnine_unit ninexnine_unit_1737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11302)
);

ninexnine_unit ninexnine_unit_1738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12302)
);

ninexnine_unit ninexnine_unit_1739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13302)
);

assign C1302=c10302+c11302+c12302+c13302;
assign A1302=(C1302>=0)?1:0;

ninexnine_unit ninexnine_unit_1740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10312)
);

ninexnine_unit ninexnine_unit_1741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11312)
);

ninexnine_unit ninexnine_unit_1742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12312)
);

ninexnine_unit ninexnine_unit_1743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13312)
);

assign C1312=c10312+c11312+c12312+c13312;
assign A1312=(C1312>=0)?1:0;

ninexnine_unit ninexnine_unit_1744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10322)
);

ninexnine_unit ninexnine_unit_1745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11322)
);

ninexnine_unit ninexnine_unit_1746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12322)
);

ninexnine_unit ninexnine_unit_1747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13322)
);

assign C1322=c10322+c11322+c12322+c13322;
assign A1322=(C1322>=0)?1:0;

ninexnine_unit ninexnine_unit_1748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10332)
);

ninexnine_unit ninexnine_unit_1749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11332)
);

ninexnine_unit ninexnine_unit_1750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12332)
);

ninexnine_unit ninexnine_unit_1751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13332)
);

assign C1332=c10332+c11332+c12332+c13332;
assign A1332=(C1332>=0)?1:0;

ninexnine_unit ninexnine_unit_1752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10342)
);

ninexnine_unit ninexnine_unit_1753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11342)
);

ninexnine_unit ninexnine_unit_1754(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12342)
);

ninexnine_unit ninexnine_unit_1755(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13342)
);

assign C1342=c10342+c11342+c12342+c13342;
assign A1342=(C1342>=0)?1:0;

ninexnine_unit ninexnine_unit_1756(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10352)
);

ninexnine_unit ninexnine_unit_1757(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11352)
);

ninexnine_unit ninexnine_unit_1758(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12352)
);

ninexnine_unit ninexnine_unit_1759(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13352)
);

assign C1352=c10352+c11352+c12352+c13352;
assign A1352=(C1352>=0)?1:0;

ninexnine_unit ninexnine_unit_1760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10362)
);

ninexnine_unit ninexnine_unit_1761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11362)
);

ninexnine_unit ninexnine_unit_1762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12362)
);

ninexnine_unit ninexnine_unit_1763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13362)
);

assign C1362=c10362+c11362+c12362+c13362;
assign A1362=(C1362>=0)?1:0;

ninexnine_unit ninexnine_unit_1764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10372)
);

ninexnine_unit ninexnine_unit_1765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11372)
);

ninexnine_unit ninexnine_unit_1766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12372)
);

ninexnine_unit ninexnine_unit_1767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13372)
);

assign C1372=c10372+c11372+c12372+c13372;
assign A1372=(C1372>=0)?1:0;

ninexnine_unit ninexnine_unit_1768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10382)
);

ninexnine_unit ninexnine_unit_1769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11382)
);

ninexnine_unit ninexnine_unit_1770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12382)
);

ninexnine_unit ninexnine_unit_1771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13382)
);

assign C1382=c10382+c11382+c12382+c13382;
assign A1382=(C1382>=0)?1:0;

ninexnine_unit ninexnine_unit_1772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10392)
);

ninexnine_unit ninexnine_unit_1773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11392)
);

ninexnine_unit ninexnine_unit_1774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12392)
);

ninexnine_unit ninexnine_unit_1775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13392)
);

assign C1392=c10392+c11392+c12392+c13392;
assign A1392=(C1392>=0)?1:0;

ninexnine_unit ninexnine_unit_1776(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c103A2)
);

ninexnine_unit ninexnine_unit_1777(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c113A2)
);

ninexnine_unit ninexnine_unit_1778(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c123A2)
);

ninexnine_unit ninexnine_unit_1779(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c133A2)
);

assign C13A2=c103A2+c113A2+c123A2+c133A2;
assign A13A2=(C13A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1780(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c103B2)
);

ninexnine_unit ninexnine_unit_1781(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c113B2)
);

ninexnine_unit ninexnine_unit_1782(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c123B2)
);

ninexnine_unit ninexnine_unit_1783(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c133B2)
);

assign C13B2=c103B2+c113B2+c123B2+c133B2;
assign A13B2=(C13B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1784(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c103C2)
);

ninexnine_unit ninexnine_unit_1785(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c113C2)
);

ninexnine_unit ninexnine_unit_1786(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c123C2)
);

ninexnine_unit ninexnine_unit_1787(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c133C2)
);

assign C13C2=c103C2+c113C2+c123C2+c133C2;
assign A13C2=(C13C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1788(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c103D2)
);

ninexnine_unit ninexnine_unit_1789(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c113D2)
);

ninexnine_unit ninexnine_unit_1790(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c123D2)
);

ninexnine_unit ninexnine_unit_1791(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c133D2)
);

assign C13D2=c103D2+c113D2+c123D2+c133D2;
assign A13D2=(C13D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10402)
);

ninexnine_unit ninexnine_unit_1793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11402)
);

ninexnine_unit ninexnine_unit_1794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12402)
);

ninexnine_unit ninexnine_unit_1795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13402)
);

assign C1402=c10402+c11402+c12402+c13402;
assign A1402=(C1402>=0)?1:0;

ninexnine_unit ninexnine_unit_1796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10412)
);

ninexnine_unit ninexnine_unit_1797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11412)
);

ninexnine_unit ninexnine_unit_1798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12412)
);

ninexnine_unit ninexnine_unit_1799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13412)
);

assign C1412=c10412+c11412+c12412+c13412;
assign A1412=(C1412>=0)?1:0;

ninexnine_unit ninexnine_unit_1800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10422)
);

ninexnine_unit ninexnine_unit_1801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11422)
);

ninexnine_unit ninexnine_unit_1802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12422)
);

ninexnine_unit ninexnine_unit_1803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13422)
);

assign C1422=c10422+c11422+c12422+c13422;
assign A1422=(C1422>=0)?1:0;

ninexnine_unit ninexnine_unit_1804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10432)
);

ninexnine_unit ninexnine_unit_1805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11432)
);

ninexnine_unit ninexnine_unit_1806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12432)
);

ninexnine_unit ninexnine_unit_1807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13432)
);

assign C1432=c10432+c11432+c12432+c13432;
assign A1432=(C1432>=0)?1:0;

ninexnine_unit ninexnine_unit_1808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10442)
);

ninexnine_unit ninexnine_unit_1809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11442)
);

ninexnine_unit ninexnine_unit_1810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12442)
);

ninexnine_unit ninexnine_unit_1811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13442)
);

assign C1442=c10442+c11442+c12442+c13442;
assign A1442=(C1442>=0)?1:0;

ninexnine_unit ninexnine_unit_1812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10452)
);

ninexnine_unit ninexnine_unit_1813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11452)
);

ninexnine_unit ninexnine_unit_1814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12452)
);

ninexnine_unit ninexnine_unit_1815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13452)
);

assign C1452=c10452+c11452+c12452+c13452;
assign A1452=(C1452>=0)?1:0;

ninexnine_unit ninexnine_unit_1816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10462)
);

ninexnine_unit ninexnine_unit_1817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11462)
);

ninexnine_unit ninexnine_unit_1818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12462)
);

ninexnine_unit ninexnine_unit_1819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13462)
);

assign C1462=c10462+c11462+c12462+c13462;
assign A1462=(C1462>=0)?1:0;

ninexnine_unit ninexnine_unit_1820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10472)
);

ninexnine_unit ninexnine_unit_1821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11472)
);

ninexnine_unit ninexnine_unit_1822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12472)
);

ninexnine_unit ninexnine_unit_1823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13472)
);

assign C1472=c10472+c11472+c12472+c13472;
assign A1472=(C1472>=0)?1:0;

ninexnine_unit ninexnine_unit_1824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10482)
);

ninexnine_unit ninexnine_unit_1825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11482)
);

ninexnine_unit ninexnine_unit_1826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12482)
);

ninexnine_unit ninexnine_unit_1827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13482)
);

assign C1482=c10482+c11482+c12482+c13482;
assign A1482=(C1482>=0)?1:0;

ninexnine_unit ninexnine_unit_1828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10492)
);

ninexnine_unit ninexnine_unit_1829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11492)
);

ninexnine_unit ninexnine_unit_1830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12492)
);

ninexnine_unit ninexnine_unit_1831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13492)
);

assign C1492=c10492+c11492+c12492+c13492;
assign A1492=(C1492>=0)?1:0;

ninexnine_unit ninexnine_unit_1832(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c104A2)
);

ninexnine_unit ninexnine_unit_1833(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c114A2)
);

ninexnine_unit ninexnine_unit_1834(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c124A2)
);

ninexnine_unit ninexnine_unit_1835(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c134A2)
);

assign C14A2=c104A2+c114A2+c124A2+c134A2;
assign A14A2=(C14A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1836(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c104B2)
);

ninexnine_unit ninexnine_unit_1837(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c114B2)
);

ninexnine_unit ninexnine_unit_1838(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c124B2)
);

ninexnine_unit ninexnine_unit_1839(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c134B2)
);

assign C14B2=c104B2+c114B2+c124B2+c134B2;
assign A14B2=(C14B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1840(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c104C2)
);

ninexnine_unit ninexnine_unit_1841(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c114C2)
);

ninexnine_unit ninexnine_unit_1842(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c124C2)
);

ninexnine_unit ninexnine_unit_1843(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c134C2)
);

assign C14C2=c104C2+c114C2+c124C2+c134C2;
assign A14C2=(C14C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1844(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c104D2)
);

ninexnine_unit ninexnine_unit_1845(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c114D2)
);

ninexnine_unit ninexnine_unit_1846(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c124D2)
);

ninexnine_unit ninexnine_unit_1847(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c134D2)
);

assign C14D2=c104D2+c114D2+c124D2+c134D2;
assign A14D2=(C14D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10502)
);

ninexnine_unit ninexnine_unit_1849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11502)
);

ninexnine_unit ninexnine_unit_1850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12502)
);

ninexnine_unit ninexnine_unit_1851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13502)
);

assign C1502=c10502+c11502+c12502+c13502;
assign A1502=(C1502>=0)?1:0;

ninexnine_unit ninexnine_unit_1852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10512)
);

ninexnine_unit ninexnine_unit_1853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11512)
);

ninexnine_unit ninexnine_unit_1854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12512)
);

ninexnine_unit ninexnine_unit_1855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13512)
);

assign C1512=c10512+c11512+c12512+c13512;
assign A1512=(C1512>=0)?1:0;

ninexnine_unit ninexnine_unit_1856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10522)
);

ninexnine_unit ninexnine_unit_1857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11522)
);

ninexnine_unit ninexnine_unit_1858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12522)
);

ninexnine_unit ninexnine_unit_1859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13522)
);

assign C1522=c10522+c11522+c12522+c13522;
assign A1522=(C1522>=0)?1:0;

ninexnine_unit ninexnine_unit_1860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10532)
);

ninexnine_unit ninexnine_unit_1861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11532)
);

ninexnine_unit ninexnine_unit_1862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12532)
);

ninexnine_unit ninexnine_unit_1863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13532)
);

assign C1532=c10532+c11532+c12532+c13532;
assign A1532=(C1532>=0)?1:0;

ninexnine_unit ninexnine_unit_1864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10542)
);

ninexnine_unit ninexnine_unit_1865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11542)
);

ninexnine_unit ninexnine_unit_1866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12542)
);

ninexnine_unit ninexnine_unit_1867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13542)
);

assign C1542=c10542+c11542+c12542+c13542;
assign A1542=(C1542>=0)?1:0;

ninexnine_unit ninexnine_unit_1868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10552)
);

ninexnine_unit ninexnine_unit_1869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11552)
);

ninexnine_unit ninexnine_unit_1870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12552)
);

ninexnine_unit ninexnine_unit_1871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13552)
);

assign C1552=c10552+c11552+c12552+c13552;
assign A1552=(C1552>=0)?1:0;

ninexnine_unit ninexnine_unit_1872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10562)
);

ninexnine_unit ninexnine_unit_1873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11562)
);

ninexnine_unit ninexnine_unit_1874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12562)
);

ninexnine_unit ninexnine_unit_1875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13562)
);

assign C1562=c10562+c11562+c12562+c13562;
assign A1562=(C1562>=0)?1:0;

ninexnine_unit ninexnine_unit_1876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10572)
);

ninexnine_unit ninexnine_unit_1877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11572)
);

ninexnine_unit ninexnine_unit_1878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12572)
);

ninexnine_unit ninexnine_unit_1879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13572)
);

assign C1572=c10572+c11572+c12572+c13572;
assign A1572=(C1572>=0)?1:0;

ninexnine_unit ninexnine_unit_1880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10582)
);

ninexnine_unit ninexnine_unit_1881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11582)
);

ninexnine_unit ninexnine_unit_1882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12582)
);

ninexnine_unit ninexnine_unit_1883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13582)
);

assign C1582=c10582+c11582+c12582+c13582;
assign A1582=(C1582>=0)?1:0;

ninexnine_unit ninexnine_unit_1884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10592)
);

ninexnine_unit ninexnine_unit_1885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11592)
);

ninexnine_unit ninexnine_unit_1886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12592)
);

ninexnine_unit ninexnine_unit_1887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13592)
);

assign C1592=c10592+c11592+c12592+c13592;
assign A1592=(C1592>=0)?1:0;

ninexnine_unit ninexnine_unit_1888(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c105A2)
);

ninexnine_unit ninexnine_unit_1889(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c115A2)
);

ninexnine_unit ninexnine_unit_1890(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c125A2)
);

ninexnine_unit ninexnine_unit_1891(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c135A2)
);

assign C15A2=c105A2+c115A2+c125A2+c135A2;
assign A15A2=(C15A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1892(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c105B2)
);

ninexnine_unit ninexnine_unit_1893(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c115B2)
);

ninexnine_unit ninexnine_unit_1894(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c125B2)
);

ninexnine_unit ninexnine_unit_1895(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c135B2)
);

assign C15B2=c105B2+c115B2+c125B2+c135B2;
assign A15B2=(C15B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1896(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c105C2)
);

ninexnine_unit ninexnine_unit_1897(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c115C2)
);

ninexnine_unit ninexnine_unit_1898(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c125C2)
);

ninexnine_unit ninexnine_unit_1899(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c135C2)
);

assign C15C2=c105C2+c115C2+c125C2+c135C2;
assign A15C2=(C15C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1900(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c105D2)
);

ninexnine_unit ninexnine_unit_1901(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c115D2)
);

ninexnine_unit ninexnine_unit_1902(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c125D2)
);

ninexnine_unit ninexnine_unit_1903(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c135D2)
);

assign C15D2=c105D2+c115D2+c125D2+c135D2;
assign A15D2=(C15D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10602)
);

ninexnine_unit ninexnine_unit_1905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11602)
);

ninexnine_unit ninexnine_unit_1906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12602)
);

ninexnine_unit ninexnine_unit_1907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13602)
);

assign C1602=c10602+c11602+c12602+c13602;
assign A1602=(C1602>=0)?1:0;

ninexnine_unit ninexnine_unit_1908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10612)
);

ninexnine_unit ninexnine_unit_1909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11612)
);

ninexnine_unit ninexnine_unit_1910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12612)
);

ninexnine_unit ninexnine_unit_1911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13612)
);

assign C1612=c10612+c11612+c12612+c13612;
assign A1612=(C1612>=0)?1:0;

ninexnine_unit ninexnine_unit_1912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10622)
);

ninexnine_unit ninexnine_unit_1913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11622)
);

ninexnine_unit ninexnine_unit_1914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12622)
);

ninexnine_unit ninexnine_unit_1915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13622)
);

assign C1622=c10622+c11622+c12622+c13622;
assign A1622=(C1622>=0)?1:0;

ninexnine_unit ninexnine_unit_1916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10632)
);

ninexnine_unit ninexnine_unit_1917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11632)
);

ninexnine_unit ninexnine_unit_1918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12632)
);

ninexnine_unit ninexnine_unit_1919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13632)
);

assign C1632=c10632+c11632+c12632+c13632;
assign A1632=(C1632>=0)?1:0;

ninexnine_unit ninexnine_unit_1920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10642)
);

ninexnine_unit ninexnine_unit_1921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11642)
);

ninexnine_unit ninexnine_unit_1922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12642)
);

ninexnine_unit ninexnine_unit_1923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13642)
);

assign C1642=c10642+c11642+c12642+c13642;
assign A1642=(C1642>=0)?1:0;

ninexnine_unit ninexnine_unit_1924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10652)
);

ninexnine_unit ninexnine_unit_1925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11652)
);

ninexnine_unit ninexnine_unit_1926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12652)
);

ninexnine_unit ninexnine_unit_1927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13652)
);

assign C1652=c10652+c11652+c12652+c13652;
assign A1652=(C1652>=0)?1:0;

ninexnine_unit ninexnine_unit_1928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10662)
);

ninexnine_unit ninexnine_unit_1929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11662)
);

ninexnine_unit ninexnine_unit_1930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12662)
);

ninexnine_unit ninexnine_unit_1931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13662)
);

assign C1662=c10662+c11662+c12662+c13662;
assign A1662=(C1662>=0)?1:0;

ninexnine_unit ninexnine_unit_1932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10672)
);

ninexnine_unit ninexnine_unit_1933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11672)
);

ninexnine_unit ninexnine_unit_1934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12672)
);

ninexnine_unit ninexnine_unit_1935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13672)
);

assign C1672=c10672+c11672+c12672+c13672;
assign A1672=(C1672>=0)?1:0;

ninexnine_unit ninexnine_unit_1936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10682)
);

ninexnine_unit ninexnine_unit_1937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11682)
);

ninexnine_unit ninexnine_unit_1938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12682)
);

ninexnine_unit ninexnine_unit_1939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13682)
);

assign C1682=c10682+c11682+c12682+c13682;
assign A1682=(C1682>=0)?1:0;

ninexnine_unit ninexnine_unit_1940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10692)
);

ninexnine_unit ninexnine_unit_1941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11692)
);

ninexnine_unit ninexnine_unit_1942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12692)
);

ninexnine_unit ninexnine_unit_1943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13692)
);

assign C1692=c10692+c11692+c12692+c13692;
assign A1692=(C1692>=0)?1:0;

ninexnine_unit ninexnine_unit_1944(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c106A2)
);

ninexnine_unit ninexnine_unit_1945(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c116A2)
);

ninexnine_unit ninexnine_unit_1946(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c126A2)
);

ninexnine_unit ninexnine_unit_1947(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c136A2)
);

assign C16A2=c106A2+c116A2+c126A2+c136A2;
assign A16A2=(C16A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1948(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c106B2)
);

ninexnine_unit ninexnine_unit_1949(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c116B2)
);

ninexnine_unit ninexnine_unit_1950(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c126B2)
);

ninexnine_unit ninexnine_unit_1951(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c136B2)
);

assign C16B2=c106B2+c116B2+c126B2+c136B2;
assign A16B2=(C16B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1952(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c106C2)
);

ninexnine_unit ninexnine_unit_1953(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c116C2)
);

ninexnine_unit ninexnine_unit_1954(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c126C2)
);

ninexnine_unit ninexnine_unit_1955(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c136C2)
);

assign C16C2=c106C2+c116C2+c126C2+c136C2;
assign A16C2=(C16C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1956(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c106D2)
);

ninexnine_unit ninexnine_unit_1957(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c116D2)
);

ninexnine_unit ninexnine_unit_1958(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c126D2)
);

ninexnine_unit ninexnine_unit_1959(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c136D2)
);

assign C16D2=c106D2+c116D2+c126D2+c136D2;
assign A16D2=(C16D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10702)
);

ninexnine_unit ninexnine_unit_1961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11702)
);

ninexnine_unit ninexnine_unit_1962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12702)
);

ninexnine_unit ninexnine_unit_1963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13702)
);

assign C1702=c10702+c11702+c12702+c13702;
assign A1702=(C1702>=0)?1:0;

ninexnine_unit ninexnine_unit_1964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10712)
);

ninexnine_unit ninexnine_unit_1965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11712)
);

ninexnine_unit ninexnine_unit_1966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12712)
);

ninexnine_unit ninexnine_unit_1967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13712)
);

assign C1712=c10712+c11712+c12712+c13712;
assign A1712=(C1712>=0)?1:0;

ninexnine_unit ninexnine_unit_1968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10722)
);

ninexnine_unit ninexnine_unit_1969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11722)
);

ninexnine_unit ninexnine_unit_1970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12722)
);

ninexnine_unit ninexnine_unit_1971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13722)
);

assign C1722=c10722+c11722+c12722+c13722;
assign A1722=(C1722>=0)?1:0;

ninexnine_unit ninexnine_unit_1972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10732)
);

ninexnine_unit ninexnine_unit_1973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11732)
);

ninexnine_unit ninexnine_unit_1974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12732)
);

ninexnine_unit ninexnine_unit_1975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13732)
);

assign C1732=c10732+c11732+c12732+c13732;
assign A1732=(C1732>=0)?1:0;

ninexnine_unit ninexnine_unit_1976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10742)
);

ninexnine_unit ninexnine_unit_1977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11742)
);

ninexnine_unit ninexnine_unit_1978(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12742)
);

ninexnine_unit ninexnine_unit_1979(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13742)
);

assign C1742=c10742+c11742+c12742+c13742;
assign A1742=(C1742>=0)?1:0;

ninexnine_unit ninexnine_unit_1980(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10752)
);

ninexnine_unit ninexnine_unit_1981(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11752)
);

ninexnine_unit ninexnine_unit_1982(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12752)
);

ninexnine_unit ninexnine_unit_1983(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13752)
);

assign C1752=c10752+c11752+c12752+c13752;
assign A1752=(C1752>=0)?1:0;

ninexnine_unit ninexnine_unit_1984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10762)
);

ninexnine_unit ninexnine_unit_1985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11762)
);

ninexnine_unit ninexnine_unit_1986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12762)
);

ninexnine_unit ninexnine_unit_1987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13762)
);

assign C1762=c10762+c11762+c12762+c13762;
assign A1762=(C1762>=0)?1:0;

ninexnine_unit ninexnine_unit_1988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10772)
);

ninexnine_unit ninexnine_unit_1989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11772)
);

ninexnine_unit ninexnine_unit_1990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12772)
);

ninexnine_unit ninexnine_unit_1991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13772)
);

assign C1772=c10772+c11772+c12772+c13772;
assign A1772=(C1772>=0)?1:0;

ninexnine_unit ninexnine_unit_1992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10782)
);

ninexnine_unit ninexnine_unit_1993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11782)
);

ninexnine_unit ninexnine_unit_1994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12782)
);

ninexnine_unit ninexnine_unit_1995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13782)
);

assign C1782=c10782+c11782+c12782+c13782;
assign A1782=(C1782>=0)?1:0;

ninexnine_unit ninexnine_unit_1996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10792)
);

ninexnine_unit ninexnine_unit_1997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11792)
);

ninexnine_unit ninexnine_unit_1998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12792)
);

ninexnine_unit ninexnine_unit_1999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13792)
);

assign C1792=c10792+c11792+c12792+c13792;
assign A1792=(C1792>=0)?1:0;

ninexnine_unit ninexnine_unit_2000(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c107A2)
);

ninexnine_unit ninexnine_unit_2001(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c117A2)
);

ninexnine_unit ninexnine_unit_2002(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c127A2)
);

ninexnine_unit ninexnine_unit_2003(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c137A2)
);

assign C17A2=c107A2+c117A2+c127A2+c137A2;
assign A17A2=(C17A2>=0)?1:0;

ninexnine_unit ninexnine_unit_2004(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c107B2)
);

ninexnine_unit ninexnine_unit_2005(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c117B2)
);

ninexnine_unit ninexnine_unit_2006(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c127B2)
);

ninexnine_unit ninexnine_unit_2007(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c137B2)
);

assign C17B2=c107B2+c117B2+c127B2+c137B2;
assign A17B2=(C17B2>=0)?1:0;

ninexnine_unit ninexnine_unit_2008(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c107C2)
);

ninexnine_unit ninexnine_unit_2009(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c117C2)
);

ninexnine_unit ninexnine_unit_2010(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c127C2)
);

ninexnine_unit ninexnine_unit_2011(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c137C2)
);

assign C17C2=c107C2+c117C2+c127C2+c137C2;
assign A17C2=(C17C2>=0)?1:0;

ninexnine_unit ninexnine_unit_2012(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c107D2)
);

ninexnine_unit ninexnine_unit_2013(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c117D2)
);

ninexnine_unit ninexnine_unit_2014(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c127D2)
);

ninexnine_unit ninexnine_unit_2015(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c137D2)
);

assign C17D2=c107D2+c117D2+c127D2+c137D2;
assign A17D2=(C17D2>=0)?1:0;

ninexnine_unit ninexnine_unit_2016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10802)
);

ninexnine_unit ninexnine_unit_2017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11802)
);

ninexnine_unit ninexnine_unit_2018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12802)
);

ninexnine_unit ninexnine_unit_2019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13802)
);

assign C1802=c10802+c11802+c12802+c13802;
assign A1802=(C1802>=0)?1:0;

ninexnine_unit ninexnine_unit_2020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10812)
);

ninexnine_unit ninexnine_unit_2021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11812)
);

ninexnine_unit ninexnine_unit_2022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12812)
);

ninexnine_unit ninexnine_unit_2023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13812)
);

assign C1812=c10812+c11812+c12812+c13812;
assign A1812=(C1812>=0)?1:0;

ninexnine_unit ninexnine_unit_2024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10822)
);

ninexnine_unit ninexnine_unit_2025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11822)
);

ninexnine_unit ninexnine_unit_2026(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12822)
);

ninexnine_unit ninexnine_unit_2027(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13822)
);

assign C1822=c10822+c11822+c12822+c13822;
assign A1822=(C1822>=0)?1:0;

ninexnine_unit ninexnine_unit_2028(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10832)
);

ninexnine_unit ninexnine_unit_2029(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11832)
);

ninexnine_unit ninexnine_unit_2030(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12832)
);

ninexnine_unit ninexnine_unit_2031(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13832)
);

assign C1832=c10832+c11832+c12832+c13832;
assign A1832=(C1832>=0)?1:0;

ninexnine_unit ninexnine_unit_2032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10842)
);

ninexnine_unit ninexnine_unit_2033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11842)
);

ninexnine_unit ninexnine_unit_2034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12842)
);

ninexnine_unit ninexnine_unit_2035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13842)
);

assign C1842=c10842+c11842+c12842+c13842;
assign A1842=(C1842>=0)?1:0;

ninexnine_unit ninexnine_unit_2036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10852)
);

ninexnine_unit ninexnine_unit_2037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11852)
);

ninexnine_unit ninexnine_unit_2038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12852)
);

ninexnine_unit ninexnine_unit_2039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13852)
);

assign C1852=c10852+c11852+c12852+c13852;
assign A1852=(C1852>=0)?1:0;

ninexnine_unit ninexnine_unit_2040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10862)
);

ninexnine_unit ninexnine_unit_2041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11862)
);

ninexnine_unit ninexnine_unit_2042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12862)
);

ninexnine_unit ninexnine_unit_2043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13862)
);

assign C1862=c10862+c11862+c12862+c13862;
assign A1862=(C1862>=0)?1:0;

ninexnine_unit ninexnine_unit_2044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10872)
);

ninexnine_unit ninexnine_unit_2045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11872)
);

ninexnine_unit ninexnine_unit_2046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12872)
);

ninexnine_unit ninexnine_unit_2047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13872)
);

assign C1872=c10872+c11872+c12872+c13872;
assign A1872=(C1872>=0)?1:0;

ninexnine_unit ninexnine_unit_2048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10882)
);

ninexnine_unit ninexnine_unit_2049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11882)
);

ninexnine_unit ninexnine_unit_2050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12882)
);

ninexnine_unit ninexnine_unit_2051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13882)
);

assign C1882=c10882+c11882+c12882+c13882;
assign A1882=(C1882>=0)?1:0;

ninexnine_unit ninexnine_unit_2052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10892)
);

ninexnine_unit ninexnine_unit_2053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11892)
);

ninexnine_unit ninexnine_unit_2054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12892)
);

ninexnine_unit ninexnine_unit_2055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13892)
);

assign C1892=c10892+c11892+c12892+c13892;
assign A1892=(C1892>=0)?1:0;

ninexnine_unit ninexnine_unit_2056(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c108A2)
);

ninexnine_unit ninexnine_unit_2057(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c118A2)
);

ninexnine_unit ninexnine_unit_2058(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c128A2)
);

ninexnine_unit ninexnine_unit_2059(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c138A2)
);

assign C18A2=c108A2+c118A2+c128A2+c138A2;
assign A18A2=(C18A2>=0)?1:0;

ninexnine_unit ninexnine_unit_2060(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c108B2)
);

ninexnine_unit ninexnine_unit_2061(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c118B2)
);

ninexnine_unit ninexnine_unit_2062(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c128B2)
);

ninexnine_unit ninexnine_unit_2063(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c138B2)
);

assign C18B2=c108B2+c118B2+c128B2+c138B2;
assign A18B2=(C18B2>=0)?1:0;

ninexnine_unit ninexnine_unit_2064(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c108C2)
);

ninexnine_unit ninexnine_unit_2065(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c118C2)
);

ninexnine_unit ninexnine_unit_2066(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c128C2)
);

ninexnine_unit ninexnine_unit_2067(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c138C2)
);

assign C18C2=c108C2+c118C2+c128C2+c138C2;
assign A18C2=(C18C2>=0)?1:0;

ninexnine_unit ninexnine_unit_2068(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c108D2)
);

ninexnine_unit ninexnine_unit_2069(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c118D2)
);

ninexnine_unit ninexnine_unit_2070(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c128D2)
);

ninexnine_unit ninexnine_unit_2071(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c138D2)
);

assign C18D2=c108D2+c118D2+c128D2+c138D2;
assign A18D2=(C18D2>=0)?1:0;

ninexnine_unit ninexnine_unit_2072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10902)
);

ninexnine_unit ninexnine_unit_2073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11902)
);

ninexnine_unit ninexnine_unit_2074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12902)
);

ninexnine_unit ninexnine_unit_2075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13902)
);

assign C1902=c10902+c11902+c12902+c13902;
assign A1902=(C1902>=0)?1:0;

ninexnine_unit ninexnine_unit_2076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10912)
);

ninexnine_unit ninexnine_unit_2077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11912)
);

ninexnine_unit ninexnine_unit_2078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12912)
);

ninexnine_unit ninexnine_unit_2079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13912)
);

assign C1912=c10912+c11912+c12912+c13912;
assign A1912=(C1912>=0)?1:0;

ninexnine_unit ninexnine_unit_2080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10922)
);

ninexnine_unit ninexnine_unit_2081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11922)
);

ninexnine_unit ninexnine_unit_2082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12922)
);

ninexnine_unit ninexnine_unit_2083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13922)
);

assign C1922=c10922+c11922+c12922+c13922;
assign A1922=(C1922>=0)?1:0;

ninexnine_unit ninexnine_unit_2084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10932)
);

ninexnine_unit ninexnine_unit_2085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11932)
);

ninexnine_unit ninexnine_unit_2086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12932)
);

ninexnine_unit ninexnine_unit_2087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13932)
);

assign C1932=c10932+c11932+c12932+c13932;
assign A1932=(C1932>=0)?1:0;

ninexnine_unit ninexnine_unit_2088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10942)
);

ninexnine_unit ninexnine_unit_2089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11942)
);

ninexnine_unit ninexnine_unit_2090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12942)
);

ninexnine_unit ninexnine_unit_2091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13942)
);

assign C1942=c10942+c11942+c12942+c13942;
assign A1942=(C1942>=0)?1:0;

ninexnine_unit ninexnine_unit_2092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10952)
);

ninexnine_unit ninexnine_unit_2093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11952)
);

ninexnine_unit ninexnine_unit_2094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12952)
);

ninexnine_unit ninexnine_unit_2095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13952)
);

assign C1952=c10952+c11952+c12952+c13952;
assign A1952=(C1952>=0)?1:0;

ninexnine_unit ninexnine_unit_2096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10962)
);

ninexnine_unit ninexnine_unit_2097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11962)
);

ninexnine_unit ninexnine_unit_2098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12962)
);

ninexnine_unit ninexnine_unit_2099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13962)
);

assign C1962=c10962+c11962+c12962+c13962;
assign A1962=(C1962>=0)?1:0;

ninexnine_unit ninexnine_unit_2100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10972)
);

ninexnine_unit ninexnine_unit_2101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11972)
);

ninexnine_unit ninexnine_unit_2102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12972)
);

ninexnine_unit ninexnine_unit_2103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13972)
);

assign C1972=c10972+c11972+c12972+c13972;
assign A1972=(C1972>=0)?1:0;

ninexnine_unit ninexnine_unit_2104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10982)
);

ninexnine_unit ninexnine_unit_2105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11982)
);

ninexnine_unit ninexnine_unit_2106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12982)
);

ninexnine_unit ninexnine_unit_2107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13982)
);

assign C1982=c10982+c11982+c12982+c13982;
assign A1982=(C1982>=0)?1:0;

ninexnine_unit ninexnine_unit_2108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10992)
);

ninexnine_unit ninexnine_unit_2109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11992)
);

ninexnine_unit ninexnine_unit_2110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12992)
);

ninexnine_unit ninexnine_unit_2111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13992)
);

assign C1992=c10992+c11992+c12992+c13992;
assign A1992=(C1992>=0)?1:0;

ninexnine_unit ninexnine_unit_2112(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c109A2)
);

ninexnine_unit ninexnine_unit_2113(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c119A2)
);

ninexnine_unit ninexnine_unit_2114(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c129A2)
);

ninexnine_unit ninexnine_unit_2115(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c139A2)
);

assign C19A2=c109A2+c119A2+c129A2+c139A2;
assign A19A2=(C19A2>=0)?1:0;

ninexnine_unit ninexnine_unit_2116(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c109B2)
);

ninexnine_unit ninexnine_unit_2117(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c119B2)
);

ninexnine_unit ninexnine_unit_2118(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c129B2)
);

ninexnine_unit ninexnine_unit_2119(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c139B2)
);

assign C19B2=c109B2+c119B2+c129B2+c139B2;
assign A19B2=(C19B2>=0)?1:0;

ninexnine_unit ninexnine_unit_2120(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c109C2)
);

ninexnine_unit ninexnine_unit_2121(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c119C2)
);

ninexnine_unit ninexnine_unit_2122(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c129C2)
);

ninexnine_unit ninexnine_unit_2123(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c139C2)
);

assign C19C2=c109C2+c119C2+c129C2+c139C2;
assign A19C2=(C19C2>=0)?1:0;

ninexnine_unit ninexnine_unit_2124(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c109D2)
);

ninexnine_unit ninexnine_unit_2125(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c119D2)
);

ninexnine_unit ninexnine_unit_2126(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c129D2)
);

ninexnine_unit ninexnine_unit_2127(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c139D2)
);

assign C19D2=c109D2+c119D2+c129D2+c139D2;
assign A19D2=(C19D2>=0)?1:0;

ninexnine_unit ninexnine_unit_2128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A02)
);

ninexnine_unit ninexnine_unit_2129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A02)
);

ninexnine_unit ninexnine_unit_2130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A02)
);

ninexnine_unit ninexnine_unit_2131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A02)
);

assign C1A02=c10A02+c11A02+c12A02+c13A02;
assign A1A02=(C1A02>=0)?1:0;

ninexnine_unit ninexnine_unit_2132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A12)
);

ninexnine_unit ninexnine_unit_2133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A12)
);

ninexnine_unit ninexnine_unit_2134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A12)
);

ninexnine_unit ninexnine_unit_2135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A12)
);

assign C1A12=c10A12+c11A12+c12A12+c13A12;
assign A1A12=(C1A12>=0)?1:0;

ninexnine_unit ninexnine_unit_2136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A22)
);

ninexnine_unit ninexnine_unit_2137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A22)
);

ninexnine_unit ninexnine_unit_2138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A22)
);

ninexnine_unit ninexnine_unit_2139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A22)
);

assign C1A22=c10A22+c11A22+c12A22+c13A22;
assign A1A22=(C1A22>=0)?1:0;

ninexnine_unit ninexnine_unit_2140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A32)
);

ninexnine_unit ninexnine_unit_2141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A32)
);

ninexnine_unit ninexnine_unit_2142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A32)
);

ninexnine_unit ninexnine_unit_2143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A32)
);

assign C1A32=c10A32+c11A32+c12A32+c13A32;
assign A1A32=(C1A32>=0)?1:0;

ninexnine_unit ninexnine_unit_2144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A42)
);

ninexnine_unit ninexnine_unit_2145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A42)
);

ninexnine_unit ninexnine_unit_2146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A42)
);

ninexnine_unit ninexnine_unit_2147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A42)
);

assign C1A42=c10A42+c11A42+c12A42+c13A42;
assign A1A42=(C1A42>=0)?1:0;

ninexnine_unit ninexnine_unit_2148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A52)
);

ninexnine_unit ninexnine_unit_2149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A52)
);

ninexnine_unit ninexnine_unit_2150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A52)
);

ninexnine_unit ninexnine_unit_2151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A52)
);

assign C1A52=c10A52+c11A52+c12A52+c13A52;
assign A1A52=(C1A52>=0)?1:0;

ninexnine_unit ninexnine_unit_2152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A62)
);

ninexnine_unit ninexnine_unit_2153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A62)
);

ninexnine_unit ninexnine_unit_2154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A62)
);

ninexnine_unit ninexnine_unit_2155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A62)
);

assign C1A62=c10A62+c11A62+c12A62+c13A62;
assign A1A62=(C1A62>=0)?1:0;

ninexnine_unit ninexnine_unit_2156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A72)
);

ninexnine_unit ninexnine_unit_2157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A72)
);

ninexnine_unit ninexnine_unit_2158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A72)
);

ninexnine_unit ninexnine_unit_2159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A72)
);

assign C1A72=c10A72+c11A72+c12A72+c13A72;
assign A1A72=(C1A72>=0)?1:0;

ninexnine_unit ninexnine_unit_2160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A82)
);

ninexnine_unit ninexnine_unit_2161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A82)
);

ninexnine_unit ninexnine_unit_2162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A82)
);

ninexnine_unit ninexnine_unit_2163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A82)
);

assign C1A82=c10A82+c11A82+c12A82+c13A82;
assign A1A82=(C1A82>=0)?1:0;

ninexnine_unit ninexnine_unit_2164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10A92)
);

ninexnine_unit ninexnine_unit_2165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11A92)
);

ninexnine_unit ninexnine_unit_2166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12A92)
);

ninexnine_unit ninexnine_unit_2167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13A92)
);

assign C1A92=c10A92+c11A92+c12A92+c13A92;
assign A1A92=(C1A92>=0)?1:0;

ninexnine_unit ninexnine_unit_2168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10AA2)
);

ninexnine_unit ninexnine_unit_2169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11AA2)
);

ninexnine_unit ninexnine_unit_2170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12AA2)
);

ninexnine_unit ninexnine_unit_2171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13AA2)
);

assign C1AA2=c10AA2+c11AA2+c12AA2+c13AA2;
assign A1AA2=(C1AA2>=0)?1:0;

ninexnine_unit ninexnine_unit_2172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10AB2)
);

ninexnine_unit ninexnine_unit_2173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11AB2)
);

ninexnine_unit ninexnine_unit_2174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12AB2)
);

ninexnine_unit ninexnine_unit_2175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13AB2)
);

assign C1AB2=c10AB2+c11AB2+c12AB2+c13AB2;
assign A1AB2=(C1AB2>=0)?1:0;

ninexnine_unit ninexnine_unit_2176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10AC2)
);

ninexnine_unit ninexnine_unit_2177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11AC2)
);

ninexnine_unit ninexnine_unit_2178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12AC2)
);

ninexnine_unit ninexnine_unit_2179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13AC2)
);

assign C1AC2=c10AC2+c11AC2+c12AC2+c13AC2;
assign A1AC2=(C1AC2>=0)?1:0;

ninexnine_unit ninexnine_unit_2180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10AD2)
);

ninexnine_unit ninexnine_unit_2181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11AD2)
);

ninexnine_unit ninexnine_unit_2182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12AD2)
);

ninexnine_unit ninexnine_unit_2183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13AD2)
);

assign C1AD2=c10AD2+c11AD2+c12AD2+c13AD2;
assign A1AD2=(C1AD2>=0)?1:0;

ninexnine_unit ninexnine_unit_2184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B02)
);

ninexnine_unit ninexnine_unit_2185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B02)
);

ninexnine_unit ninexnine_unit_2186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B02)
);

ninexnine_unit ninexnine_unit_2187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B02)
);

assign C1B02=c10B02+c11B02+c12B02+c13B02;
assign A1B02=(C1B02>=0)?1:0;

ninexnine_unit ninexnine_unit_2188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B12)
);

ninexnine_unit ninexnine_unit_2189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B12)
);

ninexnine_unit ninexnine_unit_2190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B12)
);

ninexnine_unit ninexnine_unit_2191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B12)
);

assign C1B12=c10B12+c11B12+c12B12+c13B12;
assign A1B12=(C1B12>=0)?1:0;

ninexnine_unit ninexnine_unit_2192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B22)
);

ninexnine_unit ninexnine_unit_2193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B22)
);

ninexnine_unit ninexnine_unit_2194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B22)
);

ninexnine_unit ninexnine_unit_2195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B22)
);

assign C1B22=c10B22+c11B22+c12B22+c13B22;
assign A1B22=(C1B22>=0)?1:0;

ninexnine_unit ninexnine_unit_2196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B32)
);

ninexnine_unit ninexnine_unit_2197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B32)
);

ninexnine_unit ninexnine_unit_2198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B32)
);

ninexnine_unit ninexnine_unit_2199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B32)
);

assign C1B32=c10B32+c11B32+c12B32+c13B32;
assign A1B32=(C1B32>=0)?1:0;

ninexnine_unit ninexnine_unit_2200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B42)
);

ninexnine_unit ninexnine_unit_2201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B42)
);

ninexnine_unit ninexnine_unit_2202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B42)
);

ninexnine_unit ninexnine_unit_2203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B42)
);

assign C1B42=c10B42+c11B42+c12B42+c13B42;
assign A1B42=(C1B42>=0)?1:0;

ninexnine_unit ninexnine_unit_2204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B52)
);

ninexnine_unit ninexnine_unit_2205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B52)
);

ninexnine_unit ninexnine_unit_2206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B52)
);

ninexnine_unit ninexnine_unit_2207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B52)
);

assign C1B52=c10B52+c11B52+c12B52+c13B52;
assign A1B52=(C1B52>=0)?1:0;

ninexnine_unit ninexnine_unit_2208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B62)
);

ninexnine_unit ninexnine_unit_2209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B62)
);

ninexnine_unit ninexnine_unit_2210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B62)
);

ninexnine_unit ninexnine_unit_2211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B62)
);

assign C1B62=c10B62+c11B62+c12B62+c13B62;
assign A1B62=(C1B62>=0)?1:0;

ninexnine_unit ninexnine_unit_2212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B72)
);

ninexnine_unit ninexnine_unit_2213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B72)
);

ninexnine_unit ninexnine_unit_2214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B72)
);

ninexnine_unit ninexnine_unit_2215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B72)
);

assign C1B72=c10B72+c11B72+c12B72+c13B72;
assign A1B72=(C1B72>=0)?1:0;

ninexnine_unit ninexnine_unit_2216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B82)
);

ninexnine_unit ninexnine_unit_2217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B82)
);

ninexnine_unit ninexnine_unit_2218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B82)
);

ninexnine_unit ninexnine_unit_2219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B82)
);

assign C1B82=c10B82+c11B82+c12B82+c13B82;
assign A1B82=(C1B82>=0)?1:0;

ninexnine_unit ninexnine_unit_2220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10B92)
);

ninexnine_unit ninexnine_unit_2221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11B92)
);

ninexnine_unit ninexnine_unit_2222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12B92)
);

ninexnine_unit ninexnine_unit_2223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13B92)
);

assign C1B92=c10B92+c11B92+c12B92+c13B92;
assign A1B92=(C1B92>=0)?1:0;

ninexnine_unit ninexnine_unit_2224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10BA2)
);

ninexnine_unit ninexnine_unit_2225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11BA2)
);

ninexnine_unit ninexnine_unit_2226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12BA2)
);

ninexnine_unit ninexnine_unit_2227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13BA2)
);

assign C1BA2=c10BA2+c11BA2+c12BA2+c13BA2;
assign A1BA2=(C1BA2>=0)?1:0;

ninexnine_unit ninexnine_unit_2228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10BB2)
);

ninexnine_unit ninexnine_unit_2229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11BB2)
);

ninexnine_unit ninexnine_unit_2230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12BB2)
);

ninexnine_unit ninexnine_unit_2231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13BB2)
);

assign C1BB2=c10BB2+c11BB2+c12BB2+c13BB2;
assign A1BB2=(C1BB2>=0)?1:0;

ninexnine_unit ninexnine_unit_2232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10BC2)
);

ninexnine_unit ninexnine_unit_2233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11BC2)
);

ninexnine_unit ninexnine_unit_2234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12BC2)
);

ninexnine_unit ninexnine_unit_2235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13BC2)
);

assign C1BC2=c10BC2+c11BC2+c12BC2+c13BC2;
assign A1BC2=(C1BC2>=0)?1:0;

ninexnine_unit ninexnine_unit_2236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10BD2)
);

ninexnine_unit ninexnine_unit_2237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11BD2)
);

ninexnine_unit ninexnine_unit_2238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12BD2)
);

ninexnine_unit ninexnine_unit_2239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13BD2)
);

assign C1BD2=c10BD2+c11BD2+c12BD2+c13BD2;
assign A1BD2=(C1BD2>=0)?1:0;

ninexnine_unit ninexnine_unit_2240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C02)
);

ninexnine_unit ninexnine_unit_2241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C02)
);

ninexnine_unit ninexnine_unit_2242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C02)
);

ninexnine_unit ninexnine_unit_2243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C02)
);

assign C1C02=c10C02+c11C02+c12C02+c13C02;
assign A1C02=(C1C02>=0)?1:0;

ninexnine_unit ninexnine_unit_2244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C12)
);

ninexnine_unit ninexnine_unit_2245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C12)
);

ninexnine_unit ninexnine_unit_2246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C12)
);

ninexnine_unit ninexnine_unit_2247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C12)
);

assign C1C12=c10C12+c11C12+c12C12+c13C12;
assign A1C12=(C1C12>=0)?1:0;

ninexnine_unit ninexnine_unit_2248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C22)
);

ninexnine_unit ninexnine_unit_2249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C22)
);

ninexnine_unit ninexnine_unit_2250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C22)
);

ninexnine_unit ninexnine_unit_2251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C22)
);

assign C1C22=c10C22+c11C22+c12C22+c13C22;
assign A1C22=(C1C22>=0)?1:0;

ninexnine_unit ninexnine_unit_2252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C32)
);

ninexnine_unit ninexnine_unit_2253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C32)
);

ninexnine_unit ninexnine_unit_2254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C32)
);

ninexnine_unit ninexnine_unit_2255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C32)
);

assign C1C32=c10C32+c11C32+c12C32+c13C32;
assign A1C32=(C1C32>=0)?1:0;

ninexnine_unit ninexnine_unit_2256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C42)
);

ninexnine_unit ninexnine_unit_2257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C42)
);

ninexnine_unit ninexnine_unit_2258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C42)
);

ninexnine_unit ninexnine_unit_2259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C42)
);

assign C1C42=c10C42+c11C42+c12C42+c13C42;
assign A1C42=(C1C42>=0)?1:0;

ninexnine_unit ninexnine_unit_2260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C52)
);

ninexnine_unit ninexnine_unit_2261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C52)
);

ninexnine_unit ninexnine_unit_2262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C52)
);

ninexnine_unit ninexnine_unit_2263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C52)
);

assign C1C52=c10C52+c11C52+c12C52+c13C52;
assign A1C52=(C1C52>=0)?1:0;

ninexnine_unit ninexnine_unit_2264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C62)
);

ninexnine_unit ninexnine_unit_2265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C62)
);

ninexnine_unit ninexnine_unit_2266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C62)
);

ninexnine_unit ninexnine_unit_2267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C62)
);

assign C1C62=c10C62+c11C62+c12C62+c13C62;
assign A1C62=(C1C62>=0)?1:0;

ninexnine_unit ninexnine_unit_2268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C72)
);

ninexnine_unit ninexnine_unit_2269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C72)
);

ninexnine_unit ninexnine_unit_2270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C72)
);

ninexnine_unit ninexnine_unit_2271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C72)
);

assign C1C72=c10C72+c11C72+c12C72+c13C72;
assign A1C72=(C1C72>=0)?1:0;

ninexnine_unit ninexnine_unit_2272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C82)
);

ninexnine_unit ninexnine_unit_2273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C82)
);

ninexnine_unit ninexnine_unit_2274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C82)
);

ninexnine_unit ninexnine_unit_2275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C82)
);

assign C1C82=c10C82+c11C82+c12C82+c13C82;
assign A1C82=(C1C82>=0)?1:0;

ninexnine_unit ninexnine_unit_2276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10C92)
);

ninexnine_unit ninexnine_unit_2277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11C92)
);

ninexnine_unit ninexnine_unit_2278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12C92)
);

ninexnine_unit ninexnine_unit_2279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13C92)
);

assign C1C92=c10C92+c11C92+c12C92+c13C92;
assign A1C92=(C1C92>=0)?1:0;

ninexnine_unit ninexnine_unit_2280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10CA2)
);

ninexnine_unit ninexnine_unit_2281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11CA2)
);

ninexnine_unit ninexnine_unit_2282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12CA2)
);

ninexnine_unit ninexnine_unit_2283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13CA2)
);

assign C1CA2=c10CA2+c11CA2+c12CA2+c13CA2;
assign A1CA2=(C1CA2>=0)?1:0;

ninexnine_unit ninexnine_unit_2284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10CB2)
);

ninexnine_unit ninexnine_unit_2285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11CB2)
);

ninexnine_unit ninexnine_unit_2286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12CB2)
);

ninexnine_unit ninexnine_unit_2287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13CB2)
);

assign C1CB2=c10CB2+c11CB2+c12CB2+c13CB2;
assign A1CB2=(C1CB2>=0)?1:0;

ninexnine_unit ninexnine_unit_2288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10CC2)
);

ninexnine_unit ninexnine_unit_2289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11CC2)
);

ninexnine_unit ninexnine_unit_2290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12CC2)
);

ninexnine_unit ninexnine_unit_2291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13CC2)
);

assign C1CC2=c10CC2+c11CC2+c12CC2+c13CC2;
assign A1CC2=(C1CC2>=0)?1:0;

ninexnine_unit ninexnine_unit_2292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10CD2)
);

ninexnine_unit ninexnine_unit_2293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11CD2)
);

ninexnine_unit ninexnine_unit_2294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12CD2)
);

ninexnine_unit ninexnine_unit_2295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13CD2)
);

assign C1CD2=c10CD2+c11CD2+c12CD2+c13CD2;
assign A1CD2=(C1CD2>=0)?1:0;

ninexnine_unit ninexnine_unit_2296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D02)
);

ninexnine_unit ninexnine_unit_2297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D02)
);

ninexnine_unit ninexnine_unit_2298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D02)
);

ninexnine_unit ninexnine_unit_2299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D02)
);

assign C1D02=c10D02+c11D02+c12D02+c13D02;
assign A1D02=(C1D02>=0)?1:0;

ninexnine_unit ninexnine_unit_2300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D12)
);

ninexnine_unit ninexnine_unit_2301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D12)
);

ninexnine_unit ninexnine_unit_2302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D12)
);

ninexnine_unit ninexnine_unit_2303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D12)
);

assign C1D12=c10D12+c11D12+c12D12+c13D12;
assign A1D12=(C1D12>=0)?1:0;

ninexnine_unit ninexnine_unit_2304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D22)
);

ninexnine_unit ninexnine_unit_2305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D22)
);

ninexnine_unit ninexnine_unit_2306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D22)
);

ninexnine_unit ninexnine_unit_2307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D22)
);

assign C1D22=c10D22+c11D22+c12D22+c13D22;
assign A1D22=(C1D22>=0)?1:0;

ninexnine_unit ninexnine_unit_2308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D32)
);

ninexnine_unit ninexnine_unit_2309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D32)
);

ninexnine_unit ninexnine_unit_2310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D32)
);

ninexnine_unit ninexnine_unit_2311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D32)
);

assign C1D32=c10D32+c11D32+c12D32+c13D32;
assign A1D32=(C1D32>=0)?1:0;

ninexnine_unit ninexnine_unit_2312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D42)
);

ninexnine_unit ninexnine_unit_2313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D42)
);

ninexnine_unit ninexnine_unit_2314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D42)
);

ninexnine_unit ninexnine_unit_2315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D42)
);

assign C1D42=c10D42+c11D42+c12D42+c13D42;
assign A1D42=(C1D42>=0)?1:0;

ninexnine_unit ninexnine_unit_2316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D52)
);

ninexnine_unit ninexnine_unit_2317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D52)
);

ninexnine_unit ninexnine_unit_2318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D52)
);

ninexnine_unit ninexnine_unit_2319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D52)
);

assign C1D52=c10D52+c11D52+c12D52+c13D52;
assign A1D52=(C1D52>=0)?1:0;

ninexnine_unit ninexnine_unit_2320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D62)
);

ninexnine_unit ninexnine_unit_2321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D62)
);

ninexnine_unit ninexnine_unit_2322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D62)
);

ninexnine_unit ninexnine_unit_2323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D62)
);

assign C1D62=c10D62+c11D62+c12D62+c13D62;
assign A1D62=(C1D62>=0)?1:0;

ninexnine_unit ninexnine_unit_2324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D72)
);

ninexnine_unit ninexnine_unit_2325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D72)
);

ninexnine_unit ninexnine_unit_2326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D72)
);

ninexnine_unit ninexnine_unit_2327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D72)
);

assign C1D72=c10D72+c11D72+c12D72+c13D72;
assign A1D72=(C1D72>=0)?1:0;

ninexnine_unit ninexnine_unit_2328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D82)
);

ninexnine_unit ninexnine_unit_2329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D82)
);

ninexnine_unit ninexnine_unit_2330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D82)
);

ninexnine_unit ninexnine_unit_2331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D82)
);

assign C1D82=c10D82+c11D82+c12D82+c13D82;
assign A1D82=(C1D82>=0)?1:0;

ninexnine_unit ninexnine_unit_2332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10D92)
);

ninexnine_unit ninexnine_unit_2333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11D92)
);

ninexnine_unit ninexnine_unit_2334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12D92)
);

ninexnine_unit ninexnine_unit_2335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13D92)
);

assign C1D92=c10D92+c11D92+c12D92+c13D92;
assign A1D92=(C1D92>=0)?1:0;

ninexnine_unit ninexnine_unit_2336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10DA2)
);

ninexnine_unit ninexnine_unit_2337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11DA2)
);

ninexnine_unit ninexnine_unit_2338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12DA2)
);

ninexnine_unit ninexnine_unit_2339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13DA2)
);

assign C1DA2=c10DA2+c11DA2+c12DA2+c13DA2;
assign A1DA2=(C1DA2>=0)?1:0;

ninexnine_unit ninexnine_unit_2340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10DB2)
);

ninexnine_unit ninexnine_unit_2341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11DB2)
);

ninexnine_unit ninexnine_unit_2342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12DB2)
);

ninexnine_unit ninexnine_unit_2343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13DB2)
);

assign C1DB2=c10DB2+c11DB2+c12DB2+c13DB2;
assign A1DB2=(C1DB2>=0)?1:0;

ninexnine_unit ninexnine_unit_2344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10DC2)
);

ninexnine_unit ninexnine_unit_2345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11DC2)
);

ninexnine_unit ninexnine_unit_2346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12DC2)
);

ninexnine_unit ninexnine_unit_2347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13DC2)
);

assign C1DC2=c10DC2+c11DC2+c12DC2+c13DC2;
assign A1DC2=(C1DC2>=0)?1:0;

ninexnine_unit ninexnine_unit_2348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10DD2)
);

ninexnine_unit ninexnine_unit_2349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11DD2)
);

ninexnine_unit ninexnine_unit_2350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12DD2)
);

ninexnine_unit ninexnine_unit_2351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13DD2)
);

assign C1DD2=c10DD2+c11DD2+c12DD2+c13DD2;
assign A1DD2=(C1DD2>=0)?1:0;

ninexnine_unit ninexnine_unit_2352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10003)
);

ninexnine_unit ninexnine_unit_2353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11003)
);

ninexnine_unit ninexnine_unit_2354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12003)
);

ninexnine_unit ninexnine_unit_2355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13003)
);

assign C1003=c10003+c11003+c12003+c13003;
assign A1003=(C1003>=0)?1:0;

ninexnine_unit ninexnine_unit_2356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10013)
);

ninexnine_unit ninexnine_unit_2357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11013)
);

ninexnine_unit ninexnine_unit_2358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12013)
);

ninexnine_unit ninexnine_unit_2359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13013)
);

assign C1013=c10013+c11013+c12013+c13013;
assign A1013=(C1013>=0)?1:0;

ninexnine_unit ninexnine_unit_2360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10023)
);

ninexnine_unit ninexnine_unit_2361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11023)
);

ninexnine_unit ninexnine_unit_2362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12023)
);

ninexnine_unit ninexnine_unit_2363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13023)
);

assign C1023=c10023+c11023+c12023+c13023;
assign A1023=(C1023>=0)?1:0;

ninexnine_unit ninexnine_unit_2364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10033)
);

ninexnine_unit ninexnine_unit_2365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11033)
);

ninexnine_unit ninexnine_unit_2366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12033)
);

ninexnine_unit ninexnine_unit_2367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13033)
);

assign C1033=c10033+c11033+c12033+c13033;
assign A1033=(C1033>=0)?1:0;

ninexnine_unit ninexnine_unit_2368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10043)
);

ninexnine_unit ninexnine_unit_2369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11043)
);

ninexnine_unit ninexnine_unit_2370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12043)
);

ninexnine_unit ninexnine_unit_2371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13043)
);

assign C1043=c10043+c11043+c12043+c13043;
assign A1043=(C1043>=0)?1:0;

ninexnine_unit ninexnine_unit_2372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10053)
);

ninexnine_unit ninexnine_unit_2373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11053)
);

ninexnine_unit ninexnine_unit_2374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12053)
);

ninexnine_unit ninexnine_unit_2375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13053)
);

assign C1053=c10053+c11053+c12053+c13053;
assign A1053=(C1053>=0)?1:0;

ninexnine_unit ninexnine_unit_2376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10063)
);

ninexnine_unit ninexnine_unit_2377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11063)
);

ninexnine_unit ninexnine_unit_2378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12063)
);

ninexnine_unit ninexnine_unit_2379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13063)
);

assign C1063=c10063+c11063+c12063+c13063;
assign A1063=(C1063>=0)?1:0;

ninexnine_unit ninexnine_unit_2380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10073)
);

ninexnine_unit ninexnine_unit_2381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11073)
);

ninexnine_unit ninexnine_unit_2382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12073)
);

ninexnine_unit ninexnine_unit_2383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13073)
);

assign C1073=c10073+c11073+c12073+c13073;
assign A1073=(C1073>=0)?1:0;

ninexnine_unit ninexnine_unit_2384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10083)
);

ninexnine_unit ninexnine_unit_2385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11083)
);

ninexnine_unit ninexnine_unit_2386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12083)
);

ninexnine_unit ninexnine_unit_2387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13083)
);

assign C1083=c10083+c11083+c12083+c13083;
assign A1083=(C1083>=0)?1:0;

ninexnine_unit ninexnine_unit_2388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10093)
);

ninexnine_unit ninexnine_unit_2389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11093)
);

ninexnine_unit ninexnine_unit_2390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12093)
);

ninexnine_unit ninexnine_unit_2391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13093)
);

assign C1093=c10093+c11093+c12093+c13093;
assign A1093=(C1093>=0)?1:0;

ninexnine_unit ninexnine_unit_2392(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c100A3)
);

ninexnine_unit ninexnine_unit_2393(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c110A3)
);

ninexnine_unit ninexnine_unit_2394(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c120A3)
);

ninexnine_unit ninexnine_unit_2395(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c130A3)
);

assign C10A3=c100A3+c110A3+c120A3+c130A3;
assign A10A3=(C10A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2396(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c100B3)
);

ninexnine_unit ninexnine_unit_2397(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c110B3)
);

ninexnine_unit ninexnine_unit_2398(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c120B3)
);

ninexnine_unit ninexnine_unit_2399(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c130B3)
);

assign C10B3=c100B3+c110B3+c120B3+c130B3;
assign A10B3=(C10B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2400(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c100C3)
);

ninexnine_unit ninexnine_unit_2401(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c110C3)
);

ninexnine_unit ninexnine_unit_2402(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c120C3)
);

ninexnine_unit ninexnine_unit_2403(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c130C3)
);

assign C10C3=c100C3+c110C3+c120C3+c130C3;
assign A10C3=(C10C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2404(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c100D3)
);

ninexnine_unit ninexnine_unit_2405(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c110D3)
);

ninexnine_unit ninexnine_unit_2406(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c120D3)
);

ninexnine_unit ninexnine_unit_2407(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c130D3)
);

assign C10D3=c100D3+c110D3+c120D3+c130D3;
assign A10D3=(C10D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10103)
);

ninexnine_unit ninexnine_unit_2409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11103)
);

ninexnine_unit ninexnine_unit_2410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12103)
);

ninexnine_unit ninexnine_unit_2411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13103)
);

assign C1103=c10103+c11103+c12103+c13103;
assign A1103=(C1103>=0)?1:0;

ninexnine_unit ninexnine_unit_2412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10113)
);

ninexnine_unit ninexnine_unit_2413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11113)
);

ninexnine_unit ninexnine_unit_2414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12113)
);

ninexnine_unit ninexnine_unit_2415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13113)
);

assign C1113=c10113+c11113+c12113+c13113;
assign A1113=(C1113>=0)?1:0;

ninexnine_unit ninexnine_unit_2416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10123)
);

ninexnine_unit ninexnine_unit_2417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11123)
);

ninexnine_unit ninexnine_unit_2418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12123)
);

ninexnine_unit ninexnine_unit_2419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13123)
);

assign C1123=c10123+c11123+c12123+c13123;
assign A1123=(C1123>=0)?1:0;

ninexnine_unit ninexnine_unit_2420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10133)
);

ninexnine_unit ninexnine_unit_2421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11133)
);

ninexnine_unit ninexnine_unit_2422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12133)
);

ninexnine_unit ninexnine_unit_2423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13133)
);

assign C1133=c10133+c11133+c12133+c13133;
assign A1133=(C1133>=0)?1:0;

ninexnine_unit ninexnine_unit_2424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10143)
);

ninexnine_unit ninexnine_unit_2425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11143)
);

ninexnine_unit ninexnine_unit_2426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12143)
);

ninexnine_unit ninexnine_unit_2427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13143)
);

assign C1143=c10143+c11143+c12143+c13143;
assign A1143=(C1143>=0)?1:0;

ninexnine_unit ninexnine_unit_2428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10153)
);

ninexnine_unit ninexnine_unit_2429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11153)
);

ninexnine_unit ninexnine_unit_2430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12153)
);

ninexnine_unit ninexnine_unit_2431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13153)
);

assign C1153=c10153+c11153+c12153+c13153;
assign A1153=(C1153>=0)?1:0;

ninexnine_unit ninexnine_unit_2432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10163)
);

ninexnine_unit ninexnine_unit_2433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11163)
);

ninexnine_unit ninexnine_unit_2434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12163)
);

ninexnine_unit ninexnine_unit_2435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13163)
);

assign C1163=c10163+c11163+c12163+c13163;
assign A1163=(C1163>=0)?1:0;

ninexnine_unit ninexnine_unit_2436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10173)
);

ninexnine_unit ninexnine_unit_2437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11173)
);

ninexnine_unit ninexnine_unit_2438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12173)
);

ninexnine_unit ninexnine_unit_2439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13173)
);

assign C1173=c10173+c11173+c12173+c13173;
assign A1173=(C1173>=0)?1:0;

ninexnine_unit ninexnine_unit_2440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10183)
);

ninexnine_unit ninexnine_unit_2441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11183)
);

ninexnine_unit ninexnine_unit_2442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12183)
);

ninexnine_unit ninexnine_unit_2443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13183)
);

assign C1183=c10183+c11183+c12183+c13183;
assign A1183=(C1183>=0)?1:0;

ninexnine_unit ninexnine_unit_2444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10193)
);

ninexnine_unit ninexnine_unit_2445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11193)
);

ninexnine_unit ninexnine_unit_2446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12193)
);

ninexnine_unit ninexnine_unit_2447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13193)
);

assign C1193=c10193+c11193+c12193+c13193;
assign A1193=(C1193>=0)?1:0;

ninexnine_unit ninexnine_unit_2448(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c101A3)
);

ninexnine_unit ninexnine_unit_2449(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c111A3)
);

ninexnine_unit ninexnine_unit_2450(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c121A3)
);

ninexnine_unit ninexnine_unit_2451(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c131A3)
);

assign C11A3=c101A3+c111A3+c121A3+c131A3;
assign A11A3=(C11A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2452(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c101B3)
);

ninexnine_unit ninexnine_unit_2453(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c111B3)
);

ninexnine_unit ninexnine_unit_2454(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c121B3)
);

ninexnine_unit ninexnine_unit_2455(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c131B3)
);

assign C11B3=c101B3+c111B3+c121B3+c131B3;
assign A11B3=(C11B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2456(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c101C3)
);

ninexnine_unit ninexnine_unit_2457(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c111C3)
);

ninexnine_unit ninexnine_unit_2458(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c121C3)
);

ninexnine_unit ninexnine_unit_2459(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c131C3)
);

assign C11C3=c101C3+c111C3+c121C3+c131C3;
assign A11C3=(C11C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2460(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c101D3)
);

ninexnine_unit ninexnine_unit_2461(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c111D3)
);

ninexnine_unit ninexnine_unit_2462(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c121D3)
);

ninexnine_unit ninexnine_unit_2463(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c131D3)
);

assign C11D3=c101D3+c111D3+c121D3+c131D3;
assign A11D3=(C11D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10203)
);

ninexnine_unit ninexnine_unit_2465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11203)
);

ninexnine_unit ninexnine_unit_2466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12203)
);

ninexnine_unit ninexnine_unit_2467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13203)
);

assign C1203=c10203+c11203+c12203+c13203;
assign A1203=(C1203>=0)?1:0;

ninexnine_unit ninexnine_unit_2468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10213)
);

ninexnine_unit ninexnine_unit_2469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11213)
);

ninexnine_unit ninexnine_unit_2470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12213)
);

ninexnine_unit ninexnine_unit_2471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13213)
);

assign C1213=c10213+c11213+c12213+c13213;
assign A1213=(C1213>=0)?1:0;

ninexnine_unit ninexnine_unit_2472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10223)
);

ninexnine_unit ninexnine_unit_2473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11223)
);

ninexnine_unit ninexnine_unit_2474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12223)
);

ninexnine_unit ninexnine_unit_2475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13223)
);

assign C1223=c10223+c11223+c12223+c13223;
assign A1223=(C1223>=0)?1:0;

ninexnine_unit ninexnine_unit_2476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10233)
);

ninexnine_unit ninexnine_unit_2477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11233)
);

ninexnine_unit ninexnine_unit_2478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12233)
);

ninexnine_unit ninexnine_unit_2479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13233)
);

assign C1233=c10233+c11233+c12233+c13233;
assign A1233=(C1233>=0)?1:0;

ninexnine_unit ninexnine_unit_2480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10243)
);

ninexnine_unit ninexnine_unit_2481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11243)
);

ninexnine_unit ninexnine_unit_2482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12243)
);

ninexnine_unit ninexnine_unit_2483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13243)
);

assign C1243=c10243+c11243+c12243+c13243;
assign A1243=(C1243>=0)?1:0;

ninexnine_unit ninexnine_unit_2484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10253)
);

ninexnine_unit ninexnine_unit_2485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11253)
);

ninexnine_unit ninexnine_unit_2486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12253)
);

ninexnine_unit ninexnine_unit_2487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13253)
);

assign C1253=c10253+c11253+c12253+c13253;
assign A1253=(C1253>=0)?1:0;

ninexnine_unit ninexnine_unit_2488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10263)
);

ninexnine_unit ninexnine_unit_2489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11263)
);

ninexnine_unit ninexnine_unit_2490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12263)
);

ninexnine_unit ninexnine_unit_2491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13263)
);

assign C1263=c10263+c11263+c12263+c13263;
assign A1263=(C1263>=0)?1:0;

ninexnine_unit ninexnine_unit_2492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10273)
);

ninexnine_unit ninexnine_unit_2493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11273)
);

ninexnine_unit ninexnine_unit_2494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12273)
);

ninexnine_unit ninexnine_unit_2495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13273)
);

assign C1273=c10273+c11273+c12273+c13273;
assign A1273=(C1273>=0)?1:0;

ninexnine_unit ninexnine_unit_2496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10283)
);

ninexnine_unit ninexnine_unit_2497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11283)
);

ninexnine_unit ninexnine_unit_2498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12283)
);

ninexnine_unit ninexnine_unit_2499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13283)
);

assign C1283=c10283+c11283+c12283+c13283;
assign A1283=(C1283>=0)?1:0;

ninexnine_unit ninexnine_unit_2500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10293)
);

ninexnine_unit ninexnine_unit_2501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11293)
);

ninexnine_unit ninexnine_unit_2502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12293)
);

ninexnine_unit ninexnine_unit_2503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13293)
);

assign C1293=c10293+c11293+c12293+c13293;
assign A1293=(C1293>=0)?1:0;

ninexnine_unit ninexnine_unit_2504(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c102A3)
);

ninexnine_unit ninexnine_unit_2505(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c112A3)
);

ninexnine_unit ninexnine_unit_2506(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c122A3)
);

ninexnine_unit ninexnine_unit_2507(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c132A3)
);

assign C12A3=c102A3+c112A3+c122A3+c132A3;
assign A12A3=(C12A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2508(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c102B3)
);

ninexnine_unit ninexnine_unit_2509(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c112B3)
);

ninexnine_unit ninexnine_unit_2510(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c122B3)
);

ninexnine_unit ninexnine_unit_2511(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c132B3)
);

assign C12B3=c102B3+c112B3+c122B3+c132B3;
assign A12B3=(C12B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2512(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c102C3)
);

ninexnine_unit ninexnine_unit_2513(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c112C3)
);

ninexnine_unit ninexnine_unit_2514(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c122C3)
);

ninexnine_unit ninexnine_unit_2515(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c132C3)
);

assign C12C3=c102C3+c112C3+c122C3+c132C3;
assign A12C3=(C12C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2516(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c102D3)
);

ninexnine_unit ninexnine_unit_2517(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c112D3)
);

ninexnine_unit ninexnine_unit_2518(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c122D3)
);

ninexnine_unit ninexnine_unit_2519(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c132D3)
);

assign C12D3=c102D3+c112D3+c122D3+c132D3;
assign A12D3=(C12D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10303)
);

ninexnine_unit ninexnine_unit_2521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11303)
);

ninexnine_unit ninexnine_unit_2522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12303)
);

ninexnine_unit ninexnine_unit_2523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13303)
);

assign C1303=c10303+c11303+c12303+c13303;
assign A1303=(C1303>=0)?1:0;

ninexnine_unit ninexnine_unit_2524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10313)
);

ninexnine_unit ninexnine_unit_2525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11313)
);

ninexnine_unit ninexnine_unit_2526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12313)
);

ninexnine_unit ninexnine_unit_2527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13313)
);

assign C1313=c10313+c11313+c12313+c13313;
assign A1313=(C1313>=0)?1:0;

ninexnine_unit ninexnine_unit_2528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10323)
);

ninexnine_unit ninexnine_unit_2529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11323)
);

ninexnine_unit ninexnine_unit_2530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12323)
);

ninexnine_unit ninexnine_unit_2531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13323)
);

assign C1323=c10323+c11323+c12323+c13323;
assign A1323=(C1323>=0)?1:0;

ninexnine_unit ninexnine_unit_2532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10333)
);

ninexnine_unit ninexnine_unit_2533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11333)
);

ninexnine_unit ninexnine_unit_2534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12333)
);

ninexnine_unit ninexnine_unit_2535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13333)
);

assign C1333=c10333+c11333+c12333+c13333;
assign A1333=(C1333>=0)?1:0;

ninexnine_unit ninexnine_unit_2536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10343)
);

ninexnine_unit ninexnine_unit_2537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11343)
);

ninexnine_unit ninexnine_unit_2538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12343)
);

ninexnine_unit ninexnine_unit_2539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13343)
);

assign C1343=c10343+c11343+c12343+c13343;
assign A1343=(C1343>=0)?1:0;

ninexnine_unit ninexnine_unit_2540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10353)
);

ninexnine_unit ninexnine_unit_2541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11353)
);

ninexnine_unit ninexnine_unit_2542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12353)
);

ninexnine_unit ninexnine_unit_2543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13353)
);

assign C1353=c10353+c11353+c12353+c13353;
assign A1353=(C1353>=0)?1:0;

ninexnine_unit ninexnine_unit_2544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10363)
);

ninexnine_unit ninexnine_unit_2545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11363)
);

ninexnine_unit ninexnine_unit_2546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12363)
);

ninexnine_unit ninexnine_unit_2547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13363)
);

assign C1363=c10363+c11363+c12363+c13363;
assign A1363=(C1363>=0)?1:0;

ninexnine_unit ninexnine_unit_2548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10373)
);

ninexnine_unit ninexnine_unit_2549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11373)
);

ninexnine_unit ninexnine_unit_2550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12373)
);

ninexnine_unit ninexnine_unit_2551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13373)
);

assign C1373=c10373+c11373+c12373+c13373;
assign A1373=(C1373>=0)?1:0;

ninexnine_unit ninexnine_unit_2552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10383)
);

ninexnine_unit ninexnine_unit_2553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11383)
);

ninexnine_unit ninexnine_unit_2554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12383)
);

ninexnine_unit ninexnine_unit_2555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13383)
);

assign C1383=c10383+c11383+c12383+c13383;
assign A1383=(C1383>=0)?1:0;

ninexnine_unit ninexnine_unit_2556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10393)
);

ninexnine_unit ninexnine_unit_2557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11393)
);

ninexnine_unit ninexnine_unit_2558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12393)
);

ninexnine_unit ninexnine_unit_2559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13393)
);

assign C1393=c10393+c11393+c12393+c13393;
assign A1393=(C1393>=0)?1:0;

ninexnine_unit ninexnine_unit_2560(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c103A3)
);

ninexnine_unit ninexnine_unit_2561(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c113A3)
);

ninexnine_unit ninexnine_unit_2562(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c123A3)
);

ninexnine_unit ninexnine_unit_2563(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c133A3)
);

assign C13A3=c103A3+c113A3+c123A3+c133A3;
assign A13A3=(C13A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2564(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c103B3)
);

ninexnine_unit ninexnine_unit_2565(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c113B3)
);

ninexnine_unit ninexnine_unit_2566(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c123B3)
);

ninexnine_unit ninexnine_unit_2567(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c133B3)
);

assign C13B3=c103B3+c113B3+c123B3+c133B3;
assign A13B3=(C13B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2568(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c103C3)
);

ninexnine_unit ninexnine_unit_2569(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c113C3)
);

ninexnine_unit ninexnine_unit_2570(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c123C3)
);

ninexnine_unit ninexnine_unit_2571(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c133C3)
);

assign C13C3=c103C3+c113C3+c123C3+c133C3;
assign A13C3=(C13C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2572(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c103D3)
);

ninexnine_unit ninexnine_unit_2573(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c113D3)
);

ninexnine_unit ninexnine_unit_2574(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c123D3)
);

ninexnine_unit ninexnine_unit_2575(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c133D3)
);

assign C13D3=c103D3+c113D3+c123D3+c133D3;
assign A13D3=(C13D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10403)
);

ninexnine_unit ninexnine_unit_2577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11403)
);

ninexnine_unit ninexnine_unit_2578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12403)
);

ninexnine_unit ninexnine_unit_2579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13403)
);

assign C1403=c10403+c11403+c12403+c13403;
assign A1403=(C1403>=0)?1:0;

ninexnine_unit ninexnine_unit_2580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10413)
);

ninexnine_unit ninexnine_unit_2581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11413)
);

ninexnine_unit ninexnine_unit_2582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12413)
);

ninexnine_unit ninexnine_unit_2583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13413)
);

assign C1413=c10413+c11413+c12413+c13413;
assign A1413=(C1413>=0)?1:0;

ninexnine_unit ninexnine_unit_2584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10423)
);

ninexnine_unit ninexnine_unit_2585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11423)
);

ninexnine_unit ninexnine_unit_2586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12423)
);

ninexnine_unit ninexnine_unit_2587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13423)
);

assign C1423=c10423+c11423+c12423+c13423;
assign A1423=(C1423>=0)?1:0;

ninexnine_unit ninexnine_unit_2588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10433)
);

ninexnine_unit ninexnine_unit_2589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11433)
);

ninexnine_unit ninexnine_unit_2590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12433)
);

ninexnine_unit ninexnine_unit_2591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13433)
);

assign C1433=c10433+c11433+c12433+c13433;
assign A1433=(C1433>=0)?1:0;

ninexnine_unit ninexnine_unit_2592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10443)
);

ninexnine_unit ninexnine_unit_2593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11443)
);

ninexnine_unit ninexnine_unit_2594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12443)
);

ninexnine_unit ninexnine_unit_2595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13443)
);

assign C1443=c10443+c11443+c12443+c13443;
assign A1443=(C1443>=0)?1:0;

ninexnine_unit ninexnine_unit_2596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10453)
);

ninexnine_unit ninexnine_unit_2597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11453)
);

ninexnine_unit ninexnine_unit_2598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12453)
);

ninexnine_unit ninexnine_unit_2599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13453)
);

assign C1453=c10453+c11453+c12453+c13453;
assign A1453=(C1453>=0)?1:0;

ninexnine_unit ninexnine_unit_2600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10463)
);

ninexnine_unit ninexnine_unit_2601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11463)
);

ninexnine_unit ninexnine_unit_2602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12463)
);

ninexnine_unit ninexnine_unit_2603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13463)
);

assign C1463=c10463+c11463+c12463+c13463;
assign A1463=(C1463>=0)?1:0;

ninexnine_unit ninexnine_unit_2604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10473)
);

ninexnine_unit ninexnine_unit_2605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11473)
);

ninexnine_unit ninexnine_unit_2606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12473)
);

ninexnine_unit ninexnine_unit_2607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13473)
);

assign C1473=c10473+c11473+c12473+c13473;
assign A1473=(C1473>=0)?1:0;

ninexnine_unit ninexnine_unit_2608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10483)
);

ninexnine_unit ninexnine_unit_2609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11483)
);

ninexnine_unit ninexnine_unit_2610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12483)
);

ninexnine_unit ninexnine_unit_2611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13483)
);

assign C1483=c10483+c11483+c12483+c13483;
assign A1483=(C1483>=0)?1:0;

ninexnine_unit ninexnine_unit_2612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10493)
);

ninexnine_unit ninexnine_unit_2613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11493)
);

ninexnine_unit ninexnine_unit_2614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12493)
);

ninexnine_unit ninexnine_unit_2615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13493)
);

assign C1493=c10493+c11493+c12493+c13493;
assign A1493=(C1493>=0)?1:0;

ninexnine_unit ninexnine_unit_2616(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c104A3)
);

ninexnine_unit ninexnine_unit_2617(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c114A3)
);

ninexnine_unit ninexnine_unit_2618(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c124A3)
);

ninexnine_unit ninexnine_unit_2619(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c134A3)
);

assign C14A3=c104A3+c114A3+c124A3+c134A3;
assign A14A3=(C14A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2620(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c104B3)
);

ninexnine_unit ninexnine_unit_2621(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c114B3)
);

ninexnine_unit ninexnine_unit_2622(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c124B3)
);

ninexnine_unit ninexnine_unit_2623(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c134B3)
);

assign C14B3=c104B3+c114B3+c124B3+c134B3;
assign A14B3=(C14B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2624(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c104C3)
);

ninexnine_unit ninexnine_unit_2625(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c114C3)
);

ninexnine_unit ninexnine_unit_2626(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c124C3)
);

ninexnine_unit ninexnine_unit_2627(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c134C3)
);

assign C14C3=c104C3+c114C3+c124C3+c134C3;
assign A14C3=(C14C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2628(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c104D3)
);

ninexnine_unit ninexnine_unit_2629(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c114D3)
);

ninexnine_unit ninexnine_unit_2630(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c124D3)
);

ninexnine_unit ninexnine_unit_2631(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c134D3)
);

assign C14D3=c104D3+c114D3+c124D3+c134D3;
assign A14D3=(C14D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10503)
);

ninexnine_unit ninexnine_unit_2633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11503)
);

ninexnine_unit ninexnine_unit_2634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12503)
);

ninexnine_unit ninexnine_unit_2635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13503)
);

assign C1503=c10503+c11503+c12503+c13503;
assign A1503=(C1503>=0)?1:0;

ninexnine_unit ninexnine_unit_2636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10513)
);

ninexnine_unit ninexnine_unit_2637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11513)
);

ninexnine_unit ninexnine_unit_2638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12513)
);

ninexnine_unit ninexnine_unit_2639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13513)
);

assign C1513=c10513+c11513+c12513+c13513;
assign A1513=(C1513>=0)?1:0;

ninexnine_unit ninexnine_unit_2640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10523)
);

ninexnine_unit ninexnine_unit_2641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11523)
);

ninexnine_unit ninexnine_unit_2642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12523)
);

ninexnine_unit ninexnine_unit_2643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13523)
);

assign C1523=c10523+c11523+c12523+c13523;
assign A1523=(C1523>=0)?1:0;

ninexnine_unit ninexnine_unit_2644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10533)
);

ninexnine_unit ninexnine_unit_2645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11533)
);

ninexnine_unit ninexnine_unit_2646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12533)
);

ninexnine_unit ninexnine_unit_2647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13533)
);

assign C1533=c10533+c11533+c12533+c13533;
assign A1533=(C1533>=0)?1:0;

ninexnine_unit ninexnine_unit_2648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10543)
);

ninexnine_unit ninexnine_unit_2649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11543)
);

ninexnine_unit ninexnine_unit_2650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12543)
);

ninexnine_unit ninexnine_unit_2651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13543)
);

assign C1543=c10543+c11543+c12543+c13543;
assign A1543=(C1543>=0)?1:0;

ninexnine_unit ninexnine_unit_2652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10553)
);

ninexnine_unit ninexnine_unit_2653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11553)
);

ninexnine_unit ninexnine_unit_2654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12553)
);

ninexnine_unit ninexnine_unit_2655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13553)
);

assign C1553=c10553+c11553+c12553+c13553;
assign A1553=(C1553>=0)?1:0;

ninexnine_unit ninexnine_unit_2656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10563)
);

ninexnine_unit ninexnine_unit_2657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11563)
);

ninexnine_unit ninexnine_unit_2658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12563)
);

ninexnine_unit ninexnine_unit_2659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13563)
);

assign C1563=c10563+c11563+c12563+c13563;
assign A1563=(C1563>=0)?1:0;

ninexnine_unit ninexnine_unit_2660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10573)
);

ninexnine_unit ninexnine_unit_2661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11573)
);

ninexnine_unit ninexnine_unit_2662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12573)
);

ninexnine_unit ninexnine_unit_2663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13573)
);

assign C1573=c10573+c11573+c12573+c13573;
assign A1573=(C1573>=0)?1:0;

ninexnine_unit ninexnine_unit_2664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10583)
);

ninexnine_unit ninexnine_unit_2665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11583)
);

ninexnine_unit ninexnine_unit_2666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12583)
);

ninexnine_unit ninexnine_unit_2667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13583)
);

assign C1583=c10583+c11583+c12583+c13583;
assign A1583=(C1583>=0)?1:0;

ninexnine_unit ninexnine_unit_2668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10593)
);

ninexnine_unit ninexnine_unit_2669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11593)
);

ninexnine_unit ninexnine_unit_2670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12593)
);

ninexnine_unit ninexnine_unit_2671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13593)
);

assign C1593=c10593+c11593+c12593+c13593;
assign A1593=(C1593>=0)?1:0;

ninexnine_unit ninexnine_unit_2672(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c105A3)
);

ninexnine_unit ninexnine_unit_2673(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c115A3)
);

ninexnine_unit ninexnine_unit_2674(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c125A3)
);

ninexnine_unit ninexnine_unit_2675(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c135A3)
);

assign C15A3=c105A3+c115A3+c125A3+c135A3;
assign A15A3=(C15A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2676(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c105B3)
);

ninexnine_unit ninexnine_unit_2677(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c115B3)
);

ninexnine_unit ninexnine_unit_2678(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c125B3)
);

ninexnine_unit ninexnine_unit_2679(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c135B3)
);

assign C15B3=c105B3+c115B3+c125B3+c135B3;
assign A15B3=(C15B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2680(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c105C3)
);

ninexnine_unit ninexnine_unit_2681(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c115C3)
);

ninexnine_unit ninexnine_unit_2682(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c125C3)
);

ninexnine_unit ninexnine_unit_2683(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c135C3)
);

assign C15C3=c105C3+c115C3+c125C3+c135C3;
assign A15C3=(C15C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2684(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c105D3)
);

ninexnine_unit ninexnine_unit_2685(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c115D3)
);

ninexnine_unit ninexnine_unit_2686(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c125D3)
);

ninexnine_unit ninexnine_unit_2687(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c135D3)
);

assign C15D3=c105D3+c115D3+c125D3+c135D3;
assign A15D3=(C15D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10603)
);

ninexnine_unit ninexnine_unit_2689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11603)
);

ninexnine_unit ninexnine_unit_2690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12603)
);

ninexnine_unit ninexnine_unit_2691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13603)
);

assign C1603=c10603+c11603+c12603+c13603;
assign A1603=(C1603>=0)?1:0;

ninexnine_unit ninexnine_unit_2692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10613)
);

ninexnine_unit ninexnine_unit_2693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11613)
);

ninexnine_unit ninexnine_unit_2694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12613)
);

ninexnine_unit ninexnine_unit_2695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13613)
);

assign C1613=c10613+c11613+c12613+c13613;
assign A1613=(C1613>=0)?1:0;

ninexnine_unit ninexnine_unit_2696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10623)
);

ninexnine_unit ninexnine_unit_2697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11623)
);

ninexnine_unit ninexnine_unit_2698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12623)
);

ninexnine_unit ninexnine_unit_2699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13623)
);

assign C1623=c10623+c11623+c12623+c13623;
assign A1623=(C1623>=0)?1:0;

ninexnine_unit ninexnine_unit_2700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10633)
);

ninexnine_unit ninexnine_unit_2701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11633)
);

ninexnine_unit ninexnine_unit_2702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12633)
);

ninexnine_unit ninexnine_unit_2703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13633)
);

assign C1633=c10633+c11633+c12633+c13633;
assign A1633=(C1633>=0)?1:0;

ninexnine_unit ninexnine_unit_2704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10643)
);

ninexnine_unit ninexnine_unit_2705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11643)
);

ninexnine_unit ninexnine_unit_2706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12643)
);

ninexnine_unit ninexnine_unit_2707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13643)
);

assign C1643=c10643+c11643+c12643+c13643;
assign A1643=(C1643>=0)?1:0;

ninexnine_unit ninexnine_unit_2708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10653)
);

ninexnine_unit ninexnine_unit_2709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11653)
);

ninexnine_unit ninexnine_unit_2710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12653)
);

ninexnine_unit ninexnine_unit_2711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13653)
);

assign C1653=c10653+c11653+c12653+c13653;
assign A1653=(C1653>=0)?1:0;

ninexnine_unit ninexnine_unit_2712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10663)
);

ninexnine_unit ninexnine_unit_2713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11663)
);

ninexnine_unit ninexnine_unit_2714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12663)
);

ninexnine_unit ninexnine_unit_2715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13663)
);

assign C1663=c10663+c11663+c12663+c13663;
assign A1663=(C1663>=0)?1:0;

ninexnine_unit ninexnine_unit_2716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10673)
);

ninexnine_unit ninexnine_unit_2717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11673)
);

ninexnine_unit ninexnine_unit_2718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12673)
);

ninexnine_unit ninexnine_unit_2719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13673)
);

assign C1673=c10673+c11673+c12673+c13673;
assign A1673=(C1673>=0)?1:0;

ninexnine_unit ninexnine_unit_2720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10683)
);

ninexnine_unit ninexnine_unit_2721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11683)
);

ninexnine_unit ninexnine_unit_2722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12683)
);

ninexnine_unit ninexnine_unit_2723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13683)
);

assign C1683=c10683+c11683+c12683+c13683;
assign A1683=(C1683>=0)?1:0;

ninexnine_unit ninexnine_unit_2724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10693)
);

ninexnine_unit ninexnine_unit_2725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11693)
);

ninexnine_unit ninexnine_unit_2726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12693)
);

ninexnine_unit ninexnine_unit_2727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13693)
);

assign C1693=c10693+c11693+c12693+c13693;
assign A1693=(C1693>=0)?1:0;

ninexnine_unit ninexnine_unit_2728(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c106A3)
);

ninexnine_unit ninexnine_unit_2729(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c116A3)
);

ninexnine_unit ninexnine_unit_2730(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c126A3)
);

ninexnine_unit ninexnine_unit_2731(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c136A3)
);

assign C16A3=c106A3+c116A3+c126A3+c136A3;
assign A16A3=(C16A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2732(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c106B3)
);

ninexnine_unit ninexnine_unit_2733(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c116B3)
);

ninexnine_unit ninexnine_unit_2734(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c126B3)
);

ninexnine_unit ninexnine_unit_2735(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c136B3)
);

assign C16B3=c106B3+c116B3+c126B3+c136B3;
assign A16B3=(C16B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2736(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c106C3)
);

ninexnine_unit ninexnine_unit_2737(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c116C3)
);

ninexnine_unit ninexnine_unit_2738(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c126C3)
);

ninexnine_unit ninexnine_unit_2739(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c136C3)
);

assign C16C3=c106C3+c116C3+c126C3+c136C3;
assign A16C3=(C16C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2740(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c106D3)
);

ninexnine_unit ninexnine_unit_2741(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c116D3)
);

ninexnine_unit ninexnine_unit_2742(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c126D3)
);

ninexnine_unit ninexnine_unit_2743(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c136D3)
);

assign C16D3=c106D3+c116D3+c126D3+c136D3;
assign A16D3=(C16D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10703)
);

ninexnine_unit ninexnine_unit_2745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11703)
);

ninexnine_unit ninexnine_unit_2746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12703)
);

ninexnine_unit ninexnine_unit_2747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13703)
);

assign C1703=c10703+c11703+c12703+c13703;
assign A1703=(C1703>=0)?1:0;

ninexnine_unit ninexnine_unit_2748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10713)
);

ninexnine_unit ninexnine_unit_2749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11713)
);

ninexnine_unit ninexnine_unit_2750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12713)
);

ninexnine_unit ninexnine_unit_2751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13713)
);

assign C1713=c10713+c11713+c12713+c13713;
assign A1713=(C1713>=0)?1:0;

ninexnine_unit ninexnine_unit_2752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10723)
);

ninexnine_unit ninexnine_unit_2753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11723)
);

ninexnine_unit ninexnine_unit_2754(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12723)
);

ninexnine_unit ninexnine_unit_2755(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13723)
);

assign C1723=c10723+c11723+c12723+c13723;
assign A1723=(C1723>=0)?1:0;

ninexnine_unit ninexnine_unit_2756(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10733)
);

ninexnine_unit ninexnine_unit_2757(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11733)
);

ninexnine_unit ninexnine_unit_2758(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12733)
);

ninexnine_unit ninexnine_unit_2759(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13733)
);

assign C1733=c10733+c11733+c12733+c13733;
assign A1733=(C1733>=0)?1:0;

ninexnine_unit ninexnine_unit_2760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10743)
);

ninexnine_unit ninexnine_unit_2761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11743)
);

ninexnine_unit ninexnine_unit_2762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12743)
);

ninexnine_unit ninexnine_unit_2763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13743)
);

assign C1743=c10743+c11743+c12743+c13743;
assign A1743=(C1743>=0)?1:0;

ninexnine_unit ninexnine_unit_2764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10753)
);

ninexnine_unit ninexnine_unit_2765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11753)
);

ninexnine_unit ninexnine_unit_2766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12753)
);

ninexnine_unit ninexnine_unit_2767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13753)
);

assign C1753=c10753+c11753+c12753+c13753;
assign A1753=(C1753>=0)?1:0;

ninexnine_unit ninexnine_unit_2768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10763)
);

ninexnine_unit ninexnine_unit_2769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11763)
);

ninexnine_unit ninexnine_unit_2770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12763)
);

ninexnine_unit ninexnine_unit_2771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13763)
);

assign C1763=c10763+c11763+c12763+c13763;
assign A1763=(C1763>=0)?1:0;

ninexnine_unit ninexnine_unit_2772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10773)
);

ninexnine_unit ninexnine_unit_2773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11773)
);

ninexnine_unit ninexnine_unit_2774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12773)
);

ninexnine_unit ninexnine_unit_2775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13773)
);

assign C1773=c10773+c11773+c12773+c13773;
assign A1773=(C1773>=0)?1:0;

ninexnine_unit ninexnine_unit_2776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10783)
);

ninexnine_unit ninexnine_unit_2777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11783)
);

ninexnine_unit ninexnine_unit_2778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12783)
);

ninexnine_unit ninexnine_unit_2779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13783)
);

assign C1783=c10783+c11783+c12783+c13783;
assign A1783=(C1783>=0)?1:0;

ninexnine_unit ninexnine_unit_2780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10793)
);

ninexnine_unit ninexnine_unit_2781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11793)
);

ninexnine_unit ninexnine_unit_2782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12793)
);

ninexnine_unit ninexnine_unit_2783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13793)
);

assign C1793=c10793+c11793+c12793+c13793;
assign A1793=(C1793>=0)?1:0;

ninexnine_unit ninexnine_unit_2784(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c107A3)
);

ninexnine_unit ninexnine_unit_2785(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c117A3)
);

ninexnine_unit ninexnine_unit_2786(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c127A3)
);

ninexnine_unit ninexnine_unit_2787(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c137A3)
);

assign C17A3=c107A3+c117A3+c127A3+c137A3;
assign A17A3=(C17A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2788(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c107B3)
);

ninexnine_unit ninexnine_unit_2789(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c117B3)
);

ninexnine_unit ninexnine_unit_2790(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c127B3)
);

ninexnine_unit ninexnine_unit_2791(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c137B3)
);

assign C17B3=c107B3+c117B3+c127B3+c137B3;
assign A17B3=(C17B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2792(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c107C3)
);

ninexnine_unit ninexnine_unit_2793(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c117C3)
);

ninexnine_unit ninexnine_unit_2794(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c127C3)
);

ninexnine_unit ninexnine_unit_2795(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c137C3)
);

assign C17C3=c107C3+c117C3+c127C3+c137C3;
assign A17C3=(C17C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2796(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c107D3)
);

ninexnine_unit ninexnine_unit_2797(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c117D3)
);

ninexnine_unit ninexnine_unit_2798(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c127D3)
);

ninexnine_unit ninexnine_unit_2799(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c137D3)
);

assign C17D3=c107D3+c117D3+c127D3+c137D3;
assign A17D3=(C17D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10803)
);

ninexnine_unit ninexnine_unit_2801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11803)
);

ninexnine_unit ninexnine_unit_2802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12803)
);

ninexnine_unit ninexnine_unit_2803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13803)
);

assign C1803=c10803+c11803+c12803+c13803;
assign A1803=(C1803>=0)?1:0;

ninexnine_unit ninexnine_unit_2804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10813)
);

ninexnine_unit ninexnine_unit_2805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11813)
);

ninexnine_unit ninexnine_unit_2806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12813)
);

ninexnine_unit ninexnine_unit_2807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13813)
);

assign C1813=c10813+c11813+c12813+c13813;
assign A1813=(C1813>=0)?1:0;

ninexnine_unit ninexnine_unit_2808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10823)
);

ninexnine_unit ninexnine_unit_2809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11823)
);

ninexnine_unit ninexnine_unit_2810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12823)
);

ninexnine_unit ninexnine_unit_2811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13823)
);

assign C1823=c10823+c11823+c12823+c13823;
assign A1823=(C1823>=0)?1:0;

ninexnine_unit ninexnine_unit_2812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10833)
);

ninexnine_unit ninexnine_unit_2813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11833)
);

ninexnine_unit ninexnine_unit_2814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12833)
);

ninexnine_unit ninexnine_unit_2815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13833)
);

assign C1833=c10833+c11833+c12833+c13833;
assign A1833=(C1833>=0)?1:0;

ninexnine_unit ninexnine_unit_2816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10843)
);

ninexnine_unit ninexnine_unit_2817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11843)
);

ninexnine_unit ninexnine_unit_2818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12843)
);

ninexnine_unit ninexnine_unit_2819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13843)
);

assign C1843=c10843+c11843+c12843+c13843;
assign A1843=(C1843>=0)?1:0;

ninexnine_unit ninexnine_unit_2820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10853)
);

ninexnine_unit ninexnine_unit_2821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11853)
);

ninexnine_unit ninexnine_unit_2822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12853)
);

ninexnine_unit ninexnine_unit_2823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13853)
);

assign C1853=c10853+c11853+c12853+c13853;
assign A1853=(C1853>=0)?1:0;

ninexnine_unit ninexnine_unit_2824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10863)
);

ninexnine_unit ninexnine_unit_2825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11863)
);

ninexnine_unit ninexnine_unit_2826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12863)
);

ninexnine_unit ninexnine_unit_2827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13863)
);

assign C1863=c10863+c11863+c12863+c13863;
assign A1863=(C1863>=0)?1:0;

ninexnine_unit ninexnine_unit_2828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10873)
);

ninexnine_unit ninexnine_unit_2829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11873)
);

ninexnine_unit ninexnine_unit_2830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12873)
);

ninexnine_unit ninexnine_unit_2831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13873)
);

assign C1873=c10873+c11873+c12873+c13873;
assign A1873=(C1873>=0)?1:0;

ninexnine_unit ninexnine_unit_2832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10883)
);

ninexnine_unit ninexnine_unit_2833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11883)
);

ninexnine_unit ninexnine_unit_2834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12883)
);

ninexnine_unit ninexnine_unit_2835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13883)
);

assign C1883=c10883+c11883+c12883+c13883;
assign A1883=(C1883>=0)?1:0;

ninexnine_unit ninexnine_unit_2836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10893)
);

ninexnine_unit ninexnine_unit_2837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11893)
);

ninexnine_unit ninexnine_unit_2838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12893)
);

ninexnine_unit ninexnine_unit_2839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13893)
);

assign C1893=c10893+c11893+c12893+c13893;
assign A1893=(C1893>=0)?1:0;

ninexnine_unit ninexnine_unit_2840(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c108A3)
);

ninexnine_unit ninexnine_unit_2841(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c118A3)
);

ninexnine_unit ninexnine_unit_2842(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c128A3)
);

ninexnine_unit ninexnine_unit_2843(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c138A3)
);

assign C18A3=c108A3+c118A3+c128A3+c138A3;
assign A18A3=(C18A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2844(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c108B3)
);

ninexnine_unit ninexnine_unit_2845(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c118B3)
);

ninexnine_unit ninexnine_unit_2846(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c128B3)
);

ninexnine_unit ninexnine_unit_2847(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c138B3)
);

assign C18B3=c108B3+c118B3+c128B3+c138B3;
assign A18B3=(C18B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2848(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c108C3)
);

ninexnine_unit ninexnine_unit_2849(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c118C3)
);

ninexnine_unit ninexnine_unit_2850(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c128C3)
);

ninexnine_unit ninexnine_unit_2851(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c138C3)
);

assign C18C3=c108C3+c118C3+c128C3+c138C3;
assign A18C3=(C18C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2852(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c108D3)
);

ninexnine_unit ninexnine_unit_2853(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c118D3)
);

ninexnine_unit ninexnine_unit_2854(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c128D3)
);

ninexnine_unit ninexnine_unit_2855(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c138D3)
);

assign C18D3=c108D3+c118D3+c128D3+c138D3;
assign A18D3=(C18D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10903)
);

ninexnine_unit ninexnine_unit_2857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11903)
);

ninexnine_unit ninexnine_unit_2858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12903)
);

ninexnine_unit ninexnine_unit_2859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13903)
);

assign C1903=c10903+c11903+c12903+c13903;
assign A1903=(C1903>=0)?1:0;

ninexnine_unit ninexnine_unit_2860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10913)
);

ninexnine_unit ninexnine_unit_2861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11913)
);

ninexnine_unit ninexnine_unit_2862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12913)
);

ninexnine_unit ninexnine_unit_2863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13913)
);

assign C1913=c10913+c11913+c12913+c13913;
assign A1913=(C1913>=0)?1:0;

ninexnine_unit ninexnine_unit_2864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10923)
);

ninexnine_unit ninexnine_unit_2865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11923)
);

ninexnine_unit ninexnine_unit_2866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12923)
);

ninexnine_unit ninexnine_unit_2867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13923)
);

assign C1923=c10923+c11923+c12923+c13923;
assign A1923=(C1923>=0)?1:0;

ninexnine_unit ninexnine_unit_2868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10933)
);

ninexnine_unit ninexnine_unit_2869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11933)
);

ninexnine_unit ninexnine_unit_2870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12933)
);

ninexnine_unit ninexnine_unit_2871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13933)
);

assign C1933=c10933+c11933+c12933+c13933;
assign A1933=(C1933>=0)?1:0;

ninexnine_unit ninexnine_unit_2872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10943)
);

ninexnine_unit ninexnine_unit_2873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11943)
);

ninexnine_unit ninexnine_unit_2874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12943)
);

ninexnine_unit ninexnine_unit_2875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13943)
);

assign C1943=c10943+c11943+c12943+c13943;
assign A1943=(C1943>=0)?1:0;

ninexnine_unit ninexnine_unit_2876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10953)
);

ninexnine_unit ninexnine_unit_2877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11953)
);

ninexnine_unit ninexnine_unit_2878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12953)
);

ninexnine_unit ninexnine_unit_2879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13953)
);

assign C1953=c10953+c11953+c12953+c13953;
assign A1953=(C1953>=0)?1:0;

ninexnine_unit ninexnine_unit_2880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10963)
);

ninexnine_unit ninexnine_unit_2881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11963)
);

ninexnine_unit ninexnine_unit_2882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12963)
);

ninexnine_unit ninexnine_unit_2883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13963)
);

assign C1963=c10963+c11963+c12963+c13963;
assign A1963=(C1963>=0)?1:0;

ninexnine_unit ninexnine_unit_2884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10973)
);

ninexnine_unit ninexnine_unit_2885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11973)
);

ninexnine_unit ninexnine_unit_2886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12973)
);

ninexnine_unit ninexnine_unit_2887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13973)
);

assign C1973=c10973+c11973+c12973+c13973;
assign A1973=(C1973>=0)?1:0;

ninexnine_unit ninexnine_unit_2888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10983)
);

ninexnine_unit ninexnine_unit_2889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11983)
);

ninexnine_unit ninexnine_unit_2890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12983)
);

ninexnine_unit ninexnine_unit_2891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13983)
);

assign C1983=c10983+c11983+c12983+c13983;
assign A1983=(C1983>=0)?1:0;

ninexnine_unit ninexnine_unit_2892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10993)
);

ninexnine_unit ninexnine_unit_2893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11993)
);

ninexnine_unit ninexnine_unit_2894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12993)
);

ninexnine_unit ninexnine_unit_2895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13993)
);

assign C1993=c10993+c11993+c12993+c13993;
assign A1993=(C1993>=0)?1:0;

ninexnine_unit ninexnine_unit_2896(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c109A3)
);

ninexnine_unit ninexnine_unit_2897(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c119A3)
);

ninexnine_unit ninexnine_unit_2898(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c129A3)
);

ninexnine_unit ninexnine_unit_2899(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c139A3)
);

assign C19A3=c109A3+c119A3+c129A3+c139A3;
assign A19A3=(C19A3>=0)?1:0;

ninexnine_unit ninexnine_unit_2900(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c109B3)
);

ninexnine_unit ninexnine_unit_2901(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c119B3)
);

ninexnine_unit ninexnine_unit_2902(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c129B3)
);

ninexnine_unit ninexnine_unit_2903(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c139B3)
);

assign C19B3=c109B3+c119B3+c129B3+c139B3;
assign A19B3=(C19B3>=0)?1:0;

ninexnine_unit ninexnine_unit_2904(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c109C3)
);

ninexnine_unit ninexnine_unit_2905(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c119C3)
);

ninexnine_unit ninexnine_unit_2906(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c129C3)
);

ninexnine_unit ninexnine_unit_2907(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c139C3)
);

assign C19C3=c109C3+c119C3+c129C3+c139C3;
assign A19C3=(C19C3>=0)?1:0;

ninexnine_unit ninexnine_unit_2908(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c109D3)
);

ninexnine_unit ninexnine_unit_2909(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c119D3)
);

ninexnine_unit ninexnine_unit_2910(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c129D3)
);

ninexnine_unit ninexnine_unit_2911(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c139D3)
);

assign C19D3=c109D3+c119D3+c129D3+c139D3;
assign A19D3=(C19D3>=0)?1:0;

ninexnine_unit ninexnine_unit_2912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A03)
);

ninexnine_unit ninexnine_unit_2913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A03)
);

ninexnine_unit ninexnine_unit_2914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A03)
);

ninexnine_unit ninexnine_unit_2915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A03)
);

assign C1A03=c10A03+c11A03+c12A03+c13A03;
assign A1A03=(C1A03>=0)?1:0;

ninexnine_unit ninexnine_unit_2916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A13)
);

ninexnine_unit ninexnine_unit_2917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A13)
);

ninexnine_unit ninexnine_unit_2918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A13)
);

ninexnine_unit ninexnine_unit_2919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A13)
);

assign C1A13=c10A13+c11A13+c12A13+c13A13;
assign A1A13=(C1A13>=0)?1:0;

ninexnine_unit ninexnine_unit_2920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A23)
);

ninexnine_unit ninexnine_unit_2921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A23)
);

ninexnine_unit ninexnine_unit_2922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A23)
);

ninexnine_unit ninexnine_unit_2923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A23)
);

assign C1A23=c10A23+c11A23+c12A23+c13A23;
assign A1A23=(C1A23>=0)?1:0;

ninexnine_unit ninexnine_unit_2924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A33)
);

ninexnine_unit ninexnine_unit_2925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A33)
);

ninexnine_unit ninexnine_unit_2926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A33)
);

ninexnine_unit ninexnine_unit_2927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A33)
);

assign C1A33=c10A33+c11A33+c12A33+c13A33;
assign A1A33=(C1A33>=0)?1:0;

ninexnine_unit ninexnine_unit_2928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A43)
);

ninexnine_unit ninexnine_unit_2929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A43)
);

ninexnine_unit ninexnine_unit_2930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A43)
);

ninexnine_unit ninexnine_unit_2931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A43)
);

assign C1A43=c10A43+c11A43+c12A43+c13A43;
assign A1A43=(C1A43>=0)?1:0;

ninexnine_unit ninexnine_unit_2932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A53)
);

ninexnine_unit ninexnine_unit_2933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A53)
);

ninexnine_unit ninexnine_unit_2934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A53)
);

ninexnine_unit ninexnine_unit_2935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A53)
);

assign C1A53=c10A53+c11A53+c12A53+c13A53;
assign A1A53=(C1A53>=0)?1:0;

ninexnine_unit ninexnine_unit_2936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A63)
);

ninexnine_unit ninexnine_unit_2937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A63)
);

ninexnine_unit ninexnine_unit_2938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A63)
);

ninexnine_unit ninexnine_unit_2939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A63)
);

assign C1A63=c10A63+c11A63+c12A63+c13A63;
assign A1A63=(C1A63>=0)?1:0;

ninexnine_unit ninexnine_unit_2940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A73)
);

ninexnine_unit ninexnine_unit_2941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A73)
);

ninexnine_unit ninexnine_unit_2942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A73)
);

ninexnine_unit ninexnine_unit_2943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A73)
);

assign C1A73=c10A73+c11A73+c12A73+c13A73;
assign A1A73=(C1A73>=0)?1:0;

ninexnine_unit ninexnine_unit_2944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A83)
);

ninexnine_unit ninexnine_unit_2945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A83)
);

ninexnine_unit ninexnine_unit_2946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A83)
);

ninexnine_unit ninexnine_unit_2947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A83)
);

assign C1A83=c10A83+c11A83+c12A83+c13A83;
assign A1A83=(C1A83>=0)?1:0;

ninexnine_unit ninexnine_unit_2948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10A93)
);

ninexnine_unit ninexnine_unit_2949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11A93)
);

ninexnine_unit ninexnine_unit_2950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12A93)
);

ninexnine_unit ninexnine_unit_2951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13A93)
);

assign C1A93=c10A93+c11A93+c12A93+c13A93;
assign A1A93=(C1A93>=0)?1:0;

ninexnine_unit ninexnine_unit_2952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10AA3)
);

ninexnine_unit ninexnine_unit_2953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11AA3)
);

ninexnine_unit ninexnine_unit_2954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12AA3)
);

ninexnine_unit ninexnine_unit_2955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13AA3)
);

assign C1AA3=c10AA3+c11AA3+c12AA3+c13AA3;
assign A1AA3=(C1AA3>=0)?1:0;

ninexnine_unit ninexnine_unit_2956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10AB3)
);

ninexnine_unit ninexnine_unit_2957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11AB3)
);

ninexnine_unit ninexnine_unit_2958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12AB3)
);

ninexnine_unit ninexnine_unit_2959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13AB3)
);

assign C1AB3=c10AB3+c11AB3+c12AB3+c13AB3;
assign A1AB3=(C1AB3>=0)?1:0;

ninexnine_unit ninexnine_unit_2960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10AC3)
);

ninexnine_unit ninexnine_unit_2961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11AC3)
);

ninexnine_unit ninexnine_unit_2962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12AC3)
);

ninexnine_unit ninexnine_unit_2963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13AC3)
);

assign C1AC3=c10AC3+c11AC3+c12AC3+c13AC3;
assign A1AC3=(C1AC3>=0)?1:0;

ninexnine_unit ninexnine_unit_2964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10AD3)
);

ninexnine_unit ninexnine_unit_2965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11AD3)
);

ninexnine_unit ninexnine_unit_2966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12AD3)
);

ninexnine_unit ninexnine_unit_2967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13AD3)
);

assign C1AD3=c10AD3+c11AD3+c12AD3+c13AD3;
assign A1AD3=(C1AD3>=0)?1:0;

ninexnine_unit ninexnine_unit_2968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B03)
);

ninexnine_unit ninexnine_unit_2969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B03)
);

ninexnine_unit ninexnine_unit_2970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B03)
);

ninexnine_unit ninexnine_unit_2971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B03)
);

assign C1B03=c10B03+c11B03+c12B03+c13B03;
assign A1B03=(C1B03>=0)?1:0;

ninexnine_unit ninexnine_unit_2972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B13)
);

ninexnine_unit ninexnine_unit_2973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B13)
);

ninexnine_unit ninexnine_unit_2974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B13)
);

ninexnine_unit ninexnine_unit_2975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B13)
);

assign C1B13=c10B13+c11B13+c12B13+c13B13;
assign A1B13=(C1B13>=0)?1:0;

ninexnine_unit ninexnine_unit_2976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B23)
);

ninexnine_unit ninexnine_unit_2977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B23)
);

ninexnine_unit ninexnine_unit_2978(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B23)
);

ninexnine_unit ninexnine_unit_2979(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B23)
);

assign C1B23=c10B23+c11B23+c12B23+c13B23;
assign A1B23=(C1B23>=0)?1:0;

ninexnine_unit ninexnine_unit_2980(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B33)
);

ninexnine_unit ninexnine_unit_2981(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B33)
);

ninexnine_unit ninexnine_unit_2982(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B33)
);

ninexnine_unit ninexnine_unit_2983(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B33)
);

assign C1B33=c10B33+c11B33+c12B33+c13B33;
assign A1B33=(C1B33>=0)?1:0;

ninexnine_unit ninexnine_unit_2984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B43)
);

ninexnine_unit ninexnine_unit_2985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B43)
);

ninexnine_unit ninexnine_unit_2986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B43)
);

ninexnine_unit ninexnine_unit_2987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B43)
);

assign C1B43=c10B43+c11B43+c12B43+c13B43;
assign A1B43=(C1B43>=0)?1:0;

ninexnine_unit ninexnine_unit_2988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B53)
);

ninexnine_unit ninexnine_unit_2989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B53)
);

ninexnine_unit ninexnine_unit_2990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B53)
);

ninexnine_unit ninexnine_unit_2991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B53)
);

assign C1B53=c10B53+c11B53+c12B53+c13B53;
assign A1B53=(C1B53>=0)?1:0;

ninexnine_unit ninexnine_unit_2992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B63)
);

ninexnine_unit ninexnine_unit_2993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B63)
);

ninexnine_unit ninexnine_unit_2994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B63)
);

ninexnine_unit ninexnine_unit_2995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B63)
);

assign C1B63=c10B63+c11B63+c12B63+c13B63;
assign A1B63=(C1B63>=0)?1:0;

ninexnine_unit ninexnine_unit_2996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B73)
);

ninexnine_unit ninexnine_unit_2997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B73)
);

ninexnine_unit ninexnine_unit_2998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B73)
);

ninexnine_unit ninexnine_unit_2999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B73)
);

assign C1B73=c10B73+c11B73+c12B73+c13B73;
assign A1B73=(C1B73>=0)?1:0;

ninexnine_unit ninexnine_unit_3000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B83)
);

ninexnine_unit ninexnine_unit_3001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B83)
);

ninexnine_unit ninexnine_unit_3002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B83)
);

ninexnine_unit ninexnine_unit_3003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B83)
);

assign C1B83=c10B83+c11B83+c12B83+c13B83;
assign A1B83=(C1B83>=0)?1:0;

ninexnine_unit ninexnine_unit_3004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10B93)
);

ninexnine_unit ninexnine_unit_3005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11B93)
);

ninexnine_unit ninexnine_unit_3006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12B93)
);

ninexnine_unit ninexnine_unit_3007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13B93)
);

assign C1B93=c10B93+c11B93+c12B93+c13B93;
assign A1B93=(C1B93>=0)?1:0;

ninexnine_unit ninexnine_unit_3008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10BA3)
);

ninexnine_unit ninexnine_unit_3009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11BA3)
);

ninexnine_unit ninexnine_unit_3010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12BA3)
);

ninexnine_unit ninexnine_unit_3011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13BA3)
);

assign C1BA3=c10BA3+c11BA3+c12BA3+c13BA3;
assign A1BA3=(C1BA3>=0)?1:0;

ninexnine_unit ninexnine_unit_3012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10BB3)
);

ninexnine_unit ninexnine_unit_3013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11BB3)
);

ninexnine_unit ninexnine_unit_3014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12BB3)
);

ninexnine_unit ninexnine_unit_3015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13BB3)
);

assign C1BB3=c10BB3+c11BB3+c12BB3+c13BB3;
assign A1BB3=(C1BB3>=0)?1:0;

ninexnine_unit ninexnine_unit_3016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10BC3)
);

ninexnine_unit ninexnine_unit_3017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11BC3)
);

ninexnine_unit ninexnine_unit_3018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12BC3)
);

ninexnine_unit ninexnine_unit_3019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13BC3)
);

assign C1BC3=c10BC3+c11BC3+c12BC3+c13BC3;
assign A1BC3=(C1BC3>=0)?1:0;

ninexnine_unit ninexnine_unit_3020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10BD3)
);

ninexnine_unit ninexnine_unit_3021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11BD3)
);

ninexnine_unit ninexnine_unit_3022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12BD3)
);

ninexnine_unit ninexnine_unit_3023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13BD3)
);

assign C1BD3=c10BD3+c11BD3+c12BD3+c13BD3;
assign A1BD3=(C1BD3>=0)?1:0;

ninexnine_unit ninexnine_unit_3024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C03)
);

ninexnine_unit ninexnine_unit_3025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C03)
);

ninexnine_unit ninexnine_unit_3026(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C03)
);

ninexnine_unit ninexnine_unit_3027(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C03)
);

assign C1C03=c10C03+c11C03+c12C03+c13C03;
assign A1C03=(C1C03>=0)?1:0;

ninexnine_unit ninexnine_unit_3028(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C13)
);

ninexnine_unit ninexnine_unit_3029(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C13)
);

ninexnine_unit ninexnine_unit_3030(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C13)
);

ninexnine_unit ninexnine_unit_3031(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C13)
);

assign C1C13=c10C13+c11C13+c12C13+c13C13;
assign A1C13=(C1C13>=0)?1:0;

ninexnine_unit ninexnine_unit_3032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C23)
);

ninexnine_unit ninexnine_unit_3033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C23)
);

ninexnine_unit ninexnine_unit_3034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C23)
);

ninexnine_unit ninexnine_unit_3035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C23)
);

assign C1C23=c10C23+c11C23+c12C23+c13C23;
assign A1C23=(C1C23>=0)?1:0;

ninexnine_unit ninexnine_unit_3036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C33)
);

ninexnine_unit ninexnine_unit_3037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C33)
);

ninexnine_unit ninexnine_unit_3038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C33)
);

ninexnine_unit ninexnine_unit_3039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C33)
);

assign C1C33=c10C33+c11C33+c12C33+c13C33;
assign A1C33=(C1C33>=0)?1:0;

ninexnine_unit ninexnine_unit_3040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C43)
);

ninexnine_unit ninexnine_unit_3041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C43)
);

ninexnine_unit ninexnine_unit_3042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C43)
);

ninexnine_unit ninexnine_unit_3043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C43)
);

assign C1C43=c10C43+c11C43+c12C43+c13C43;
assign A1C43=(C1C43>=0)?1:0;

ninexnine_unit ninexnine_unit_3044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C53)
);

ninexnine_unit ninexnine_unit_3045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C53)
);

ninexnine_unit ninexnine_unit_3046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C53)
);

ninexnine_unit ninexnine_unit_3047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C53)
);

assign C1C53=c10C53+c11C53+c12C53+c13C53;
assign A1C53=(C1C53>=0)?1:0;

ninexnine_unit ninexnine_unit_3048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C63)
);

ninexnine_unit ninexnine_unit_3049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C63)
);

ninexnine_unit ninexnine_unit_3050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C63)
);

ninexnine_unit ninexnine_unit_3051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C63)
);

assign C1C63=c10C63+c11C63+c12C63+c13C63;
assign A1C63=(C1C63>=0)?1:0;

ninexnine_unit ninexnine_unit_3052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C73)
);

ninexnine_unit ninexnine_unit_3053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C73)
);

ninexnine_unit ninexnine_unit_3054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C73)
);

ninexnine_unit ninexnine_unit_3055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C73)
);

assign C1C73=c10C73+c11C73+c12C73+c13C73;
assign A1C73=(C1C73>=0)?1:0;

ninexnine_unit ninexnine_unit_3056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C83)
);

ninexnine_unit ninexnine_unit_3057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C83)
);

ninexnine_unit ninexnine_unit_3058(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C83)
);

ninexnine_unit ninexnine_unit_3059(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C83)
);

assign C1C83=c10C83+c11C83+c12C83+c13C83;
assign A1C83=(C1C83>=0)?1:0;

ninexnine_unit ninexnine_unit_3060(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10C93)
);

ninexnine_unit ninexnine_unit_3061(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11C93)
);

ninexnine_unit ninexnine_unit_3062(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12C93)
);

ninexnine_unit ninexnine_unit_3063(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13C93)
);

assign C1C93=c10C93+c11C93+c12C93+c13C93;
assign A1C93=(C1C93>=0)?1:0;

ninexnine_unit ninexnine_unit_3064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10CA3)
);

ninexnine_unit ninexnine_unit_3065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11CA3)
);

ninexnine_unit ninexnine_unit_3066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12CA3)
);

ninexnine_unit ninexnine_unit_3067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13CA3)
);

assign C1CA3=c10CA3+c11CA3+c12CA3+c13CA3;
assign A1CA3=(C1CA3>=0)?1:0;

ninexnine_unit ninexnine_unit_3068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10CB3)
);

ninexnine_unit ninexnine_unit_3069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11CB3)
);

ninexnine_unit ninexnine_unit_3070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12CB3)
);

ninexnine_unit ninexnine_unit_3071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13CB3)
);

assign C1CB3=c10CB3+c11CB3+c12CB3+c13CB3;
assign A1CB3=(C1CB3>=0)?1:0;

ninexnine_unit ninexnine_unit_3072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10CC3)
);

ninexnine_unit ninexnine_unit_3073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11CC3)
);

ninexnine_unit ninexnine_unit_3074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12CC3)
);

ninexnine_unit ninexnine_unit_3075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13CC3)
);

assign C1CC3=c10CC3+c11CC3+c12CC3+c13CC3;
assign A1CC3=(C1CC3>=0)?1:0;

ninexnine_unit ninexnine_unit_3076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10CD3)
);

ninexnine_unit ninexnine_unit_3077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11CD3)
);

ninexnine_unit ninexnine_unit_3078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12CD3)
);

ninexnine_unit ninexnine_unit_3079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13CD3)
);

assign C1CD3=c10CD3+c11CD3+c12CD3+c13CD3;
assign A1CD3=(C1CD3>=0)?1:0;

ninexnine_unit ninexnine_unit_3080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D03)
);

ninexnine_unit ninexnine_unit_3081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D03)
);

ninexnine_unit ninexnine_unit_3082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D03)
);

ninexnine_unit ninexnine_unit_3083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D03)
);

assign C1D03=c10D03+c11D03+c12D03+c13D03;
assign A1D03=(C1D03>=0)?1:0;

ninexnine_unit ninexnine_unit_3084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D13)
);

ninexnine_unit ninexnine_unit_3085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D13)
);

ninexnine_unit ninexnine_unit_3086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D13)
);

ninexnine_unit ninexnine_unit_3087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D13)
);

assign C1D13=c10D13+c11D13+c12D13+c13D13;
assign A1D13=(C1D13>=0)?1:0;

ninexnine_unit ninexnine_unit_3088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D23)
);

ninexnine_unit ninexnine_unit_3089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D23)
);

ninexnine_unit ninexnine_unit_3090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D23)
);

ninexnine_unit ninexnine_unit_3091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D23)
);

assign C1D23=c10D23+c11D23+c12D23+c13D23;
assign A1D23=(C1D23>=0)?1:0;

ninexnine_unit ninexnine_unit_3092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D33)
);

ninexnine_unit ninexnine_unit_3093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D33)
);

ninexnine_unit ninexnine_unit_3094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D33)
);

ninexnine_unit ninexnine_unit_3095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D33)
);

assign C1D33=c10D33+c11D33+c12D33+c13D33;
assign A1D33=(C1D33>=0)?1:0;

ninexnine_unit ninexnine_unit_3096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D43)
);

ninexnine_unit ninexnine_unit_3097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D43)
);

ninexnine_unit ninexnine_unit_3098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D43)
);

ninexnine_unit ninexnine_unit_3099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D43)
);

assign C1D43=c10D43+c11D43+c12D43+c13D43;
assign A1D43=(C1D43>=0)?1:0;

ninexnine_unit ninexnine_unit_3100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D53)
);

ninexnine_unit ninexnine_unit_3101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D53)
);

ninexnine_unit ninexnine_unit_3102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D53)
);

ninexnine_unit ninexnine_unit_3103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D53)
);

assign C1D53=c10D53+c11D53+c12D53+c13D53;
assign A1D53=(C1D53>=0)?1:0;

ninexnine_unit ninexnine_unit_3104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D63)
);

ninexnine_unit ninexnine_unit_3105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D63)
);

ninexnine_unit ninexnine_unit_3106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D63)
);

ninexnine_unit ninexnine_unit_3107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D63)
);

assign C1D63=c10D63+c11D63+c12D63+c13D63;
assign A1D63=(C1D63>=0)?1:0;

ninexnine_unit ninexnine_unit_3108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D73)
);

ninexnine_unit ninexnine_unit_3109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D73)
);

ninexnine_unit ninexnine_unit_3110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D73)
);

ninexnine_unit ninexnine_unit_3111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D73)
);

assign C1D73=c10D73+c11D73+c12D73+c13D73;
assign A1D73=(C1D73>=0)?1:0;

ninexnine_unit ninexnine_unit_3112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D83)
);

ninexnine_unit ninexnine_unit_3113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D83)
);

ninexnine_unit ninexnine_unit_3114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D83)
);

ninexnine_unit ninexnine_unit_3115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D83)
);

assign C1D83=c10D83+c11D83+c12D83+c13D83;
assign A1D83=(C1D83>=0)?1:0;

ninexnine_unit ninexnine_unit_3116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10D93)
);

ninexnine_unit ninexnine_unit_3117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11D93)
);

ninexnine_unit ninexnine_unit_3118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12D93)
);

ninexnine_unit ninexnine_unit_3119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13D93)
);

assign C1D93=c10D93+c11D93+c12D93+c13D93;
assign A1D93=(C1D93>=0)?1:0;

ninexnine_unit ninexnine_unit_3120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10DA3)
);

ninexnine_unit ninexnine_unit_3121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11DA3)
);

ninexnine_unit ninexnine_unit_3122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12DA3)
);

ninexnine_unit ninexnine_unit_3123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13DA3)
);

assign C1DA3=c10DA3+c11DA3+c12DA3+c13DA3;
assign A1DA3=(C1DA3>=0)?1:0;

ninexnine_unit ninexnine_unit_3124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10DB3)
);

ninexnine_unit ninexnine_unit_3125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11DB3)
);

ninexnine_unit ninexnine_unit_3126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12DB3)
);

ninexnine_unit ninexnine_unit_3127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13DB3)
);

assign C1DB3=c10DB3+c11DB3+c12DB3+c13DB3;
assign A1DB3=(C1DB3>=0)?1:0;

ninexnine_unit ninexnine_unit_3128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10DC3)
);

ninexnine_unit ninexnine_unit_3129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11DC3)
);

ninexnine_unit ninexnine_unit_3130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12DC3)
);

ninexnine_unit ninexnine_unit_3131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13DC3)
);

assign C1DC3=c10DC3+c11DC3+c12DC3+c13DC3;
assign A1DC3=(C1DC3>=0)?1:0;

ninexnine_unit ninexnine_unit_3132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10DD3)
);

ninexnine_unit ninexnine_unit_3133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11DD3)
);

ninexnine_unit ninexnine_unit_3134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12DD3)
);

ninexnine_unit ninexnine_unit_3135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13DD3)
);

assign C1DD3=c10DD3+c11DD3+c12DD3+c13DD3;
assign A1DD3=(C1DD3>=0)?1:0;

ninexnine_unit ninexnine_unit_3136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10004)
);

ninexnine_unit ninexnine_unit_3137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11004)
);

ninexnine_unit ninexnine_unit_3138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12004)
);

ninexnine_unit ninexnine_unit_3139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13004)
);

assign C1004=c10004+c11004+c12004+c13004;
assign A1004=(C1004>=0)?1:0;

ninexnine_unit ninexnine_unit_3140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10014)
);

ninexnine_unit ninexnine_unit_3141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11014)
);

ninexnine_unit ninexnine_unit_3142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12014)
);

ninexnine_unit ninexnine_unit_3143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13014)
);

assign C1014=c10014+c11014+c12014+c13014;
assign A1014=(C1014>=0)?1:0;

ninexnine_unit ninexnine_unit_3144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10024)
);

ninexnine_unit ninexnine_unit_3145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11024)
);

ninexnine_unit ninexnine_unit_3146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12024)
);

ninexnine_unit ninexnine_unit_3147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13024)
);

assign C1024=c10024+c11024+c12024+c13024;
assign A1024=(C1024>=0)?1:0;

ninexnine_unit ninexnine_unit_3148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10034)
);

ninexnine_unit ninexnine_unit_3149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11034)
);

ninexnine_unit ninexnine_unit_3150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12034)
);

ninexnine_unit ninexnine_unit_3151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13034)
);

assign C1034=c10034+c11034+c12034+c13034;
assign A1034=(C1034>=0)?1:0;

ninexnine_unit ninexnine_unit_3152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10044)
);

ninexnine_unit ninexnine_unit_3153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11044)
);

ninexnine_unit ninexnine_unit_3154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12044)
);

ninexnine_unit ninexnine_unit_3155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13044)
);

assign C1044=c10044+c11044+c12044+c13044;
assign A1044=(C1044>=0)?1:0;

ninexnine_unit ninexnine_unit_3156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10054)
);

ninexnine_unit ninexnine_unit_3157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11054)
);

ninexnine_unit ninexnine_unit_3158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12054)
);

ninexnine_unit ninexnine_unit_3159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13054)
);

assign C1054=c10054+c11054+c12054+c13054;
assign A1054=(C1054>=0)?1:0;

ninexnine_unit ninexnine_unit_3160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10064)
);

ninexnine_unit ninexnine_unit_3161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11064)
);

ninexnine_unit ninexnine_unit_3162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12064)
);

ninexnine_unit ninexnine_unit_3163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13064)
);

assign C1064=c10064+c11064+c12064+c13064;
assign A1064=(C1064>=0)?1:0;

ninexnine_unit ninexnine_unit_3164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10074)
);

ninexnine_unit ninexnine_unit_3165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11074)
);

ninexnine_unit ninexnine_unit_3166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12074)
);

ninexnine_unit ninexnine_unit_3167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13074)
);

assign C1074=c10074+c11074+c12074+c13074;
assign A1074=(C1074>=0)?1:0;

ninexnine_unit ninexnine_unit_3168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10084)
);

ninexnine_unit ninexnine_unit_3169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11084)
);

ninexnine_unit ninexnine_unit_3170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12084)
);

ninexnine_unit ninexnine_unit_3171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13084)
);

assign C1084=c10084+c11084+c12084+c13084;
assign A1084=(C1084>=0)?1:0;

ninexnine_unit ninexnine_unit_3172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10094)
);

ninexnine_unit ninexnine_unit_3173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11094)
);

ninexnine_unit ninexnine_unit_3174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12094)
);

ninexnine_unit ninexnine_unit_3175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13094)
);

assign C1094=c10094+c11094+c12094+c13094;
assign A1094=(C1094>=0)?1:0;

ninexnine_unit ninexnine_unit_3176(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c100A4)
);

ninexnine_unit ninexnine_unit_3177(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c110A4)
);

ninexnine_unit ninexnine_unit_3178(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c120A4)
);

ninexnine_unit ninexnine_unit_3179(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c130A4)
);

assign C10A4=c100A4+c110A4+c120A4+c130A4;
assign A10A4=(C10A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3180(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c100B4)
);

ninexnine_unit ninexnine_unit_3181(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c110B4)
);

ninexnine_unit ninexnine_unit_3182(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c120B4)
);

ninexnine_unit ninexnine_unit_3183(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c130B4)
);

assign C10B4=c100B4+c110B4+c120B4+c130B4;
assign A10B4=(C10B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3184(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c100C4)
);

ninexnine_unit ninexnine_unit_3185(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c110C4)
);

ninexnine_unit ninexnine_unit_3186(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c120C4)
);

ninexnine_unit ninexnine_unit_3187(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c130C4)
);

assign C10C4=c100C4+c110C4+c120C4+c130C4;
assign A10C4=(C10C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3188(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c100D4)
);

ninexnine_unit ninexnine_unit_3189(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c110D4)
);

ninexnine_unit ninexnine_unit_3190(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c120D4)
);

ninexnine_unit ninexnine_unit_3191(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c130D4)
);

assign C10D4=c100D4+c110D4+c120D4+c130D4;
assign A10D4=(C10D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10104)
);

ninexnine_unit ninexnine_unit_3193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11104)
);

ninexnine_unit ninexnine_unit_3194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12104)
);

ninexnine_unit ninexnine_unit_3195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13104)
);

assign C1104=c10104+c11104+c12104+c13104;
assign A1104=(C1104>=0)?1:0;

ninexnine_unit ninexnine_unit_3196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10114)
);

ninexnine_unit ninexnine_unit_3197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11114)
);

ninexnine_unit ninexnine_unit_3198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12114)
);

ninexnine_unit ninexnine_unit_3199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13114)
);

assign C1114=c10114+c11114+c12114+c13114;
assign A1114=(C1114>=0)?1:0;

ninexnine_unit ninexnine_unit_3200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10124)
);

ninexnine_unit ninexnine_unit_3201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11124)
);

ninexnine_unit ninexnine_unit_3202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12124)
);

ninexnine_unit ninexnine_unit_3203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13124)
);

assign C1124=c10124+c11124+c12124+c13124;
assign A1124=(C1124>=0)?1:0;

ninexnine_unit ninexnine_unit_3204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10134)
);

ninexnine_unit ninexnine_unit_3205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11134)
);

ninexnine_unit ninexnine_unit_3206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12134)
);

ninexnine_unit ninexnine_unit_3207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13134)
);

assign C1134=c10134+c11134+c12134+c13134;
assign A1134=(C1134>=0)?1:0;

ninexnine_unit ninexnine_unit_3208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10144)
);

ninexnine_unit ninexnine_unit_3209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11144)
);

ninexnine_unit ninexnine_unit_3210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12144)
);

ninexnine_unit ninexnine_unit_3211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13144)
);

assign C1144=c10144+c11144+c12144+c13144;
assign A1144=(C1144>=0)?1:0;

ninexnine_unit ninexnine_unit_3212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10154)
);

ninexnine_unit ninexnine_unit_3213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11154)
);

ninexnine_unit ninexnine_unit_3214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12154)
);

ninexnine_unit ninexnine_unit_3215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13154)
);

assign C1154=c10154+c11154+c12154+c13154;
assign A1154=(C1154>=0)?1:0;

ninexnine_unit ninexnine_unit_3216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10164)
);

ninexnine_unit ninexnine_unit_3217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11164)
);

ninexnine_unit ninexnine_unit_3218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12164)
);

ninexnine_unit ninexnine_unit_3219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13164)
);

assign C1164=c10164+c11164+c12164+c13164;
assign A1164=(C1164>=0)?1:0;

ninexnine_unit ninexnine_unit_3220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10174)
);

ninexnine_unit ninexnine_unit_3221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11174)
);

ninexnine_unit ninexnine_unit_3222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12174)
);

ninexnine_unit ninexnine_unit_3223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13174)
);

assign C1174=c10174+c11174+c12174+c13174;
assign A1174=(C1174>=0)?1:0;

ninexnine_unit ninexnine_unit_3224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10184)
);

ninexnine_unit ninexnine_unit_3225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11184)
);

ninexnine_unit ninexnine_unit_3226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12184)
);

ninexnine_unit ninexnine_unit_3227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13184)
);

assign C1184=c10184+c11184+c12184+c13184;
assign A1184=(C1184>=0)?1:0;

ninexnine_unit ninexnine_unit_3228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10194)
);

ninexnine_unit ninexnine_unit_3229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11194)
);

ninexnine_unit ninexnine_unit_3230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12194)
);

ninexnine_unit ninexnine_unit_3231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13194)
);

assign C1194=c10194+c11194+c12194+c13194;
assign A1194=(C1194>=0)?1:0;

ninexnine_unit ninexnine_unit_3232(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c101A4)
);

ninexnine_unit ninexnine_unit_3233(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c111A4)
);

ninexnine_unit ninexnine_unit_3234(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c121A4)
);

ninexnine_unit ninexnine_unit_3235(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c131A4)
);

assign C11A4=c101A4+c111A4+c121A4+c131A4;
assign A11A4=(C11A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3236(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c101B4)
);

ninexnine_unit ninexnine_unit_3237(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c111B4)
);

ninexnine_unit ninexnine_unit_3238(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c121B4)
);

ninexnine_unit ninexnine_unit_3239(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c131B4)
);

assign C11B4=c101B4+c111B4+c121B4+c131B4;
assign A11B4=(C11B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3240(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c101C4)
);

ninexnine_unit ninexnine_unit_3241(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c111C4)
);

ninexnine_unit ninexnine_unit_3242(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c121C4)
);

ninexnine_unit ninexnine_unit_3243(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c131C4)
);

assign C11C4=c101C4+c111C4+c121C4+c131C4;
assign A11C4=(C11C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3244(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c101D4)
);

ninexnine_unit ninexnine_unit_3245(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c111D4)
);

ninexnine_unit ninexnine_unit_3246(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c121D4)
);

ninexnine_unit ninexnine_unit_3247(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c131D4)
);

assign C11D4=c101D4+c111D4+c121D4+c131D4;
assign A11D4=(C11D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10204)
);

ninexnine_unit ninexnine_unit_3249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11204)
);

ninexnine_unit ninexnine_unit_3250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12204)
);

ninexnine_unit ninexnine_unit_3251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13204)
);

assign C1204=c10204+c11204+c12204+c13204;
assign A1204=(C1204>=0)?1:0;

ninexnine_unit ninexnine_unit_3252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10214)
);

ninexnine_unit ninexnine_unit_3253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11214)
);

ninexnine_unit ninexnine_unit_3254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12214)
);

ninexnine_unit ninexnine_unit_3255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13214)
);

assign C1214=c10214+c11214+c12214+c13214;
assign A1214=(C1214>=0)?1:0;

ninexnine_unit ninexnine_unit_3256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10224)
);

ninexnine_unit ninexnine_unit_3257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11224)
);

ninexnine_unit ninexnine_unit_3258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12224)
);

ninexnine_unit ninexnine_unit_3259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13224)
);

assign C1224=c10224+c11224+c12224+c13224;
assign A1224=(C1224>=0)?1:0;

ninexnine_unit ninexnine_unit_3260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10234)
);

ninexnine_unit ninexnine_unit_3261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11234)
);

ninexnine_unit ninexnine_unit_3262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12234)
);

ninexnine_unit ninexnine_unit_3263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13234)
);

assign C1234=c10234+c11234+c12234+c13234;
assign A1234=(C1234>=0)?1:0;

ninexnine_unit ninexnine_unit_3264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10244)
);

ninexnine_unit ninexnine_unit_3265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11244)
);

ninexnine_unit ninexnine_unit_3266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12244)
);

ninexnine_unit ninexnine_unit_3267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13244)
);

assign C1244=c10244+c11244+c12244+c13244;
assign A1244=(C1244>=0)?1:0;

ninexnine_unit ninexnine_unit_3268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10254)
);

ninexnine_unit ninexnine_unit_3269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11254)
);

ninexnine_unit ninexnine_unit_3270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12254)
);

ninexnine_unit ninexnine_unit_3271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13254)
);

assign C1254=c10254+c11254+c12254+c13254;
assign A1254=(C1254>=0)?1:0;

ninexnine_unit ninexnine_unit_3272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10264)
);

ninexnine_unit ninexnine_unit_3273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11264)
);

ninexnine_unit ninexnine_unit_3274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12264)
);

ninexnine_unit ninexnine_unit_3275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13264)
);

assign C1264=c10264+c11264+c12264+c13264;
assign A1264=(C1264>=0)?1:0;

ninexnine_unit ninexnine_unit_3276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10274)
);

ninexnine_unit ninexnine_unit_3277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11274)
);

ninexnine_unit ninexnine_unit_3278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12274)
);

ninexnine_unit ninexnine_unit_3279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13274)
);

assign C1274=c10274+c11274+c12274+c13274;
assign A1274=(C1274>=0)?1:0;

ninexnine_unit ninexnine_unit_3280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10284)
);

ninexnine_unit ninexnine_unit_3281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11284)
);

ninexnine_unit ninexnine_unit_3282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12284)
);

ninexnine_unit ninexnine_unit_3283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13284)
);

assign C1284=c10284+c11284+c12284+c13284;
assign A1284=(C1284>=0)?1:0;

ninexnine_unit ninexnine_unit_3284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10294)
);

ninexnine_unit ninexnine_unit_3285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11294)
);

ninexnine_unit ninexnine_unit_3286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12294)
);

ninexnine_unit ninexnine_unit_3287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13294)
);

assign C1294=c10294+c11294+c12294+c13294;
assign A1294=(C1294>=0)?1:0;

ninexnine_unit ninexnine_unit_3288(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c102A4)
);

ninexnine_unit ninexnine_unit_3289(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c112A4)
);

ninexnine_unit ninexnine_unit_3290(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c122A4)
);

ninexnine_unit ninexnine_unit_3291(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c132A4)
);

assign C12A4=c102A4+c112A4+c122A4+c132A4;
assign A12A4=(C12A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3292(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c102B4)
);

ninexnine_unit ninexnine_unit_3293(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c112B4)
);

ninexnine_unit ninexnine_unit_3294(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c122B4)
);

ninexnine_unit ninexnine_unit_3295(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c132B4)
);

assign C12B4=c102B4+c112B4+c122B4+c132B4;
assign A12B4=(C12B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3296(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c102C4)
);

ninexnine_unit ninexnine_unit_3297(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c112C4)
);

ninexnine_unit ninexnine_unit_3298(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c122C4)
);

ninexnine_unit ninexnine_unit_3299(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c132C4)
);

assign C12C4=c102C4+c112C4+c122C4+c132C4;
assign A12C4=(C12C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3300(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c102D4)
);

ninexnine_unit ninexnine_unit_3301(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c112D4)
);

ninexnine_unit ninexnine_unit_3302(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c122D4)
);

ninexnine_unit ninexnine_unit_3303(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c132D4)
);

assign C12D4=c102D4+c112D4+c122D4+c132D4;
assign A12D4=(C12D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10304)
);

ninexnine_unit ninexnine_unit_3305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11304)
);

ninexnine_unit ninexnine_unit_3306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12304)
);

ninexnine_unit ninexnine_unit_3307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13304)
);

assign C1304=c10304+c11304+c12304+c13304;
assign A1304=(C1304>=0)?1:0;

ninexnine_unit ninexnine_unit_3308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10314)
);

ninexnine_unit ninexnine_unit_3309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11314)
);

ninexnine_unit ninexnine_unit_3310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12314)
);

ninexnine_unit ninexnine_unit_3311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13314)
);

assign C1314=c10314+c11314+c12314+c13314;
assign A1314=(C1314>=0)?1:0;

ninexnine_unit ninexnine_unit_3312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10324)
);

ninexnine_unit ninexnine_unit_3313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11324)
);

ninexnine_unit ninexnine_unit_3314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12324)
);

ninexnine_unit ninexnine_unit_3315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13324)
);

assign C1324=c10324+c11324+c12324+c13324;
assign A1324=(C1324>=0)?1:0;

ninexnine_unit ninexnine_unit_3316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10334)
);

ninexnine_unit ninexnine_unit_3317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11334)
);

ninexnine_unit ninexnine_unit_3318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12334)
);

ninexnine_unit ninexnine_unit_3319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13334)
);

assign C1334=c10334+c11334+c12334+c13334;
assign A1334=(C1334>=0)?1:0;

ninexnine_unit ninexnine_unit_3320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10344)
);

ninexnine_unit ninexnine_unit_3321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11344)
);

ninexnine_unit ninexnine_unit_3322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12344)
);

ninexnine_unit ninexnine_unit_3323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13344)
);

assign C1344=c10344+c11344+c12344+c13344;
assign A1344=(C1344>=0)?1:0;

ninexnine_unit ninexnine_unit_3324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10354)
);

ninexnine_unit ninexnine_unit_3325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11354)
);

ninexnine_unit ninexnine_unit_3326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12354)
);

ninexnine_unit ninexnine_unit_3327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13354)
);

assign C1354=c10354+c11354+c12354+c13354;
assign A1354=(C1354>=0)?1:0;

ninexnine_unit ninexnine_unit_3328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10364)
);

ninexnine_unit ninexnine_unit_3329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11364)
);

ninexnine_unit ninexnine_unit_3330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12364)
);

ninexnine_unit ninexnine_unit_3331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13364)
);

assign C1364=c10364+c11364+c12364+c13364;
assign A1364=(C1364>=0)?1:0;

ninexnine_unit ninexnine_unit_3332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10374)
);

ninexnine_unit ninexnine_unit_3333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11374)
);

ninexnine_unit ninexnine_unit_3334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12374)
);

ninexnine_unit ninexnine_unit_3335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13374)
);

assign C1374=c10374+c11374+c12374+c13374;
assign A1374=(C1374>=0)?1:0;

ninexnine_unit ninexnine_unit_3336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10384)
);

ninexnine_unit ninexnine_unit_3337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11384)
);

ninexnine_unit ninexnine_unit_3338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12384)
);

ninexnine_unit ninexnine_unit_3339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13384)
);

assign C1384=c10384+c11384+c12384+c13384;
assign A1384=(C1384>=0)?1:0;

ninexnine_unit ninexnine_unit_3340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10394)
);

ninexnine_unit ninexnine_unit_3341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11394)
);

ninexnine_unit ninexnine_unit_3342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12394)
);

ninexnine_unit ninexnine_unit_3343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13394)
);

assign C1394=c10394+c11394+c12394+c13394;
assign A1394=(C1394>=0)?1:0;

ninexnine_unit ninexnine_unit_3344(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c103A4)
);

ninexnine_unit ninexnine_unit_3345(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c113A4)
);

ninexnine_unit ninexnine_unit_3346(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c123A4)
);

ninexnine_unit ninexnine_unit_3347(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c133A4)
);

assign C13A4=c103A4+c113A4+c123A4+c133A4;
assign A13A4=(C13A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3348(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c103B4)
);

ninexnine_unit ninexnine_unit_3349(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c113B4)
);

ninexnine_unit ninexnine_unit_3350(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c123B4)
);

ninexnine_unit ninexnine_unit_3351(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c133B4)
);

assign C13B4=c103B4+c113B4+c123B4+c133B4;
assign A13B4=(C13B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3352(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c103C4)
);

ninexnine_unit ninexnine_unit_3353(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c113C4)
);

ninexnine_unit ninexnine_unit_3354(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c123C4)
);

ninexnine_unit ninexnine_unit_3355(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c133C4)
);

assign C13C4=c103C4+c113C4+c123C4+c133C4;
assign A13C4=(C13C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3356(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c103D4)
);

ninexnine_unit ninexnine_unit_3357(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c113D4)
);

ninexnine_unit ninexnine_unit_3358(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c123D4)
);

ninexnine_unit ninexnine_unit_3359(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c133D4)
);

assign C13D4=c103D4+c113D4+c123D4+c133D4;
assign A13D4=(C13D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10404)
);

ninexnine_unit ninexnine_unit_3361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11404)
);

ninexnine_unit ninexnine_unit_3362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12404)
);

ninexnine_unit ninexnine_unit_3363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13404)
);

assign C1404=c10404+c11404+c12404+c13404;
assign A1404=(C1404>=0)?1:0;

ninexnine_unit ninexnine_unit_3364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10414)
);

ninexnine_unit ninexnine_unit_3365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11414)
);

ninexnine_unit ninexnine_unit_3366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12414)
);

ninexnine_unit ninexnine_unit_3367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13414)
);

assign C1414=c10414+c11414+c12414+c13414;
assign A1414=(C1414>=0)?1:0;

ninexnine_unit ninexnine_unit_3368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10424)
);

ninexnine_unit ninexnine_unit_3369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11424)
);

ninexnine_unit ninexnine_unit_3370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12424)
);

ninexnine_unit ninexnine_unit_3371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13424)
);

assign C1424=c10424+c11424+c12424+c13424;
assign A1424=(C1424>=0)?1:0;

ninexnine_unit ninexnine_unit_3372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10434)
);

ninexnine_unit ninexnine_unit_3373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11434)
);

ninexnine_unit ninexnine_unit_3374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12434)
);

ninexnine_unit ninexnine_unit_3375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13434)
);

assign C1434=c10434+c11434+c12434+c13434;
assign A1434=(C1434>=0)?1:0;

ninexnine_unit ninexnine_unit_3376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10444)
);

ninexnine_unit ninexnine_unit_3377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11444)
);

ninexnine_unit ninexnine_unit_3378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12444)
);

ninexnine_unit ninexnine_unit_3379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13444)
);

assign C1444=c10444+c11444+c12444+c13444;
assign A1444=(C1444>=0)?1:0;

ninexnine_unit ninexnine_unit_3380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10454)
);

ninexnine_unit ninexnine_unit_3381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11454)
);

ninexnine_unit ninexnine_unit_3382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12454)
);

ninexnine_unit ninexnine_unit_3383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13454)
);

assign C1454=c10454+c11454+c12454+c13454;
assign A1454=(C1454>=0)?1:0;

ninexnine_unit ninexnine_unit_3384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10464)
);

ninexnine_unit ninexnine_unit_3385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11464)
);

ninexnine_unit ninexnine_unit_3386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12464)
);

ninexnine_unit ninexnine_unit_3387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13464)
);

assign C1464=c10464+c11464+c12464+c13464;
assign A1464=(C1464>=0)?1:0;

ninexnine_unit ninexnine_unit_3388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10474)
);

ninexnine_unit ninexnine_unit_3389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11474)
);

ninexnine_unit ninexnine_unit_3390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12474)
);

ninexnine_unit ninexnine_unit_3391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13474)
);

assign C1474=c10474+c11474+c12474+c13474;
assign A1474=(C1474>=0)?1:0;

ninexnine_unit ninexnine_unit_3392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10484)
);

ninexnine_unit ninexnine_unit_3393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11484)
);

ninexnine_unit ninexnine_unit_3394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12484)
);

ninexnine_unit ninexnine_unit_3395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13484)
);

assign C1484=c10484+c11484+c12484+c13484;
assign A1484=(C1484>=0)?1:0;

ninexnine_unit ninexnine_unit_3396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10494)
);

ninexnine_unit ninexnine_unit_3397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11494)
);

ninexnine_unit ninexnine_unit_3398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12494)
);

ninexnine_unit ninexnine_unit_3399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13494)
);

assign C1494=c10494+c11494+c12494+c13494;
assign A1494=(C1494>=0)?1:0;

ninexnine_unit ninexnine_unit_3400(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c104A4)
);

ninexnine_unit ninexnine_unit_3401(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c114A4)
);

ninexnine_unit ninexnine_unit_3402(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c124A4)
);

ninexnine_unit ninexnine_unit_3403(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c134A4)
);

assign C14A4=c104A4+c114A4+c124A4+c134A4;
assign A14A4=(C14A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3404(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c104B4)
);

ninexnine_unit ninexnine_unit_3405(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c114B4)
);

ninexnine_unit ninexnine_unit_3406(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c124B4)
);

ninexnine_unit ninexnine_unit_3407(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c134B4)
);

assign C14B4=c104B4+c114B4+c124B4+c134B4;
assign A14B4=(C14B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3408(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c104C4)
);

ninexnine_unit ninexnine_unit_3409(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c114C4)
);

ninexnine_unit ninexnine_unit_3410(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c124C4)
);

ninexnine_unit ninexnine_unit_3411(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c134C4)
);

assign C14C4=c104C4+c114C4+c124C4+c134C4;
assign A14C4=(C14C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3412(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c104D4)
);

ninexnine_unit ninexnine_unit_3413(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c114D4)
);

ninexnine_unit ninexnine_unit_3414(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c124D4)
);

ninexnine_unit ninexnine_unit_3415(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c134D4)
);

assign C14D4=c104D4+c114D4+c124D4+c134D4;
assign A14D4=(C14D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10504)
);

ninexnine_unit ninexnine_unit_3417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11504)
);

ninexnine_unit ninexnine_unit_3418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12504)
);

ninexnine_unit ninexnine_unit_3419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13504)
);

assign C1504=c10504+c11504+c12504+c13504;
assign A1504=(C1504>=0)?1:0;

ninexnine_unit ninexnine_unit_3420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10514)
);

ninexnine_unit ninexnine_unit_3421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11514)
);

ninexnine_unit ninexnine_unit_3422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12514)
);

ninexnine_unit ninexnine_unit_3423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13514)
);

assign C1514=c10514+c11514+c12514+c13514;
assign A1514=(C1514>=0)?1:0;

ninexnine_unit ninexnine_unit_3424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10524)
);

ninexnine_unit ninexnine_unit_3425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11524)
);

ninexnine_unit ninexnine_unit_3426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12524)
);

ninexnine_unit ninexnine_unit_3427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13524)
);

assign C1524=c10524+c11524+c12524+c13524;
assign A1524=(C1524>=0)?1:0;

ninexnine_unit ninexnine_unit_3428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10534)
);

ninexnine_unit ninexnine_unit_3429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11534)
);

ninexnine_unit ninexnine_unit_3430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12534)
);

ninexnine_unit ninexnine_unit_3431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13534)
);

assign C1534=c10534+c11534+c12534+c13534;
assign A1534=(C1534>=0)?1:0;

ninexnine_unit ninexnine_unit_3432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10544)
);

ninexnine_unit ninexnine_unit_3433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11544)
);

ninexnine_unit ninexnine_unit_3434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12544)
);

ninexnine_unit ninexnine_unit_3435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13544)
);

assign C1544=c10544+c11544+c12544+c13544;
assign A1544=(C1544>=0)?1:0;

ninexnine_unit ninexnine_unit_3436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10554)
);

ninexnine_unit ninexnine_unit_3437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11554)
);

ninexnine_unit ninexnine_unit_3438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12554)
);

ninexnine_unit ninexnine_unit_3439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13554)
);

assign C1554=c10554+c11554+c12554+c13554;
assign A1554=(C1554>=0)?1:0;

ninexnine_unit ninexnine_unit_3440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10564)
);

ninexnine_unit ninexnine_unit_3441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11564)
);

ninexnine_unit ninexnine_unit_3442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12564)
);

ninexnine_unit ninexnine_unit_3443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13564)
);

assign C1564=c10564+c11564+c12564+c13564;
assign A1564=(C1564>=0)?1:0;

ninexnine_unit ninexnine_unit_3444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10574)
);

ninexnine_unit ninexnine_unit_3445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11574)
);

ninexnine_unit ninexnine_unit_3446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12574)
);

ninexnine_unit ninexnine_unit_3447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13574)
);

assign C1574=c10574+c11574+c12574+c13574;
assign A1574=(C1574>=0)?1:0;

ninexnine_unit ninexnine_unit_3448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10584)
);

ninexnine_unit ninexnine_unit_3449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11584)
);

ninexnine_unit ninexnine_unit_3450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12584)
);

ninexnine_unit ninexnine_unit_3451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13584)
);

assign C1584=c10584+c11584+c12584+c13584;
assign A1584=(C1584>=0)?1:0;

ninexnine_unit ninexnine_unit_3452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10594)
);

ninexnine_unit ninexnine_unit_3453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11594)
);

ninexnine_unit ninexnine_unit_3454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12594)
);

ninexnine_unit ninexnine_unit_3455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13594)
);

assign C1594=c10594+c11594+c12594+c13594;
assign A1594=(C1594>=0)?1:0;

ninexnine_unit ninexnine_unit_3456(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c105A4)
);

ninexnine_unit ninexnine_unit_3457(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c115A4)
);

ninexnine_unit ninexnine_unit_3458(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c125A4)
);

ninexnine_unit ninexnine_unit_3459(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c135A4)
);

assign C15A4=c105A4+c115A4+c125A4+c135A4;
assign A15A4=(C15A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3460(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c105B4)
);

ninexnine_unit ninexnine_unit_3461(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c115B4)
);

ninexnine_unit ninexnine_unit_3462(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c125B4)
);

ninexnine_unit ninexnine_unit_3463(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c135B4)
);

assign C15B4=c105B4+c115B4+c125B4+c135B4;
assign A15B4=(C15B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3464(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c105C4)
);

ninexnine_unit ninexnine_unit_3465(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c115C4)
);

ninexnine_unit ninexnine_unit_3466(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c125C4)
);

ninexnine_unit ninexnine_unit_3467(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c135C4)
);

assign C15C4=c105C4+c115C4+c125C4+c135C4;
assign A15C4=(C15C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3468(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c105D4)
);

ninexnine_unit ninexnine_unit_3469(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c115D4)
);

ninexnine_unit ninexnine_unit_3470(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c125D4)
);

ninexnine_unit ninexnine_unit_3471(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c135D4)
);

assign C15D4=c105D4+c115D4+c125D4+c135D4;
assign A15D4=(C15D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10604)
);

ninexnine_unit ninexnine_unit_3473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11604)
);

ninexnine_unit ninexnine_unit_3474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12604)
);

ninexnine_unit ninexnine_unit_3475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13604)
);

assign C1604=c10604+c11604+c12604+c13604;
assign A1604=(C1604>=0)?1:0;

ninexnine_unit ninexnine_unit_3476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10614)
);

ninexnine_unit ninexnine_unit_3477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11614)
);

ninexnine_unit ninexnine_unit_3478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12614)
);

ninexnine_unit ninexnine_unit_3479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13614)
);

assign C1614=c10614+c11614+c12614+c13614;
assign A1614=(C1614>=0)?1:0;

ninexnine_unit ninexnine_unit_3480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10624)
);

ninexnine_unit ninexnine_unit_3481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11624)
);

ninexnine_unit ninexnine_unit_3482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12624)
);

ninexnine_unit ninexnine_unit_3483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13624)
);

assign C1624=c10624+c11624+c12624+c13624;
assign A1624=(C1624>=0)?1:0;

ninexnine_unit ninexnine_unit_3484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10634)
);

ninexnine_unit ninexnine_unit_3485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11634)
);

ninexnine_unit ninexnine_unit_3486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12634)
);

ninexnine_unit ninexnine_unit_3487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13634)
);

assign C1634=c10634+c11634+c12634+c13634;
assign A1634=(C1634>=0)?1:0;

ninexnine_unit ninexnine_unit_3488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10644)
);

ninexnine_unit ninexnine_unit_3489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11644)
);

ninexnine_unit ninexnine_unit_3490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12644)
);

ninexnine_unit ninexnine_unit_3491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13644)
);

assign C1644=c10644+c11644+c12644+c13644;
assign A1644=(C1644>=0)?1:0;

ninexnine_unit ninexnine_unit_3492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10654)
);

ninexnine_unit ninexnine_unit_3493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11654)
);

ninexnine_unit ninexnine_unit_3494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12654)
);

ninexnine_unit ninexnine_unit_3495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13654)
);

assign C1654=c10654+c11654+c12654+c13654;
assign A1654=(C1654>=0)?1:0;

ninexnine_unit ninexnine_unit_3496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10664)
);

ninexnine_unit ninexnine_unit_3497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11664)
);

ninexnine_unit ninexnine_unit_3498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12664)
);

ninexnine_unit ninexnine_unit_3499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13664)
);

assign C1664=c10664+c11664+c12664+c13664;
assign A1664=(C1664>=0)?1:0;

ninexnine_unit ninexnine_unit_3500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10674)
);

ninexnine_unit ninexnine_unit_3501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11674)
);

ninexnine_unit ninexnine_unit_3502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12674)
);

ninexnine_unit ninexnine_unit_3503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13674)
);

assign C1674=c10674+c11674+c12674+c13674;
assign A1674=(C1674>=0)?1:0;

ninexnine_unit ninexnine_unit_3504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10684)
);

ninexnine_unit ninexnine_unit_3505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11684)
);

ninexnine_unit ninexnine_unit_3506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12684)
);

ninexnine_unit ninexnine_unit_3507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13684)
);

assign C1684=c10684+c11684+c12684+c13684;
assign A1684=(C1684>=0)?1:0;

ninexnine_unit ninexnine_unit_3508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10694)
);

ninexnine_unit ninexnine_unit_3509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11694)
);

ninexnine_unit ninexnine_unit_3510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12694)
);

ninexnine_unit ninexnine_unit_3511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13694)
);

assign C1694=c10694+c11694+c12694+c13694;
assign A1694=(C1694>=0)?1:0;

ninexnine_unit ninexnine_unit_3512(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c106A4)
);

ninexnine_unit ninexnine_unit_3513(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c116A4)
);

ninexnine_unit ninexnine_unit_3514(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c126A4)
);

ninexnine_unit ninexnine_unit_3515(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c136A4)
);

assign C16A4=c106A4+c116A4+c126A4+c136A4;
assign A16A4=(C16A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3516(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c106B4)
);

ninexnine_unit ninexnine_unit_3517(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c116B4)
);

ninexnine_unit ninexnine_unit_3518(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c126B4)
);

ninexnine_unit ninexnine_unit_3519(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c136B4)
);

assign C16B4=c106B4+c116B4+c126B4+c136B4;
assign A16B4=(C16B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3520(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c106C4)
);

ninexnine_unit ninexnine_unit_3521(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c116C4)
);

ninexnine_unit ninexnine_unit_3522(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c126C4)
);

ninexnine_unit ninexnine_unit_3523(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c136C4)
);

assign C16C4=c106C4+c116C4+c126C4+c136C4;
assign A16C4=(C16C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3524(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c106D4)
);

ninexnine_unit ninexnine_unit_3525(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c116D4)
);

ninexnine_unit ninexnine_unit_3526(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c126D4)
);

ninexnine_unit ninexnine_unit_3527(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c136D4)
);

assign C16D4=c106D4+c116D4+c126D4+c136D4;
assign A16D4=(C16D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10704)
);

ninexnine_unit ninexnine_unit_3529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11704)
);

ninexnine_unit ninexnine_unit_3530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12704)
);

ninexnine_unit ninexnine_unit_3531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13704)
);

assign C1704=c10704+c11704+c12704+c13704;
assign A1704=(C1704>=0)?1:0;

ninexnine_unit ninexnine_unit_3532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10714)
);

ninexnine_unit ninexnine_unit_3533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11714)
);

ninexnine_unit ninexnine_unit_3534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12714)
);

ninexnine_unit ninexnine_unit_3535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13714)
);

assign C1714=c10714+c11714+c12714+c13714;
assign A1714=(C1714>=0)?1:0;

ninexnine_unit ninexnine_unit_3536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10724)
);

ninexnine_unit ninexnine_unit_3537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11724)
);

ninexnine_unit ninexnine_unit_3538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12724)
);

ninexnine_unit ninexnine_unit_3539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13724)
);

assign C1724=c10724+c11724+c12724+c13724;
assign A1724=(C1724>=0)?1:0;

ninexnine_unit ninexnine_unit_3540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10734)
);

ninexnine_unit ninexnine_unit_3541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11734)
);

ninexnine_unit ninexnine_unit_3542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12734)
);

ninexnine_unit ninexnine_unit_3543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13734)
);

assign C1734=c10734+c11734+c12734+c13734;
assign A1734=(C1734>=0)?1:0;

ninexnine_unit ninexnine_unit_3544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10744)
);

ninexnine_unit ninexnine_unit_3545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11744)
);

ninexnine_unit ninexnine_unit_3546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12744)
);

ninexnine_unit ninexnine_unit_3547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13744)
);

assign C1744=c10744+c11744+c12744+c13744;
assign A1744=(C1744>=0)?1:0;

ninexnine_unit ninexnine_unit_3548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10754)
);

ninexnine_unit ninexnine_unit_3549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11754)
);

ninexnine_unit ninexnine_unit_3550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12754)
);

ninexnine_unit ninexnine_unit_3551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13754)
);

assign C1754=c10754+c11754+c12754+c13754;
assign A1754=(C1754>=0)?1:0;

ninexnine_unit ninexnine_unit_3552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10764)
);

ninexnine_unit ninexnine_unit_3553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11764)
);

ninexnine_unit ninexnine_unit_3554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12764)
);

ninexnine_unit ninexnine_unit_3555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13764)
);

assign C1764=c10764+c11764+c12764+c13764;
assign A1764=(C1764>=0)?1:0;

ninexnine_unit ninexnine_unit_3556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10774)
);

ninexnine_unit ninexnine_unit_3557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11774)
);

ninexnine_unit ninexnine_unit_3558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12774)
);

ninexnine_unit ninexnine_unit_3559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13774)
);

assign C1774=c10774+c11774+c12774+c13774;
assign A1774=(C1774>=0)?1:0;

ninexnine_unit ninexnine_unit_3560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10784)
);

ninexnine_unit ninexnine_unit_3561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11784)
);

ninexnine_unit ninexnine_unit_3562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12784)
);

ninexnine_unit ninexnine_unit_3563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13784)
);

assign C1784=c10784+c11784+c12784+c13784;
assign A1784=(C1784>=0)?1:0;

ninexnine_unit ninexnine_unit_3564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10794)
);

ninexnine_unit ninexnine_unit_3565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11794)
);

ninexnine_unit ninexnine_unit_3566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12794)
);

ninexnine_unit ninexnine_unit_3567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13794)
);

assign C1794=c10794+c11794+c12794+c13794;
assign A1794=(C1794>=0)?1:0;

ninexnine_unit ninexnine_unit_3568(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c107A4)
);

ninexnine_unit ninexnine_unit_3569(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c117A4)
);

ninexnine_unit ninexnine_unit_3570(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c127A4)
);

ninexnine_unit ninexnine_unit_3571(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c137A4)
);

assign C17A4=c107A4+c117A4+c127A4+c137A4;
assign A17A4=(C17A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3572(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c107B4)
);

ninexnine_unit ninexnine_unit_3573(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c117B4)
);

ninexnine_unit ninexnine_unit_3574(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c127B4)
);

ninexnine_unit ninexnine_unit_3575(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c137B4)
);

assign C17B4=c107B4+c117B4+c127B4+c137B4;
assign A17B4=(C17B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3576(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c107C4)
);

ninexnine_unit ninexnine_unit_3577(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c117C4)
);

ninexnine_unit ninexnine_unit_3578(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c127C4)
);

ninexnine_unit ninexnine_unit_3579(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c137C4)
);

assign C17C4=c107C4+c117C4+c127C4+c137C4;
assign A17C4=(C17C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3580(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c107D4)
);

ninexnine_unit ninexnine_unit_3581(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c117D4)
);

ninexnine_unit ninexnine_unit_3582(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c127D4)
);

ninexnine_unit ninexnine_unit_3583(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c137D4)
);

assign C17D4=c107D4+c117D4+c127D4+c137D4;
assign A17D4=(C17D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10804)
);

ninexnine_unit ninexnine_unit_3585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11804)
);

ninexnine_unit ninexnine_unit_3586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12804)
);

ninexnine_unit ninexnine_unit_3587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13804)
);

assign C1804=c10804+c11804+c12804+c13804;
assign A1804=(C1804>=0)?1:0;

ninexnine_unit ninexnine_unit_3588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10814)
);

ninexnine_unit ninexnine_unit_3589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11814)
);

ninexnine_unit ninexnine_unit_3590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12814)
);

ninexnine_unit ninexnine_unit_3591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13814)
);

assign C1814=c10814+c11814+c12814+c13814;
assign A1814=(C1814>=0)?1:0;

ninexnine_unit ninexnine_unit_3592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10824)
);

ninexnine_unit ninexnine_unit_3593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11824)
);

ninexnine_unit ninexnine_unit_3594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12824)
);

ninexnine_unit ninexnine_unit_3595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13824)
);

assign C1824=c10824+c11824+c12824+c13824;
assign A1824=(C1824>=0)?1:0;

ninexnine_unit ninexnine_unit_3596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10834)
);

ninexnine_unit ninexnine_unit_3597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11834)
);

ninexnine_unit ninexnine_unit_3598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12834)
);

ninexnine_unit ninexnine_unit_3599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13834)
);

assign C1834=c10834+c11834+c12834+c13834;
assign A1834=(C1834>=0)?1:0;

ninexnine_unit ninexnine_unit_3600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10844)
);

ninexnine_unit ninexnine_unit_3601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11844)
);

ninexnine_unit ninexnine_unit_3602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12844)
);

ninexnine_unit ninexnine_unit_3603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13844)
);

assign C1844=c10844+c11844+c12844+c13844;
assign A1844=(C1844>=0)?1:0;

ninexnine_unit ninexnine_unit_3604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10854)
);

ninexnine_unit ninexnine_unit_3605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11854)
);

ninexnine_unit ninexnine_unit_3606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12854)
);

ninexnine_unit ninexnine_unit_3607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13854)
);

assign C1854=c10854+c11854+c12854+c13854;
assign A1854=(C1854>=0)?1:0;

ninexnine_unit ninexnine_unit_3608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10864)
);

ninexnine_unit ninexnine_unit_3609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11864)
);

ninexnine_unit ninexnine_unit_3610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12864)
);

ninexnine_unit ninexnine_unit_3611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13864)
);

assign C1864=c10864+c11864+c12864+c13864;
assign A1864=(C1864>=0)?1:0;

ninexnine_unit ninexnine_unit_3612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10874)
);

ninexnine_unit ninexnine_unit_3613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11874)
);

ninexnine_unit ninexnine_unit_3614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12874)
);

ninexnine_unit ninexnine_unit_3615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13874)
);

assign C1874=c10874+c11874+c12874+c13874;
assign A1874=(C1874>=0)?1:0;

ninexnine_unit ninexnine_unit_3616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10884)
);

ninexnine_unit ninexnine_unit_3617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11884)
);

ninexnine_unit ninexnine_unit_3618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12884)
);

ninexnine_unit ninexnine_unit_3619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13884)
);

assign C1884=c10884+c11884+c12884+c13884;
assign A1884=(C1884>=0)?1:0;

ninexnine_unit ninexnine_unit_3620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10894)
);

ninexnine_unit ninexnine_unit_3621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11894)
);

ninexnine_unit ninexnine_unit_3622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12894)
);

ninexnine_unit ninexnine_unit_3623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13894)
);

assign C1894=c10894+c11894+c12894+c13894;
assign A1894=(C1894>=0)?1:0;

ninexnine_unit ninexnine_unit_3624(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c108A4)
);

ninexnine_unit ninexnine_unit_3625(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c118A4)
);

ninexnine_unit ninexnine_unit_3626(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c128A4)
);

ninexnine_unit ninexnine_unit_3627(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c138A4)
);

assign C18A4=c108A4+c118A4+c128A4+c138A4;
assign A18A4=(C18A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3628(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c108B4)
);

ninexnine_unit ninexnine_unit_3629(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c118B4)
);

ninexnine_unit ninexnine_unit_3630(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c128B4)
);

ninexnine_unit ninexnine_unit_3631(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c138B4)
);

assign C18B4=c108B4+c118B4+c128B4+c138B4;
assign A18B4=(C18B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3632(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c108C4)
);

ninexnine_unit ninexnine_unit_3633(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c118C4)
);

ninexnine_unit ninexnine_unit_3634(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c128C4)
);

ninexnine_unit ninexnine_unit_3635(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c138C4)
);

assign C18C4=c108C4+c118C4+c128C4+c138C4;
assign A18C4=(C18C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3636(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c108D4)
);

ninexnine_unit ninexnine_unit_3637(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c118D4)
);

ninexnine_unit ninexnine_unit_3638(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c128D4)
);

ninexnine_unit ninexnine_unit_3639(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c138D4)
);

assign C18D4=c108D4+c118D4+c128D4+c138D4;
assign A18D4=(C18D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10904)
);

ninexnine_unit ninexnine_unit_3641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11904)
);

ninexnine_unit ninexnine_unit_3642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12904)
);

ninexnine_unit ninexnine_unit_3643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13904)
);

assign C1904=c10904+c11904+c12904+c13904;
assign A1904=(C1904>=0)?1:0;

ninexnine_unit ninexnine_unit_3644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10914)
);

ninexnine_unit ninexnine_unit_3645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11914)
);

ninexnine_unit ninexnine_unit_3646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12914)
);

ninexnine_unit ninexnine_unit_3647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13914)
);

assign C1914=c10914+c11914+c12914+c13914;
assign A1914=(C1914>=0)?1:0;

ninexnine_unit ninexnine_unit_3648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10924)
);

ninexnine_unit ninexnine_unit_3649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11924)
);

ninexnine_unit ninexnine_unit_3650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12924)
);

ninexnine_unit ninexnine_unit_3651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13924)
);

assign C1924=c10924+c11924+c12924+c13924;
assign A1924=(C1924>=0)?1:0;

ninexnine_unit ninexnine_unit_3652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10934)
);

ninexnine_unit ninexnine_unit_3653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11934)
);

ninexnine_unit ninexnine_unit_3654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12934)
);

ninexnine_unit ninexnine_unit_3655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13934)
);

assign C1934=c10934+c11934+c12934+c13934;
assign A1934=(C1934>=0)?1:0;

ninexnine_unit ninexnine_unit_3656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10944)
);

ninexnine_unit ninexnine_unit_3657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11944)
);

ninexnine_unit ninexnine_unit_3658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12944)
);

ninexnine_unit ninexnine_unit_3659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13944)
);

assign C1944=c10944+c11944+c12944+c13944;
assign A1944=(C1944>=0)?1:0;

ninexnine_unit ninexnine_unit_3660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10954)
);

ninexnine_unit ninexnine_unit_3661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11954)
);

ninexnine_unit ninexnine_unit_3662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12954)
);

ninexnine_unit ninexnine_unit_3663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13954)
);

assign C1954=c10954+c11954+c12954+c13954;
assign A1954=(C1954>=0)?1:0;

ninexnine_unit ninexnine_unit_3664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10964)
);

ninexnine_unit ninexnine_unit_3665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11964)
);

ninexnine_unit ninexnine_unit_3666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12964)
);

ninexnine_unit ninexnine_unit_3667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13964)
);

assign C1964=c10964+c11964+c12964+c13964;
assign A1964=(C1964>=0)?1:0;

ninexnine_unit ninexnine_unit_3668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10974)
);

ninexnine_unit ninexnine_unit_3669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11974)
);

ninexnine_unit ninexnine_unit_3670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12974)
);

ninexnine_unit ninexnine_unit_3671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13974)
);

assign C1974=c10974+c11974+c12974+c13974;
assign A1974=(C1974>=0)?1:0;

ninexnine_unit ninexnine_unit_3672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10984)
);

ninexnine_unit ninexnine_unit_3673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11984)
);

ninexnine_unit ninexnine_unit_3674(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12984)
);

ninexnine_unit ninexnine_unit_3675(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13984)
);

assign C1984=c10984+c11984+c12984+c13984;
assign A1984=(C1984>=0)?1:0;

ninexnine_unit ninexnine_unit_3676(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10994)
);

ninexnine_unit ninexnine_unit_3677(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11994)
);

ninexnine_unit ninexnine_unit_3678(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12994)
);

ninexnine_unit ninexnine_unit_3679(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13994)
);

assign C1994=c10994+c11994+c12994+c13994;
assign A1994=(C1994>=0)?1:0;

ninexnine_unit ninexnine_unit_3680(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c109A4)
);

ninexnine_unit ninexnine_unit_3681(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c119A4)
);

ninexnine_unit ninexnine_unit_3682(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c129A4)
);

ninexnine_unit ninexnine_unit_3683(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c139A4)
);

assign C19A4=c109A4+c119A4+c129A4+c139A4;
assign A19A4=(C19A4>=0)?1:0;

ninexnine_unit ninexnine_unit_3684(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c109B4)
);

ninexnine_unit ninexnine_unit_3685(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c119B4)
);

ninexnine_unit ninexnine_unit_3686(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c129B4)
);

ninexnine_unit ninexnine_unit_3687(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c139B4)
);

assign C19B4=c109B4+c119B4+c129B4+c139B4;
assign A19B4=(C19B4>=0)?1:0;

ninexnine_unit ninexnine_unit_3688(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c109C4)
);

ninexnine_unit ninexnine_unit_3689(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c119C4)
);

ninexnine_unit ninexnine_unit_3690(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c129C4)
);

ninexnine_unit ninexnine_unit_3691(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c139C4)
);

assign C19C4=c109C4+c119C4+c129C4+c139C4;
assign A19C4=(C19C4>=0)?1:0;

ninexnine_unit ninexnine_unit_3692(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c109D4)
);

ninexnine_unit ninexnine_unit_3693(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c119D4)
);

ninexnine_unit ninexnine_unit_3694(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c129D4)
);

ninexnine_unit ninexnine_unit_3695(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c139D4)
);

assign C19D4=c109D4+c119D4+c129D4+c139D4;
assign A19D4=(C19D4>=0)?1:0;

ninexnine_unit ninexnine_unit_3696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A04)
);

ninexnine_unit ninexnine_unit_3697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A04)
);

ninexnine_unit ninexnine_unit_3698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A04)
);

ninexnine_unit ninexnine_unit_3699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A04)
);

assign C1A04=c10A04+c11A04+c12A04+c13A04;
assign A1A04=(C1A04>=0)?1:0;

ninexnine_unit ninexnine_unit_3700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A14)
);

ninexnine_unit ninexnine_unit_3701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A14)
);

ninexnine_unit ninexnine_unit_3702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A14)
);

ninexnine_unit ninexnine_unit_3703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A14)
);

assign C1A14=c10A14+c11A14+c12A14+c13A14;
assign A1A14=(C1A14>=0)?1:0;

ninexnine_unit ninexnine_unit_3704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A24)
);

ninexnine_unit ninexnine_unit_3705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A24)
);

ninexnine_unit ninexnine_unit_3706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A24)
);

ninexnine_unit ninexnine_unit_3707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A24)
);

assign C1A24=c10A24+c11A24+c12A24+c13A24;
assign A1A24=(C1A24>=0)?1:0;

ninexnine_unit ninexnine_unit_3708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A34)
);

ninexnine_unit ninexnine_unit_3709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A34)
);

ninexnine_unit ninexnine_unit_3710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A34)
);

ninexnine_unit ninexnine_unit_3711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A34)
);

assign C1A34=c10A34+c11A34+c12A34+c13A34;
assign A1A34=(C1A34>=0)?1:0;

ninexnine_unit ninexnine_unit_3712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A44)
);

ninexnine_unit ninexnine_unit_3713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A44)
);

ninexnine_unit ninexnine_unit_3714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A44)
);

ninexnine_unit ninexnine_unit_3715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A44)
);

assign C1A44=c10A44+c11A44+c12A44+c13A44;
assign A1A44=(C1A44>=0)?1:0;

ninexnine_unit ninexnine_unit_3716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A54)
);

ninexnine_unit ninexnine_unit_3717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A54)
);

ninexnine_unit ninexnine_unit_3718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A54)
);

ninexnine_unit ninexnine_unit_3719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A54)
);

assign C1A54=c10A54+c11A54+c12A54+c13A54;
assign A1A54=(C1A54>=0)?1:0;

ninexnine_unit ninexnine_unit_3720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A64)
);

ninexnine_unit ninexnine_unit_3721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A64)
);

ninexnine_unit ninexnine_unit_3722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A64)
);

ninexnine_unit ninexnine_unit_3723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A64)
);

assign C1A64=c10A64+c11A64+c12A64+c13A64;
assign A1A64=(C1A64>=0)?1:0;

ninexnine_unit ninexnine_unit_3724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A74)
);

ninexnine_unit ninexnine_unit_3725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A74)
);

ninexnine_unit ninexnine_unit_3726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A74)
);

ninexnine_unit ninexnine_unit_3727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A74)
);

assign C1A74=c10A74+c11A74+c12A74+c13A74;
assign A1A74=(C1A74>=0)?1:0;

ninexnine_unit ninexnine_unit_3728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A84)
);

ninexnine_unit ninexnine_unit_3729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A84)
);

ninexnine_unit ninexnine_unit_3730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A84)
);

ninexnine_unit ninexnine_unit_3731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A84)
);

assign C1A84=c10A84+c11A84+c12A84+c13A84;
assign A1A84=(C1A84>=0)?1:0;

ninexnine_unit ninexnine_unit_3732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10A94)
);

ninexnine_unit ninexnine_unit_3733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11A94)
);

ninexnine_unit ninexnine_unit_3734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12A94)
);

ninexnine_unit ninexnine_unit_3735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13A94)
);

assign C1A94=c10A94+c11A94+c12A94+c13A94;
assign A1A94=(C1A94>=0)?1:0;

ninexnine_unit ninexnine_unit_3736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10AA4)
);

ninexnine_unit ninexnine_unit_3737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11AA4)
);

ninexnine_unit ninexnine_unit_3738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12AA4)
);

ninexnine_unit ninexnine_unit_3739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13AA4)
);

assign C1AA4=c10AA4+c11AA4+c12AA4+c13AA4;
assign A1AA4=(C1AA4>=0)?1:0;

ninexnine_unit ninexnine_unit_3740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10AB4)
);

ninexnine_unit ninexnine_unit_3741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11AB4)
);

ninexnine_unit ninexnine_unit_3742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12AB4)
);

ninexnine_unit ninexnine_unit_3743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13AB4)
);

assign C1AB4=c10AB4+c11AB4+c12AB4+c13AB4;
assign A1AB4=(C1AB4>=0)?1:0;

ninexnine_unit ninexnine_unit_3744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10AC4)
);

ninexnine_unit ninexnine_unit_3745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11AC4)
);

ninexnine_unit ninexnine_unit_3746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12AC4)
);

ninexnine_unit ninexnine_unit_3747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13AC4)
);

assign C1AC4=c10AC4+c11AC4+c12AC4+c13AC4;
assign A1AC4=(C1AC4>=0)?1:0;

ninexnine_unit ninexnine_unit_3748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10AD4)
);

ninexnine_unit ninexnine_unit_3749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11AD4)
);

ninexnine_unit ninexnine_unit_3750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12AD4)
);

ninexnine_unit ninexnine_unit_3751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13AD4)
);

assign C1AD4=c10AD4+c11AD4+c12AD4+c13AD4;
assign A1AD4=(C1AD4>=0)?1:0;

ninexnine_unit ninexnine_unit_3752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B04)
);

ninexnine_unit ninexnine_unit_3753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B04)
);

ninexnine_unit ninexnine_unit_3754(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B04)
);

ninexnine_unit ninexnine_unit_3755(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B04)
);

assign C1B04=c10B04+c11B04+c12B04+c13B04;
assign A1B04=(C1B04>=0)?1:0;

ninexnine_unit ninexnine_unit_3756(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B14)
);

ninexnine_unit ninexnine_unit_3757(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B14)
);

ninexnine_unit ninexnine_unit_3758(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B14)
);

ninexnine_unit ninexnine_unit_3759(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B14)
);

assign C1B14=c10B14+c11B14+c12B14+c13B14;
assign A1B14=(C1B14>=0)?1:0;

ninexnine_unit ninexnine_unit_3760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B24)
);

ninexnine_unit ninexnine_unit_3761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B24)
);

ninexnine_unit ninexnine_unit_3762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B24)
);

ninexnine_unit ninexnine_unit_3763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B24)
);

assign C1B24=c10B24+c11B24+c12B24+c13B24;
assign A1B24=(C1B24>=0)?1:0;

ninexnine_unit ninexnine_unit_3764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B34)
);

ninexnine_unit ninexnine_unit_3765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B34)
);

ninexnine_unit ninexnine_unit_3766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B34)
);

ninexnine_unit ninexnine_unit_3767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B34)
);

assign C1B34=c10B34+c11B34+c12B34+c13B34;
assign A1B34=(C1B34>=0)?1:0;

ninexnine_unit ninexnine_unit_3768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B44)
);

ninexnine_unit ninexnine_unit_3769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B44)
);

ninexnine_unit ninexnine_unit_3770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B44)
);

ninexnine_unit ninexnine_unit_3771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B44)
);

assign C1B44=c10B44+c11B44+c12B44+c13B44;
assign A1B44=(C1B44>=0)?1:0;

ninexnine_unit ninexnine_unit_3772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B54)
);

ninexnine_unit ninexnine_unit_3773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B54)
);

ninexnine_unit ninexnine_unit_3774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B54)
);

ninexnine_unit ninexnine_unit_3775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B54)
);

assign C1B54=c10B54+c11B54+c12B54+c13B54;
assign A1B54=(C1B54>=0)?1:0;

ninexnine_unit ninexnine_unit_3776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B64)
);

ninexnine_unit ninexnine_unit_3777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B64)
);

ninexnine_unit ninexnine_unit_3778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B64)
);

ninexnine_unit ninexnine_unit_3779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B64)
);

assign C1B64=c10B64+c11B64+c12B64+c13B64;
assign A1B64=(C1B64>=0)?1:0;

ninexnine_unit ninexnine_unit_3780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B74)
);

ninexnine_unit ninexnine_unit_3781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B74)
);

ninexnine_unit ninexnine_unit_3782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B74)
);

ninexnine_unit ninexnine_unit_3783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B74)
);

assign C1B74=c10B74+c11B74+c12B74+c13B74;
assign A1B74=(C1B74>=0)?1:0;

ninexnine_unit ninexnine_unit_3784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B84)
);

ninexnine_unit ninexnine_unit_3785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B84)
);

ninexnine_unit ninexnine_unit_3786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B84)
);

ninexnine_unit ninexnine_unit_3787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B84)
);

assign C1B84=c10B84+c11B84+c12B84+c13B84;
assign A1B84=(C1B84>=0)?1:0;

ninexnine_unit ninexnine_unit_3788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10B94)
);

ninexnine_unit ninexnine_unit_3789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11B94)
);

ninexnine_unit ninexnine_unit_3790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12B94)
);

ninexnine_unit ninexnine_unit_3791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13B94)
);

assign C1B94=c10B94+c11B94+c12B94+c13B94;
assign A1B94=(C1B94>=0)?1:0;

ninexnine_unit ninexnine_unit_3792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10BA4)
);

ninexnine_unit ninexnine_unit_3793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11BA4)
);

ninexnine_unit ninexnine_unit_3794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12BA4)
);

ninexnine_unit ninexnine_unit_3795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13BA4)
);

assign C1BA4=c10BA4+c11BA4+c12BA4+c13BA4;
assign A1BA4=(C1BA4>=0)?1:0;

ninexnine_unit ninexnine_unit_3796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10BB4)
);

ninexnine_unit ninexnine_unit_3797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11BB4)
);

ninexnine_unit ninexnine_unit_3798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12BB4)
);

ninexnine_unit ninexnine_unit_3799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13BB4)
);

assign C1BB4=c10BB4+c11BB4+c12BB4+c13BB4;
assign A1BB4=(C1BB4>=0)?1:0;

ninexnine_unit ninexnine_unit_3800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10BC4)
);

ninexnine_unit ninexnine_unit_3801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11BC4)
);

ninexnine_unit ninexnine_unit_3802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12BC4)
);

ninexnine_unit ninexnine_unit_3803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13BC4)
);

assign C1BC4=c10BC4+c11BC4+c12BC4+c13BC4;
assign A1BC4=(C1BC4>=0)?1:0;

ninexnine_unit ninexnine_unit_3804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10BD4)
);

ninexnine_unit ninexnine_unit_3805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11BD4)
);

ninexnine_unit ninexnine_unit_3806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12BD4)
);

ninexnine_unit ninexnine_unit_3807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13BD4)
);

assign C1BD4=c10BD4+c11BD4+c12BD4+c13BD4;
assign A1BD4=(C1BD4>=0)?1:0;

ninexnine_unit ninexnine_unit_3808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C04)
);

ninexnine_unit ninexnine_unit_3809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C04)
);

ninexnine_unit ninexnine_unit_3810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C04)
);

ninexnine_unit ninexnine_unit_3811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C04)
);

assign C1C04=c10C04+c11C04+c12C04+c13C04;
assign A1C04=(C1C04>=0)?1:0;

ninexnine_unit ninexnine_unit_3812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C14)
);

ninexnine_unit ninexnine_unit_3813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C14)
);

ninexnine_unit ninexnine_unit_3814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C14)
);

ninexnine_unit ninexnine_unit_3815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C14)
);

assign C1C14=c10C14+c11C14+c12C14+c13C14;
assign A1C14=(C1C14>=0)?1:0;

ninexnine_unit ninexnine_unit_3816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C24)
);

ninexnine_unit ninexnine_unit_3817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C24)
);

ninexnine_unit ninexnine_unit_3818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C24)
);

ninexnine_unit ninexnine_unit_3819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C24)
);

assign C1C24=c10C24+c11C24+c12C24+c13C24;
assign A1C24=(C1C24>=0)?1:0;

ninexnine_unit ninexnine_unit_3820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C34)
);

ninexnine_unit ninexnine_unit_3821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C34)
);

ninexnine_unit ninexnine_unit_3822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C34)
);

ninexnine_unit ninexnine_unit_3823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C34)
);

assign C1C34=c10C34+c11C34+c12C34+c13C34;
assign A1C34=(C1C34>=0)?1:0;

ninexnine_unit ninexnine_unit_3824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C44)
);

ninexnine_unit ninexnine_unit_3825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C44)
);

ninexnine_unit ninexnine_unit_3826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C44)
);

ninexnine_unit ninexnine_unit_3827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C44)
);

assign C1C44=c10C44+c11C44+c12C44+c13C44;
assign A1C44=(C1C44>=0)?1:0;

ninexnine_unit ninexnine_unit_3828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C54)
);

ninexnine_unit ninexnine_unit_3829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C54)
);

ninexnine_unit ninexnine_unit_3830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C54)
);

ninexnine_unit ninexnine_unit_3831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C54)
);

assign C1C54=c10C54+c11C54+c12C54+c13C54;
assign A1C54=(C1C54>=0)?1:0;

ninexnine_unit ninexnine_unit_3832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C64)
);

ninexnine_unit ninexnine_unit_3833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C64)
);

ninexnine_unit ninexnine_unit_3834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C64)
);

ninexnine_unit ninexnine_unit_3835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C64)
);

assign C1C64=c10C64+c11C64+c12C64+c13C64;
assign A1C64=(C1C64>=0)?1:0;

ninexnine_unit ninexnine_unit_3836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C74)
);

ninexnine_unit ninexnine_unit_3837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C74)
);

ninexnine_unit ninexnine_unit_3838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C74)
);

ninexnine_unit ninexnine_unit_3839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C74)
);

assign C1C74=c10C74+c11C74+c12C74+c13C74;
assign A1C74=(C1C74>=0)?1:0;

ninexnine_unit ninexnine_unit_3840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C84)
);

ninexnine_unit ninexnine_unit_3841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C84)
);

ninexnine_unit ninexnine_unit_3842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C84)
);

ninexnine_unit ninexnine_unit_3843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C84)
);

assign C1C84=c10C84+c11C84+c12C84+c13C84;
assign A1C84=(C1C84>=0)?1:0;

ninexnine_unit ninexnine_unit_3844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10C94)
);

ninexnine_unit ninexnine_unit_3845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11C94)
);

ninexnine_unit ninexnine_unit_3846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12C94)
);

ninexnine_unit ninexnine_unit_3847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13C94)
);

assign C1C94=c10C94+c11C94+c12C94+c13C94;
assign A1C94=(C1C94>=0)?1:0;

ninexnine_unit ninexnine_unit_3848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10CA4)
);

ninexnine_unit ninexnine_unit_3849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11CA4)
);

ninexnine_unit ninexnine_unit_3850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12CA4)
);

ninexnine_unit ninexnine_unit_3851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13CA4)
);

assign C1CA4=c10CA4+c11CA4+c12CA4+c13CA4;
assign A1CA4=(C1CA4>=0)?1:0;

ninexnine_unit ninexnine_unit_3852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10CB4)
);

ninexnine_unit ninexnine_unit_3853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11CB4)
);

ninexnine_unit ninexnine_unit_3854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12CB4)
);

ninexnine_unit ninexnine_unit_3855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13CB4)
);

assign C1CB4=c10CB4+c11CB4+c12CB4+c13CB4;
assign A1CB4=(C1CB4>=0)?1:0;

ninexnine_unit ninexnine_unit_3856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10CC4)
);

ninexnine_unit ninexnine_unit_3857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11CC4)
);

ninexnine_unit ninexnine_unit_3858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12CC4)
);

ninexnine_unit ninexnine_unit_3859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13CC4)
);

assign C1CC4=c10CC4+c11CC4+c12CC4+c13CC4;
assign A1CC4=(C1CC4>=0)?1:0;

ninexnine_unit ninexnine_unit_3860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10CD4)
);

ninexnine_unit ninexnine_unit_3861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11CD4)
);

ninexnine_unit ninexnine_unit_3862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12CD4)
);

ninexnine_unit ninexnine_unit_3863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13CD4)
);

assign C1CD4=c10CD4+c11CD4+c12CD4+c13CD4;
assign A1CD4=(C1CD4>=0)?1:0;

ninexnine_unit ninexnine_unit_3864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D04)
);

ninexnine_unit ninexnine_unit_3865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D04)
);

ninexnine_unit ninexnine_unit_3866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D04)
);

ninexnine_unit ninexnine_unit_3867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D04)
);

assign C1D04=c10D04+c11D04+c12D04+c13D04;
assign A1D04=(C1D04>=0)?1:0;

ninexnine_unit ninexnine_unit_3868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D14)
);

ninexnine_unit ninexnine_unit_3869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D14)
);

ninexnine_unit ninexnine_unit_3870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D14)
);

ninexnine_unit ninexnine_unit_3871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D14)
);

assign C1D14=c10D14+c11D14+c12D14+c13D14;
assign A1D14=(C1D14>=0)?1:0;

ninexnine_unit ninexnine_unit_3872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D24)
);

ninexnine_unit ninexnine_unit_3873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D24)
);

ninexnine_unit ninexnine_unit_3874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D24)
);

ninexnine_unit ninexnine_unit_3875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D24)
);

assign C1D24=c10D24+c11D24+c12D24+c13D24;
assign A1D24=(C1D24>=0)?1:0;

ninexnine_unit ninexnine_unit_3876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D34)
);

ninexnine_unit ninexnine_unit_3877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D34)
);

ninexnine_unit ninexnine_unit_3878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D34)
);

ninexnine_unit ninexnine_unit_3879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D34)
);

assign C1D34=c10D34+c11D34+c12D34+c13D34;
assign A1D34=(C1D34>=0)?1:0;

ninexnine_unit ninexnine_unit_3880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D44)
);

ninexnine_unit ninexnine_unit_3881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D44)
);

ninexnine_unit ninexnine_unit_3882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D44)
);

ninexnine_unit ninexnine_unit_3883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D44)
);

assign C1D44=c10D44+c11D44+c12D44+c13D44;
assign A1D44=(C1D44>=0)?1:0;

ninexnine_unit ninexnine_unit_3884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D54)
);

ninexnine_unit ninexnine_unit_3885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D54)
);

ninexnine_unit ninexnine_unit_3886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D54)
);

ninexnine_unit ninexnine_unit_3887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D54)
);

assign C1D54=c10D54+c11D54+c12D54+c13D54;
assign A1D54=(C1D54>=0)?1:0;

ninexnine_unit ninexnine_unit_3888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D64)
);

ninexnine_unit ninexnine_unit_3889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D64)
);

ninexnine_unit ninexnine_unit_3890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D64)
);

ninexnine_unit ninexnine_unit_3891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D64)
);

assign C1D64=c10D64+c11D64+c12D64+c13D64;
assign A1D64=(C1D64>=0)?1:0;

ninexnine_unit ninexnine_unit_3892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D74)
);

ninexnine_unit ninexnine_unit_3893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D74)
);

ninexnine_unit ninexnine_unit_3894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D74)
);

ninexnine_unit ninexnine_unit_3895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D74)
);

assign C1D74=c10D74+c11D74+c12D74+c13D74;
assign A1D74=(C1D74>=0)?1:0;

ninexnine_unit ninexnine_unit_3896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D84)
);

ninexnine_unit ninexnine_unit_3897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D84)
);

ninexnine_unit ninexnine_unit_3898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D84)
);

ninexnine_unit ninexnine_unit_3899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D84)
);

assign C1D84=c10D84+c11D84+c12D84+c13D84;
assign A1D84=(C1D84>=0)?1:0;

ninexnine_unit ninexnine_unit_3900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10D94)
);

ninexnine_unit ninexnine_unit_3901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11D94)
);

ninexnine_unit ninexnine_unit_3902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12D94)
);

ninexnine_unit ninexnine_unit_3903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13D94)
);

assign C1D94=c10D94+c11D94+c12D94+c13D94;
assign A1D94=(C1D94>=0)?1:0;

ninexnine_unit ninexnine_unit_3904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10DA4)
);

ninexnine_unit ninexnine_unit_3905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11DA4)
);

ninexnine_unit ninexnine_unit_3906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12DA4)
);

ninexnine_unit ninexnine_unit_3907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13DA4)
);

assign C1DA4=c10DA4+c11DA4+c12DA4+c13DA4;
assign A1DA4=(C1DA4>=0)?1:0;

ninexnine_unit ninexnine_unit_3908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10DB4)
);

ninexnine_unit ninexnine_unit_3909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11DB4)
);

ninexnine_unit ninexnine_unit_3910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12DB4)
);

ninexnine_unit ninexnine_unit_3911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13DB4)
);

assign C1DB4=c10DB4+c11DB4+c12DB4+c13DB4;
assign A1DB4=(C1DB4>=0)?1:0;

ninexnine_unit ninexnine_unit_3912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10DC4)
);

ninexnine_unit ninexnine_unit_3913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11DC4)
);

ninexnine_unit ninexnine_unit_3914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12DC4)
);

ninexnine_unit ninexnine_unit_3915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13DC4)
);

assign C1DC4=c10DC4+c11DC4+c12DC4+c13DC4;
assign A1DC4=(C1DC4>=0)?1:0;

ninexnine_unit ninexnine_unit_3916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10DD4)
);

ninexnine_unit ninexnine_unit_3917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11DD4)
);

ninexnine_unit ninexnine_unit_3918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12DD4)
);

ninexnine_unit ninexnine_unit_3919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13DD4)
);

assign C1DD4=c10DD4+c11DD4+c12DD4+c13DD4;
assign A1DD4=(C1DD4>=0)?1:0;

ninexnine_unit ninexnine_unit_3920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10005)
);

ninexnine_unit ninexnine_unit_3921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11005)
);

ninexnine_unit ninexnine_unit_3922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12005)
);

ninexnine_unit ninexnine_unit_3923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13005)
);

assign C1005=c10005+c11005+c12005+c13005;
assign A1005=(C1005>=0)?1:0;

ninexnine_unit ninexnine_unit_3924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10015)
);

ninexnine_unit ninexnine_unit_3925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11015)
);

ninexnine_unit ninexnine_unit_3926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12015)
);

ninexnine_unit ninexnine_unit_3927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13015)
);

assign C1015=c10015+c11015+c12015+c13015;
assign A1015=(C1015>=0)?1:0;

ninexnine_unit ninexnine_unit_3928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10025)
);

ninexnine_unit ninexnine_unit_3929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11025)
);

ninexnine_unit ninexnine_unit_3930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12025)
);

ninexnine_unit ninexnine_unit_3931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13025)
);

assign C1025=c10025+c11025+c12025+c13025;
assign A1025=(C1025>=0)?1:0;

ninexnine_unit ninexnine_unit_3932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10035)
);

ninexnine_unit ninexnine_unit_3933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11035)
);

ninexnine_unit ninexnine_unit_3934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12035)
);

ninexnine_unit ninexnine_unit_3935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13035)
);

assign C1035=c10035+c11035+c12035+c13035;
assign A1035=(C1035>=0)?1:0;

ninexnine_unit ninexnine_unit_3936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10045)
);

ninexnine_unit ninexnine_unit_3937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11045)
);

ninexnine_unit ninexnine_unit_3938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12045)
);

ninexnine_unit ninexnine_unit_3939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13045)
);

assign C1045=c10045+c11045+c12045+c13045;
assign A1045=(C1045>=0)?1:0;

ninexnine_unit ninexnine_unit_3940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10055)
);

ninexnine_unit ninexnine_unit_3941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11055)
);

ninexnine_unit ninexnine_unit_3942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12055)
);

ninexnine_unit ninexnine_unit_3943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13055)
);

assign C1055=c10055+c11055+c12055+c13055;
assign A1055=(C1055>=0)?1:0;

ninexnine_unit ninexnine_unit_3944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10065)
);

ninexnine_unit ninexnine_unit_3945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11065)
);

ninexnine_unit ninexnine_unit_3946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12065)
);

ninexnine_unit ninexnine_unit_3947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13065)
);

assign C1065=c10065+c11065+c12065+c13065;
assign A1065=(C1065>=0)?1:0;

ninexnine_unit ninexnine_unit_3948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10075)
);

ninexnine_unit ninexnine_unit_3949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11075)
);

ninexnine_unit ninexnine_unit_3950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12075)
);

ninexnine_unit ninexnine_unit_3951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13075)
);

assign C1075=c10075+c11075+c12075+c13075;
assign A1075=(C1075>=0)?1:0;

ninexnine_unit ninexnine_unit_3952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10085)
);

ninexnine_unit ninexnine_unit_3953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11085)
);

ninexnine_unit ninexnine_unit_3954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12085)
);

ninexnine_unit ninexnine_unit_3955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13085)
);

assign C1085=c10085+c11085+c12085+c13085;
assign A1085=(C1085>=0)?1:0;

ninexnine_unit ninexnine_unit_3956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10095)
);

ninexnine_unit ninexnine_unit_3957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11095)
);

ninexnine_unit ninexnine_unit_3958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12095)
);

ninexnine_unit ninexnine_unit_3959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13095)
);

assign C1095=c10095+c11095+c12095+c13095;
assign A1095=(C1095>=0)?1:0;

ninexnine_unit ninexnine_unit_3960(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c100A5)
);

ninexnine_unit ninexnine_unit_3961(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c110A5)
);

ninexnine_unit ninexnine_unit_3962(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c120A5)
);

ninexnine_unit ninexnine_unit_3963(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c130A5)
);

assign C10A5=c100A5+c110A5+c120A5+c130A5;
assign A10A5=(C10A5>=0)?1:0;

ninexnine_unit ninexnine_unit_3964(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c100B5)
);

ninexnine_unit ninexnine_unit_3965(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c110B5)
);

ninexnine_unit ninexnine_unit_3966(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c120B5)
);

ninexnine_unit ninexnine_unit_3967(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c130B5)
);

assign C10B5=c100B5+c110B5+c120B5+c130B5;
assign A10B5=(C10B5>=0)?1:0;

ninexnine_unit ninexnine_unit_3968(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c100C5)
);

ninexnine_unit ninexnine_unit_3969(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c110C5)
);

ninexnine_unit ninexnine_unit_3970(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c120C5)
);

ninexnine_unit ninexnine_unit_3971(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c130C5)
);

assign C10C5=c100C5+c110C5+c120C5+c130C5;
assign A10C5=(C10C5>=0)?1:0;

ninexnine_unit ninexnine_unit_3972(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c100D5)
);

ninexnine_unit ninexnine_unit_3973(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c110D5)
);

ninexnine_unit ninexnine_unit_3974(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c120D5)
);

ninexnine_unit ninexnine_unit_3975(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c130D5)
);

assign C10D5=c100D5+c110D5+c120D5+c130D5;
assign A10D5=(C10D5>=0)?1:0;

ninexnine_unit ninexnine_unit_3976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10105)
);

ninexnine_unit ninexnine_unit_3977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11105)
);

ninexnine_unit ninexnine_unit_3978(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12105)
);

ninexnine_unit ninexnine_unit_3979(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13105)
);

assign C1105=c10105+c11105+c12105+c13105;
assign A1105=(C1105>=0)?1:0;

ninexnine_unit ninexnine_unit_3980(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10115)
);

ninexnine_unit ninexnine_unit_3981(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11115)
);

ninexnine_unit ninexnine_unit_3982(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12115)
);

ninexnine_unit ninexnine_unit_3983(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13115)
);

assign C1115=c10115+c11115+c12115+c13115;
assign A1115=(C1115>=0)?1:0;

ninexnine_unit ninexnine_unit_3984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10125)
);

ninexnine_unit ninexnine_unit_3985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11125)
);

ninexnine_unit ninexnine_unit_3986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12125)
);

ninexnine_unit ninexnine_unit_3987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13125)
);

assign C1125=c10125+c11125+c12125+c13125;
assign A1125=(C1125>=0)?1:0;

ninexnine_unit ninexnine_unit_3988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10135)
);

ninexnine_unit ninexnine_unit_3989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11135)
);

ninexnine_unit ninexnine_unit_3990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12135)
);

ninexnine_unit ninexnine_unit_3991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13135)
);

assign C1135=c10135+c11135+c12135+c13135;
assign A1135=(C1135>=0)?1:0;

ninexnine_unit ninexnine_unit_3992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10145)
);

ninexnine_unit ninexnine_unit_3993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11145)
);

ninexnine_unit ninexnine_unit_3994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12145)
);

ninexnine_unit ninexnine_unit_3995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13145)
);

assign C1145=c10145+c11145+c12145+c13145;
assign A1145=(C1145>=0)?1:0;

ninexnine_unit ninexnine_unit_3996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10155)
);

ninexnine_unit ninexnine_unit_3997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11155)
);

ninexnine_unit ninexnine_unit_3998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12155)
);

ninexnine_unit ninexnine_unit_3999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13155)
);

assign C1155=c10155+c11155+c12155+c13155;
assign A1155=(C1155>=0)?1:0;

ninexnine_unit ninexnine_unit_4000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10165)
);

ninexnine_unit ninexnine_unit_4001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11165)
);

ninexnine_unit ninexnine_unit_4002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12165)
);

ninexnine_unit ninexnine_unit_4003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13165)
);

assign C1165=c10165+c11165+c12165+c13165;
assign A1165=(C1165>=0)?1:0;

ninexnine_unit ninexnine_unit_4004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10175)
);

ninexnine_unit ninexnine_unit_4005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11175)
);

ninexnine_unit ninexnine_unit_4006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12175)
);

ninexnine_unit ninexnine_unit_4007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13175)
);

assign C1175=c10175+c11175+c12175+c13175;
assign A1175=(C1175>=0)?1:0;

ninexnine_unit ninexnine_unit_4008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10185)
);

ninexnine_unit ninexnine_unit_4009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11185)
);

ninexnine_unit ninexnine_unit_4010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12185)
);

ninexnine_unit ninexnine_unit_4011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13185)
);

assign C1185=c10185+c11185+c12185+c13185;
assign A1185=(C1185>=0)?1:0;

ninexnine_unit ninexnine_unit_4012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10195)
);

ninexnine_unit ninexnine_unit_4013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11195)
);

ninexnine_unit ninexnine_unit_4014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12195)
);

ninexnine_unit ninexnine_unit_4015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13195)
);

assign C1195=c10195+c11195+c12195+c13195;
assign A1195=(C1195>=0)?1:0;

ninexnine_unit ninexnine_unit_4016(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c101A5)
);

ninexnine_unit ninexnine_unit_4017(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c111A5)
);

ninexnine_unit ninexnine_unit_4018(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c121A5)
);

ninexnine_unit ninexnine_unit_4019(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c131A5)
);

assign C11A5=c101A5+c111A5+c121A5+c131A5;
assign A11A5=(C11A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4020(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c101B5)
);

ninexnine_unit ninexnine_unit_4021(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c111B5)
);

ninexnine_unit ninexnine_unit_4022(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c121B5)
);

ninexnine_unit ninexnine_unit_4023(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c131B5)
);

assign C11B5=c101B5+c111B5+c121B5+c131B5;
assign A11B5=(C11B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4024(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c101C5)
);

ninexnine_unit ninexnine_unit_4025(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c111C5)
);

ninexnine_unit ninexnine_unit_4026(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c121C5)
);

ninexnine_unit ninexnine_unit_4027(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c131C5)
);

assign C11C5=c101C5+c111C5+c121C5+c131C5;
assign A11C5=(C11C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4028(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c101D5)
);

ninexnine_unit ninexnine_unit_4029(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c111D5)
);

ninexnine_unit ninexnine_unit_4030(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c121D5)
);

ninexnine_unit ninexnine_unit_4031(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c131D5)
);

assign C11D5=c101D5+c111D5+c121D5+c131D5;
assign A11D5=(C11D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10205)
);

ninexnine_unit ninexnine_unit_4033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11205)
);

ninexnine_unit ninexnine_unit_4034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12205)
);

ninexnine_unit ninexnine_unit_4035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13205)
);

assign C1205=c10205+c11205+c12205+c13205;
assign A1205=(C1205>=0)?1:0;

ninexnine_unit ninexnine_unit_4036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10215)
);

ninexnine_unit ninexnine_unit_4037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11215)
);

ninexnine_unit ninexnine_unit_4038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12215)
);

ninexnine_unit ninexnine_unit_4039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13215)
);

assign C1215=c10215+c11215+c12215+c13215;
assign A1215=(C1215>=0)?1:0;

ninexnine_unit ninexnine_unit_4040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10225)
);

ninexnine_unit ninexnine_unit_4041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11225)
);

ninexnine_unit ninexnine_unit_4042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12225)
);

ninexnine_unit ninexnine_unit_4043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13225)
);

assign C1225=c10225+c11225+c12225+c13225;
assign A1225=(C1225>=0)?1:0;

ninexnine_unit ninexnine_unit_4044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10235)
);

ninexnine_unit ninexnine_unit_4045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11235)
);

ninexnine_unit ninexnine_unit_4046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12235)
);

ninexnine_unit ninexnine_unit_4047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13235)
);

assign C1235=c10235+c11235+c12235+c13235;
assign A1235=(C1235>=0)?1:0;

ninexnine_unit ninexnine_unit_4048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10245)
);

ninexnine_unit ninexnine_unit_4049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11245)
);

ninexnine_unit ninexnine_unit_4050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12245)
);

ninexnine_unit ninexnine_unit_4051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13245)
);

assign C1245=c10245+c11245+c12245+c13245;
assign A1245=(C1245>=0)?1:0;

ninexnine_unit ninexnine_unit_4052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10255)
);

ninexnine_unit ninexnine_unit_4053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11255)
);

ninexnine_unit ninexnine_unit_4054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12255)
);

ninexnine_unit ninexnine_unit_4055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13255)
);

assign C1255=c10255+c11255+c12255+c13255;
assign A1255=(C1255>=0)?1:0;

ninexnine_unit ninexnine_unit_4056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10265)
);

ninexnine_unit ninexnine_unit_4057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11265)
);

ninexnine_unit ninexnine_unit_4058(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12265)
);

ninexnine_unit ninexnine_unit_4059(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13265)
);

assign C1265=c10265+c11265+c12265+c13265;
assign A1265=(C1265>=0)?1:0;

ninexnine_unit ninexnine_unit_4060(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10275)
);

ninexnine_unit ninexnine_unit_4061(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11275)
);

ninexnine_unit ninexnine_unit_4062(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12275)
);

ninexnine_unit ninexnine_unit_4063(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13275)
);

assign C1275=c10275+c11275+c12275+c13275;
assign A1275=(C1275>=0)?1:0;

ninexnine_unit ninexnine_unit_4064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10285)
);

ninexnine_unit ninexnine_unit_4065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11285)
);

ninexnine_unit ninexnine_unit_4066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12285)
);

ninexnine_unit ninexnine_unit_4067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13285)
);

assign C1285=c10285+c11285+c12285+c13285;
assign A1285=(C1285>=0)?1:0;

ninexnine_unit ninexnine_unit_4068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10295)
);

ninexnine_unit ninexnine_unit_4069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11295)
);

ninexnine_unit ninexnine_unit_4070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12295)
);

ninexnine_unit ninexnine_unit_4071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13295)
);

assign C1295=c10295+c11295+c12295+c13295;
assign A1295=(C1295>=0)?1:0;

ninexnine_unit ninexnine_unit_4072(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c102A5)
);

ninexnine_unit ninexnine_unit_4073(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c112A5)
);

ninexnine_unit ninexnine_unit_4074(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c122A5)
);

ninexnine_unit ninexnine_unit_4075(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c132A5)
);

assign C12A5=c102A5+c112A5+c122A5+c132A5;
assign A12A5=(C12A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4076(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c102B5)
);

ninexnine_unit ninexnine_unit_4077(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c112B5)
);

ninexnine_unit ninexnine_unit_4078(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c122B5)
);

ninexnine_unit ninexnine_unit_4079(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c132B5)
);

assign C12B5=c102B5+c112B5+c122B5+c132B5;
assign A12B5=(C12B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4080(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c102C5)
);

ninexnine_unit ninexnine_unit_4081(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c112C5)
);

ninexnine_unit ninexnine_unit_4082(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c122C5)
);

ninexnine_unit ninexnine_unit_4083(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c132C5)
);

assign C12C5=c102C5+c112C5+c122C5+c132C5;
assign A12C5=(C12C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4084(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c102D5)
);

ninexnine_unit ninexnine_unit_4085(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c112D5)
);

ninexnine_unit ninexnine_unit_4086(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c122D5)
);

ninexnine_unit ninexnine_unit_4087(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c132D5)
);

assign C12D5=c102D5+c112D5+c122D5+c132D5;
assign A12D5=(C12D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10305)
);

ninexnine_unit ninexnine_unit_4089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11305)
);

ninexnine_unit ninexnine_unit_4090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12305)
);

ninexnine_unit ninexnine_unit_4091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13305)
);

assign C1305=c10305+c11305+c12305+c13305;
assign A1305=(C1305>=0)?1:0;

ninexnine_unit ninexnine_unit_4092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10315)
);

ninexnine_unit ninexnine_unit_4093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11315)
);

ninexnine_unit ninexnine_unit_4094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12315)
);

ninexnine_unit ninexnine_unit_4095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13315)
);

assign C1315=c10315+c11315+c12315+c13315;
assign A1315=(C1315>=0)?1:0;

ninexnine_unit ninexnine_unit_4096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10325)
);

ninexnine_unit ninexnine_unit_4097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11325)
);

ninexnine_unit ninexnine_unit_4098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12325)
);

ninexnine_unit ninexnine_unit_4099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13325)
);

assign C1325=c10325+c11325+c12325+c13325;
assign A1325=(C1325>=0)?1:0;

ninexnine_unit ninexnine_unit_4100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10335)
);

ninexnine_unit ninexnine_unit_4101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11335)
);

ninexnine_unit ninexnine_unit_4102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12335)
);

ninexnine_unit ninexnine_unit_4103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13335)
);

assign C1335=c10335+c11335+c12335+c13335;
assign A1335=(C1335>=0)?1:0;

ninexnine_unit ninexnine_unit_4104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10345)
);

ninexnine_unit ninexnine_unit_4105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11345)
);

ninexnine_unit ninexnine_unit_4106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12345)
);

ninexnine_unit ninexnine_unit_4107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13345)
);

assign C1345=c10345+c11345+c12345+c13345;
assign A1345=(C1345>=0)?1:0;

ninexnine_unit ninexnine_unit_4108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10355)
);

ninexnine_unit ninexnine_unit_4109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11355)
);

ninexnine_unit ninexnine_unit_4110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12355)
);

ninexnine_unit ninexnine_unit_4111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13355)
);

assign C1355=c10355+c11355+c12355+c13355;
assign A1355=(C1355>=0)?1:0;

ninexnine_unit ninexnine_unit_4112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10365)
);

ninexnine_unit ninexnine_unit_4113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11365)
);

ninexnine_unit ninexnine_unit_4114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12365)
);

ninexnine_unit ninexnine_unit_4115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13365)
);

assign C1365=c10365+c11365+c12365+c13365;
assign A1365=(C1365>=0)?1:0;

ninexnine_unit ninexnine_unit_4116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10375)
);

ninexnine_unit ninexnine_unit_4117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11375)
);

ninexnine_unit ninexnine_unit_4118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12375)
);

ninexnine_unit ninexnine_unit_4119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13375)
);

assign C1375=c10375+c11375+c12375+c13375;
assign A1375=(C1375>=0)?1:0;

ninexnine_unit ninexnine_unit_4120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10385)
);

ninexnine_unit ninexnine_unit_4121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11385)
);

ninexnine_unit ninexnine_unit_4122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12385)
);

ninexnine_unit ninexnine_unit_4123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13385)
);

assign C1385=c10385+c11385+c12385+c13385;
assign A1385=(C1385>=0)?1:0;

ninexnine_unit ninexnine_unit_4124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10395)
);

ninexnine_unit ninexnine_unit_4125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11395)
);

ninexnine_unit ninexnine_unit_4126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12395)
);

ninexnine_unit ninexnine_unit_4127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13395)
);

assign C1395=c10395+c11395+c12395+c13395;
assign A1395=(C1395>=0)?1:0;

ninexnine_unit ninexnine_unit_4128(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c103A5)
);

ninexnine_unit ninexnine_unit_4129(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c113A5)
);

ninexnine_unit ninexnine_unit_4130(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c123A5)
);

ninexnine_unit ninexnine_unit_4131(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c133A5)
);

assign C13A5=c103A5+c113A5+c123A5+c133A5;
assign A13A5=(C13A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4132(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c103B5)
);

ninexnine_unit ninexnine_unit_4133(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c113B5)
);

ninexnine_unit ninexnine_unit_4134(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c123B5)
);

ninexnine_unit ninexnine_unit_4135(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c133B5)
);

assign C13B5=c103B5+c113B5+c123B5+c133B5;
assign A13B5=(C13B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4136(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c103C5)
);

ninexnine_unit ninexnine_unit_4137(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c113C5)
);

ninexnine_unit ninexnine_unit_4138(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c123C5)
);

ninexnine_unit ninexnine_unit_4139(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c133C5)
);

assign C13C5=c103C5+c113C5+c123C5+c133C5;
assign A13C5=(C13C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4140(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c103D5)
);

ninexnine_unit ninexnine_unit_4141(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c113D5)
);

ninexnine_unit ninexnine_unit_4142(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c123D5)
);

ninexnine_unit ninexnine_unit_4143(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c133D5)
);

assign C13D5=c103D5+c113D5+c123D5+c133D5;
assign A13D5=(C13D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10405)
);

ninexnine_unit ninexnine_unit_4145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11405)
);

ninexnine_unit ninexnine_unit_4146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12405)
);

ninexnine_unit ninexnine_unit_4147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13405)
);

assign C1405=c10405+c11405+c12405+c13405;
assign A1405=(C1405>=0)?1:0;

ninexnine_unit ninexnine_unit_4148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10415)
);

ninexnine_unit ninexnine_unit_4149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11415)
);

ninexnine_unit ninexnine_unit_4150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12415)
);

ninexnine_unit ninexnine_unit_4151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13415)
);

assign C1415=c10415+c11415+c12415+c13415;
assign A1415=(C1415>=0)?1:0;

ninexnine_unit ninexnine_unit_4152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10425)
);

ninexnine_unit ninexnine_unit_4153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11425)
);

ninexnine_unit ninexnine_unit_4154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12425)
);

ninexnine_unit ninexnine_unit_4155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13425)
);

assign C1425=c10425+c11425+c12425+c13425;
assign A1425=(C1425>=0)?1:0;

ninexnine_unit ninexnine_unit_4156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10435)
);

ninexnine_unit ninexnine_unit_4157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11435)
);

ninexnine_unit ninexnine_unit_4158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12435)
);

ninexnine_unit ninexnine_unit_4159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13435)
);

assign C1435=c10435+c11435+c12435+c13435;
assign A1435=(C1435>=0)?1:0;

ninexnine_unit ninexnine_unit_4160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10445)
);

ninexnine_unit ninexnine_unit_4161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11445)
);

ninexnine_unit ninexnine_unit_4162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12445)
);

ninexnine_unit ninexnine_unit_4163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13445)
);

assign C1445=c10445+c11445+c12445+c13445;
assign A1445=(C1445>=0)?1:0;

ninexnine_unit ninexnine_unit_4164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10455)
);

ninexnine_unit ninexnine_unit_4165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11455)
);

ninexnine_unit ninexnine_unit_4166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12455)
);

ninexnine_unit ninexnine_unit_4167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13455)
);

assign C1455=c10455+c11455+c12455+c13455;
assign A1455=(C1455>=0)?1:0;

ninexnine_unit ninexnine_unit_4168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10465)
);

ninexnine_unit ninexnine_unit_4169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11465)
);

ninexnine_unit ninexnine_unit_4170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12465)
);

ninexnine_unit ninexnine_unit_4171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13465)
);

assign C1465=c10465+c11465+c12465+c13465;
assign A1465=(C1465>=0)?1:0;

ninexnine_unit ninexnine_unit_4172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10475)
);

ninexnine_unit ninexnine_unit_4173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11475)
);

ninexnine_unit ninexnine_unit_4174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12475)
);

ninexnine_unit ninexnine_unit_4175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13475)
);

assign C1475=c10475+c11475+c12475+c13475;
assign A1475=(C1475>=0)?1:0;

ninexnine_unit ninexnine_unit_4176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10485)
);

ninexnine_unit ninexnine_unit_4177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11485)
);

ninexnine_unit ninexnine_unit_4178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12485)
);

ninexnine_unit ninexnine_unit_4179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13485)
);

assign C1485=c10485+c11485+c12485+c13485;
assign A1485=(C1485>=0)?1:0;

ninexnine_unit ninexnine_unit_4180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10495)
);

ninexnine_unit ninexnine_unit_4181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11495)
);

ninexnine_unit ninexnine_unit_4182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12495)
);

ninexnine_unit ninexnine_unit_4183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13495)
);

assign C1495=c10495+c11495+c12495+c13495;
assign A1495=(C1495>=0)?1:0;

ninexnine_unit ninexnine_unit_4184(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c104A5)
);

ninexnine_unit ninexnine_unit_4185(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c114A5)
);

ninexnine_unit ninexnine_unit_4186(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c124A5)
);

ninexnine_unit ninexnine_unit_4187(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c134A5)
);

assign C14A5=c104A5+c114A5+c124A5+c134A5;
assign A14A5=(C14A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4188(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c104B5)
);

ninexnine_unit ninexnine_unit_4189(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c114B5)
);

ninexnine_unit ninexnine_unit_4190(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c124B5)
);

ninexnine_unit ninexnine_unit_4191(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c134B5)
);

assign C14B5=c104B5+c114B5+c124B5+c134B5;
assign A14B5=(C14B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4192(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c104C5)
);

ninexnine_unit ninexnine_unit_4193(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c114C5)
);

ninexnine_unit ninexnine_unit_4194(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c124C5)
);

ninexnine_unit ninexnine_unit_4195(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c134C5)
);

assign C14C5=c104C5+c114C5+c124C5+c134C5;
assign A14C5=(C14C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4196(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c104D5)
);

ninexnine_unit ninexnine_unit_4197(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c114D5)
);

ninexnine_unit ninexnine_unit_4198(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c124D5)
);

ninexnine_unit ninexnine_unit_4199(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c134D5)
);

assign C14D5=c104D5+c114D5+c124D5+c134D5;
assign A14D5=(C14D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10505)
);

ninexnine_unit ninexnine_unit_4201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11505)
);

ninexnine_unit ninexnine_unit_4202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12505)
);

ninexnine_unit ninexnine_unit_4203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13505)
);

assign C1505=c10505+c11505+c12505+c13505;
assign A1505=(C1505>=0)?1:0;

ninexnine_unit ninexnine_unit_4204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10515)
);

ninexnine_unit ninexnine_unit_4205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11515)
);

ninexnine_unit ninexnine_unit_4206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12515)
);

ninexnine_unit ninexnine_unit_4207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13515)
);

assign C1515=c10515+c11515+c12515+c13515;
assign A1515=(C1515>=0)?1:0;

ninexnine_unit ninexnine_unit_4208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10525)
);

ninexnine_unit ninexnine_unit_4209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11525)
);

ninexnine_unit ninexnine_unit_4210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12525)
);

ninexnine_unit ninexnine_unit_4211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13525)
);

assign C1525=c10525+c11525+c12525+c13525;
assign A1525=(C1525>=0)?1:0;

ninexnine_unit ninexnine_unit_4212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10535)
);

ninexnine_unit ninexnine_unit_4213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11535)
);

ninexnine_unit ninexnine_unit_4214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12535)
);

ninexnine_unit ninexnine_unit_4215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13535)
);

assign C1535=c10535+c11535+c12535+c13535;
assign A1535=(C1535>=0)?1:0;

ninexnine_unit ninexnine_unit_4216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10545)
);

ninexnine_unit ninexnine_unit_4217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11545)
);

ninexnine_unit ninexnine_unit_4218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12545)
);

ninexnine_unit ninexnine_unit_4219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13545)
);

assign C1545=c10545+c11545+c12545+c13545;
assign A1545=(C1545>=0)?1:0;

ninexnine_unit ninexnine_unit_4220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10555)
);

ninexnine_unit ninexnine_unit_4221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11555)
);

ninexnine_unit ninexnine_unit_4222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12555)
);

ninexnine_unit ninexnine_unit_4223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13555)
);

assign C1555=c10555+c11555+c12555+c13555;
assign A1555=(C1555>=0)?1:0;

ninexnine_unit ninexnine_unit_4224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10565)
);

ninexnine_unit ninexnine_unit_4225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11565)
);

ninexnine_unit ninexnine_unit_4226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12565)
);

ninexnine_unit ninexnine_unit_4227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13565)
);

assign C1565=c10565+c11565+c12565+c13565;
assign A1565=(C1565>=0)?1:0;

ninexnine_unit ninexnine_unit_4228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10575)
);

ninexnine_unit ninexnine_unit_4229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11575)
);

ninexnine_unit ninexnine_unit_4230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12575)
);

ninexnine_unit ninexnine_unit_4231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13575)
);

assign C1575=c10575+c11575+c12575+c13575;
assign A1575=(C1575>=0)?1:0;

ninexnine_unit ninexnine_unit_4232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10585)
);

ninexnine_unit ninexnine_unit_4233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11585)
);

ninexnine_unit ninexnine_unit_4234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12585)
);

ninexnine_unit ninexnine_unit_4235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13585)
);

assign C1585=c10585+c11585+c12585+c13585;
assign A1585=(C1585>=0)?1:0;

ninexnine_unit ninexnine_unit_4236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10595)
);

ninexnine_unit ninexnine_unit_4237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11595)
);

ninexnine_unit ninexnine_unit_4238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12595)
);

ninexnine_unit ninexnine_unit_4239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13595)
);

assign C1595=c10595+c11595+c12595+c13595;
assign A1595=(C1595>=0)?1:0;

ninexnine_unit ninexnine_unit_4240(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c105A5)
);

ninexnine_unit ninexnine_unit_4241(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c115A5)
);

ninexnine_unit ninexnine_unit_4242(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c125A5)
);

ninexnine_unit ninexnine_unit_4243(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c135A5)
);

assign C15A5=c105A5+c115A5+c125A5+c135A5;
assign A15A5=(C15A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4244(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c105B5)
);

ninexnine_unit ninexnine_unit_4245(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c115B5)
);

ninexnine_unit ninexnine_unit_4246(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c125B5)
);

ninexnine_unit ninexnine_unit_4247(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c135B5)
);

assign C15B5=c105B5+c115B5+c125B5+c135B5;
assign A15B5=(C15B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4248(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c105C5)
);

ninexnine_unit ninexnine_unit_4249(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c115C5)
);

ninexnine_unit ninexnine_unit_4250(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c125C5)
);

ninexnine_unit ninexnine_unit_4251(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c135C5)
);

assign C15C5=c105C5+c115C5+c125C5+c135C5;
assign A15C5=(C15C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4252(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c105D5)
);

ninexnine_unit ninexnine_unit_4253(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c115D5)
);

ninexnine_unit ninexnine_unit_4254(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c125D5)
);

ninexnine_unit ninexnine_unit_4255(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c135D5)
);

assign C15D5=c105D5+c115D5+c125D5+c135D5;
assign A15D5=(C15D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10605)
);

ninexnine_unit ninexnine_unit_4257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11605)
);

ninexnine_unit ninexnine_unit_4258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12605)
);

ninexnine_unit ninexnine_unit_4259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13605)
);

assign C1605=c10605+c11605+c12605+c13605;
assign A1605=(C1605>=0)?1:0;

ninexnine_unit ninexnine_unit_4260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10615)
);

ninexnine_unit ninexnine_unit_4261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11615)
);

ninexnine_unit ninexnine_unit_4262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12615)
);

ninexnine_unit ninexnine_unit_4263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13615)
);

assign C1615=c10615+c11615+c12615+c13615;
assign A1615=(C1615>=0)?1:0;

ninexnine_unit ninexnine_unit_4264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10625)
);

ninexnine_unit ninexnine_unit_4265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11625)
);

ninexnine_unit ninexnine_unit_4266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12625)
);

ninexnine_unit ninexnine_unit_4267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13625)
);

assign C1625=c10625+c11625+c12625+c13625;
assign A1625=(C1625>=0)?1:0;

ninexnine_unit ninexnine_unit_4268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10635)
);

ninexnine_unit ninexnine_unit_4269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11635)
);

ninexnine_unit ninexnine_unit_4270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12635)
);

ninexnine_unit ninexnine_unit_4271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13635)
);

assign C1635=c10635+c11635+c12635+c13635;
assign A1635=(C1635>=0)?1:0;

ninexnine_unit ninexnine_unit_4272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10645)
);

ninexnine_unit ninexnine_unit_4273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11645)
);

ninexnine_unit ninexnine_unit_4274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12645)
);

ninexnine_unit ninexnine_unit_4275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13645)
);

assign C1645=c10645+c11645+c12645+c13645;
assign A1645=(C1645>=0)?1:0;

ninexnine_unit ninexnine_unit_4276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10655)
);

ninexnine_unit ninexnine_unit_4277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11655)
);

ninexnine_unit ninexnine_unit_4278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12655)
);

ninexnine_unit ninexnine_unit_4279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13655)
);

assign C1655=c10655+c11655+c12655+c13655;
assign A1655=(C1655>=0)?1:0;

ninexnine_unit ninexnine_unit_4280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10665)
);

ninexnine_unit ninexnine_unit_4281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11665)
);

ninexnine_unit ninexnine_unit_4282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12665)
);

ninexnine_unit ninexnine_unit_4283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13665)
);

assign C1665=c10665+c11665+c12665+c13665;
assign A1665=(C1665>=0)?1:0;

ninexnine_unit ninexnine_unit_4284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10675)
);

ninexnine_unit ninexnine_unit_4285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11675)
);

ninexnine_unit ninexnine_unit_4286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12675)
);

ninexnine_unit ninexnine_unit_4287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13675)
);

assign C1675=c10675+c11675+c12675+c13675;
assign A1675=(C1675>=0)?1:0;

ninexnine_unit ninexnine_unit_4288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10685)
);

ninexnine_unit ninexnine_unit_4289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11685)
);

ninexnine_unit ninexnine_unit_4290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12685)
);

ninexnine_unit ninexnine_unit_4291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13685)
);

assign C1685=c10685+c11685+c12685+c13685;
assign A1685=(C1685>=0)?1:0;

ninexnine_unit ninexnine_unit_4292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10695)
);

ninexnine_unit ninexnine_unit_4293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11695)
);

ninexnine_unit ninexnine_unit_4294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12695)
);

ninexnine_unit ninexnine_unit_4295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13695)
);

assign C1695=c10695+c11695+c12695+c13695;
assign A1695=(C1695>=0)?1:0;

ninexnine_unit ninexnine_unit_4296(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c106A5)
);

ninexnine_unit ninexnine_unit_4297(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c116A5)
);

ninexnine_unit ninexnine_unit_4298(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c126A5)
);

ninexnine_unit ninexnine_unit_4299(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c136A5)
);

assign C16A5=c106A5+c116A5+c126A5+c136A5;
assign A16A5=(C16A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4300(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c106B5)
);

ninexnine_unit ninexnine_unit_4301(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c116B5)
);

ninexnine_unit ninexnine_unit_4302(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c126B5)
);

ninexnine_unit ninexnine_unit_4303(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c136B5)
);

assign C16B5=c106B5+c116B5+c126B5+c136B5;
assign A16B5=(C16B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4304(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c106C5)
);

ninexnine_unit ninexnine_unit_4305(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c116C5)
);

ninexnine_unit ninexnine_unit_4306(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c126C5)
);

ninexnine_unit ninexnine_unit_4307(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c136C5)
);

assign C16C5=c106C5+c116C5+c126C5+c136C5;
assign A16C5=(C16C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4308(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c106D5)
);

ninexnine_unit ninexnine_unit_4309(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c116D5)
);

ninexnine_unit ninexnine_unit_4310(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c126D5)
);

ninexnine_unit ninexnine_unit_4311(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c136D5)
);

assign C16D5=c106D5+c116D5+c126D5+c136D5;
assign A16D5=(C16D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10705)
);

ninexnine_unit ninexnine_unit_4313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11705)
);

ninexnine_unit ninexnine_unit_4314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12705)
);

ninexnine_unit ninexnine_unit_4315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13705)
);

assign C1705=c10705+c11705+c12705+c13705;
assign A1705=(C1705>=0)?1:0;

ninexnine_unit ninexnine_unit_4316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10715)
);

ninexnine_unit ninexnine_unit_4317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11715)
);

ninexnine_unit ninexnine_unit_4318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12715)
);

ninexnine_unit ninexnine_unit_4319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13715)
);

assign C1715=c10715+c11715+c12715+c13715;
assign A1715=(C1715>=0)?1:0;

ninexnine_unit ninexnine_unit_4320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10725)
);

ninexnine_unit ninexnine_unit_4321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11725)
);

ninexnine_unit ninexnine_unit_4322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12725)
);

ninexnine_unit ninexnine_unit_4323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13725)
);

assign C1725=c10725+c11725+c12725+c13725;
assign A1725=(C1725>=0)?1:0;

ninexnine_unit ninexnine_unit_4324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10735)
);

ninexnine_unit ninexnine_unit_4325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11735)
);

ninexnine_unit ninexnine_unit_4326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12735)
);

ninexnine_unit ninexnine_unit_4327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13735)
);

assign C1735=c10735+c11735+c12735+c13735;
assign A1735=(C1735>=0)?1:0;

ninexnine_unit ninexnine_unit_4328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10745)
);

ninexnine_unit ninexnine_unit_4329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11745)
);

ninexnine_unit ninexnine_unit_4330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12745)
);

ninexnine_unit ninexnine_unit_4331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13745)
);

assign C1745=c10745+c11745+c12745+c13745;
assign A1745=(C1745>=0)?1:0;

ninexnine_unit ninexnine_unit_4332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10755)
);

ninexnine_unit ninexnine_unit_4333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11755)
);

ninexnine_unit ninexnine_unit_4334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12755)
);

ninexnine_unit ninexnine_unit_4335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13755)
);

assign C1755=c10755+c11755+c12755+c13755;
assign A1755=(C1755>=0)?1:0;

ninexnine_unit ninexnine_unit_4336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10765)
);

ninexnine_unit ninexnine_unit_4337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11765)
);

ninexnine_unit ninexnine_unit_4338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12765)
);

ninexnine_unit ninexnine_unit_4339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13765)
);

assign C1765=c10765+c11765+c12765+c13765;
assign A1765=(C1765>=0)?1:0;

ninexnine_unit ninexnine_unit_4340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10775)
);

ninexnine_unit ninexnine_unit_4341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11775)
);

ninexnine_unit ninexnine_unit_4342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12775)
);

ninexnine_unit ninexnine_unit_4343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13775)
);

assign C1775=c10775+c11775+c12775+c13775;
assign A1775=(C1775>=0)?1:0;

ninexnine_unit ninexnine_unit_4344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10785)
);

ninexnine_unit ninexnine_unit_4345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11785)
);

ninexnine_unit ninexnine_unit_4346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12785)
);

ninexnine_unit ninexnine_unit_4347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13785)
);

assign C1785=c10785+c11785+c12785+c13785;
assign A1785=(C1785>=0)?1:0;

ninexnine_unit ninexnine_unit_4348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10795)
);

ninexnine_unit ninexnine_unit_4349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11795)
);

ninexnine_unit ninexnine_unit_4350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12795)
);

ninexnine_unit ninexnine_unit_4351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13795)
);

assign C1795=c10795+c11795+c12795+c13795;
assign A1795=(C1795>=0)?1:0;

ninexnine_unit ninexnine_unit_4352(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c107A5)
);

ninexnine_unit ninexnine_unit_4353(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c117A5)
);

ninexnine_unit ninexnine_unit_4354(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c127A5)
);

ninexnine_unit ninexnine_unit_4355(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c137A5)
);

assign C17A5=c107A5+c117A5+c127A5+c137A5;
assign A17A5=(C17A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4356(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c107B5)
);

ninexnine_unit ninexnine_unit_4357(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c117B5)
);

ninexnine_unit ninexnine_unit_4358(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c127B5)
);

ninexnine_unit ninexnine_unit_4359(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c137B5)
);

assign C17B5=c107B5+c117B5+c127B5+c137B5;
assign A17B5=(C17B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4360(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c107C5)
);

ninexnine_unit ninexnine_unit_4361(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c117C5)
);

ninexnine_unit ninexnine_unit_4362(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c127C5)
);

ninexnine_unit ninexnine_unit_4363(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c137C5)
);

assign C17C5=c107C5+c117C5+c127C5+c137C5;
assign A17C5=(C17C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4364(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c107D5)
);

ninexnine_unit ninexnine_unit_4365(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c117D5)
);

ninexnine_unit ninexnine_unit_4366(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c127D5)
);

ninexnine_unit ninexnine_unit_4367(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c137D5)
);

assign C17D5=c107D5+c117D5+c127D5+c137D5;
assign A17D5=(C17D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10805)
);

ninexnine_unit ninexnine_unit_4369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11805)
);

ninexnine_unit ninexnine_unit_4370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12805)
);

ninexnine_unit ninexnine_unit_4371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13805)
);

assign C1805=c10805+c11805+c12805+c13805;
assign A1805=(C1805>=0)?1:0;

ninexnine_unit ninexnine_unit_4372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10815)
);

ninexnine_unit ninexnine_unit_4373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11815)
);

ninexnine_unit ninexnine_unit_4374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12815)
);

ninexnine_unit ninexnine_unit_4375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13815)
);

assign C1815=c10815+c11815+c12815+c13815;
assign A1815=(C1815>=0)?1:0;

ninexnine_unit ninexnine_unit_4376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10825)
);

ninexnine_unit ninexnine_unit_4377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11825)
);

ninexnine_unit ninexnine_unit_4378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12825)
);

ninexnine_unit ninexnine_unit_4379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13825)
);

assign C1825=c10825+c11825+c12825+c13825;
assign A1825=(C1825>=0)?1:0;

ninexnine_unit ninexnine_unit_4380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10835)
);

ninexnine_unit ninexnine_unit_4381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11835)
);

ninexnine_unit ninexnine_unit_4382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12835)
);

ninexnine_unit ninexnine_unit_4383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13835)
);

assign C1835=c10835+c11835+c12835+c13835;
assign A1835=(C1835>=0)?1:0;

ninexnine_unit ninexnine_unit_4384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10845)
);

ninexnine_unit ninexnine_unit_4385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11845)
);

ninexnine_unit ninexnine_unit_4386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12845)
);

ninexnine_unit ninexnine_unit_4387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13845)
);

assign C1845=c10845+c11845+c12845+c13845;
assign A1845=(C1845>=0)?1:0;

ninexnine_unit ninexnine_unit_4388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10855)
);

ninexnine_unit ninexnine_unit_4389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11855)
);

ninexnine_unit ninexnine_unit_4390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12855)
);

ninexnine_unit ninexnine_unit_4391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13855)
);

assign C1855=c10855+c11855+c12855+c13855;
assign A1855=(C1855>=0)?1:0;

ninexnine_unit ninexnine_unit_4392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10865)
);

ninexnine_unit ninexnine_unit_4393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11865)
);

ninexnine_unit ninexnine_unit_4394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12865)
);

ninexnine_unit ninexnine_unit_4395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13865)
);

assign C1865=c10865+c11865+c12865+c13865;
assign A1865=(C1865>=0)?1:0;

ninexnine_unit ninexnine_unit_4396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10875)
);

ninexnine_unit ninexnine_unit_4397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11875)
);

ninexnine_unit ninexnine_unit_4398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12875)
);

ninexnine_unit ninexnine_unit_4399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13875)
);

assign C1875=c10875+c11875+c12875+c13875;
assign A1875=(C1875>=0)?1:0;

ninexnine_unit ninexnine_unit_4400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10885)
);

ninexnine_unit ninexnine_unit_4401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11885)
);

ninexnine_unit ninexnine_unit_4402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12885)
);

ninexnine_unit ninexnine_unit_4403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13885)
);

assign C1885=c10885+c11885+c12885+c13885;
assign A1885=(C1885>=0)?1:0;

ninexnine_unit ninexnine_unit_4404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10895)
);

ninexnine_unit ninexnine_unit_4405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11895)
);

ninexnine_unit ninexnine_unit_4406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12895)
);

ninexnine_unit ninexnine_unit_4407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13895)
);

assign C1895=c10895+c11895+c12895+c13895;
assign A1895=(C1895>=0)?1:0;

ninexnine_unit ninexnine_unit_4408(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c108A5)
);

ninexnine_unit ninexnine_unit_4409(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c118A5)
);

ninexnine_unit ninexnine_unit_4410(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c128A5)
);

ninexnine_unit ninexnine_unit_4411(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c138A5)
);

assign C18A5=c108A5+c118A5+c128A5+c138A5;
assign A18A5=(C18A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4412(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c108B5)
);

ninexnine_unit ninexnine_unit_4413(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c118B5)
);

ninexnine_unit ninexnine_unit_4414(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c128B5)
);

ninexnine_unit ninexnine_unit_4415(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c138B5)
);

assign C18B5=c108B5+c118B5+c128B5+c138B5;
assign A18B5=(C18B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4416(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c108C5)
);

ninexnine_unit ninexnine_unit_4417(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c118C5)
);

ninexnine_unit ninexnine_unit_4418(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c128C5)
);

ninexnine_unit ninexnine_unit_4419(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c138C5)
);

assign C18C5=c108C5+c118C5+c128C5+c138C5;
assign A18C5=(C18C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4420(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c108D5)
);

ninexnine_unit ninexnine_unit_4421(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c118D5)
);

ninexnine_unit ninexnine_unit_4422(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c128D5)
);

ninexnine_unit ninexnine_unit_4423(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c138D5)
);

assign C18D5=c108D5+c118D5+c128D5+c138D5;
assign A18D5=(C18D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10905)
);

ninexnine_unit ninexnine_unit_4425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11905)
);

ninexnine_unit ninexnine_unit_4426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12905)
);

ninexnine_unit ninexnine_unit_4427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13905)
);

assign C1905=c10905+c11905+c12905+c13905;
assign A1905=(C1905>=0)?1:0;

ninexnine_unit ninexnine_unit_4428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10915)
);

ninexnine_unit ninexnine_unit_4429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11915)
);

ninexnine_unit ninexnine_unit_4430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12915)
);

ninexnine_unit ninexnine_unit_4431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13915)
);

assign C1915=c10915+c11915+c12915+c13915;
assign A1915=(C1915>=0)?1:0;

ninexnine_unit ninexnine_unit_4432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10925)
);

ninexnine_unit ninexnine_unit_4433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11925)
);

ninexnine_unit ninexnine_unit_4434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12925)
);

ninexnine_unit ninexnine_unit_4435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13925)
);

assign C1925=c10925+c11925+c12925+c13925;
assign A1925=(C1925>=0)?1:0;

ninexnine_unit ninexnine_unit_4436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10935)
);

ninexnine_unit ninexnine_unit_4437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11935)
);

ninexnine_unit ninexnine_unit_4438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12935)
);

ninexnine_unit ninexnine_unit_4439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13935)
);

assign C1935=c10935+c11935+c12935+c13935;
assign A1935=(C1935>=0)?1:0;

ninexnine_unit ninexnine_unit_4440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10945)
);

ninexnine_unit ninexnine_unit_4441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11945)
);

ninexnine_unit ninexnine_unit_4442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12945)
);

ninexnine_unit ninexnine_unit_4443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13945)
);

assign C1945=c10945+c11945+c12945+c13945;
assign A1945=(C1945>=0)?1:0;

ninexnine_unit ninexnine_unit_4444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10955)
);

ninexnine_unit ninexnine_unit_4445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11955)
);

ninexnine_unit ninexnine_unit_4446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12955)
);

ninexnine_unit ninexnine_unit_4447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13955)
);

assign C1955=c10955+c11955+c12955+c13955;
assign A1955=(C1955>=0)?1:0;

ninexnine_unit ninexnine_unit_4448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10965)
);

ninexnine_unit ninexnine_unit_4449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11965)
);

ninexnine_unit ninexnine_unit_4450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12965)
);

ninexnine_unit ninexnine_unit_4451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13965)
);

assign C1965=c10965+c11965+c12965+c13965;
assign A1965=(C1965>=0)?1:0;

ninexnine_unit ninexnine_unit_4452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10975)
);

ninexnine_unit ninexnine_unit_4453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11975)
);

ninexnine_unit ninexnine_unit_4454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12975)
);

ninexnine_unit ninexnine_unit_4455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13975)
);

assign C1975=c10975+c11975+c12975+c13975;
assign A1975=(C1975>=0)?1:0;

ninexnine_unit ninexnine_unit_4456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10985)
);

ninexnine_unit ninexnine_unit_4457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11985)
);

ninexnine_unit ninexnine_unit_4458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12985)
);

ninexnine_unit ninexnine_unit_4459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13985)
);

assign C1985=c10985+c11985+c12985+c13985;
assign A1985=(C1985>=0)?1:0;

ninexnine_unit ninexnine_unit_4460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10995)
);

ninexnine_unit ninexnine_unit_4461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11995)
);

ninexnine_unit ninexnine_unit_4462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12995)
);

ninexnine_unit ninexnine_unit_4463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13995)
);

assign C1995=c10995+c11995+c12995+c13995;
assign A1995=(C1995>=0)?1:0;

ninexnine_unit ninexnine_unit_4464(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c109A5)
);

ninexnine_unit ninexnine_unit_4465(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c119A5)
);

ninexnine_unit ninexnine_unit_4466(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c129A5)
);

ninexnine_unit ninexnine_unit_4467(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c139A5)
);

assign C19A5=c109A5+c119A5+c129A5+c139A5;
assign A19A5=(C19A5>=0)?1:0;

ninexnine_unit ninexnine_unit_4468(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c109B5)
);

ninexnine_unit ninexnine_unit_4469(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c119B5)
);

ninexnine_unit ninexnine_unit_4470(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c129B5)
);

ninexnine_unit ninexnine_unit_4471(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c139B5)
);

assign C19B5=c109B5+c119B5+c129B5+c139B5;
assign A19B5=(C19B5>=0)?1:0;

ninexnine_unit ninexnine_unit_4472(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c109C5)
);

ninexnine_unit ninexnine_unit_4473(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c119C5)
);

ninexnine_unit ninexnine_unit_4474(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c129C5)
);

ninexnine_unit ninexnine_unit_4475(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c139C5)
);

assign C19C5=c109C5+c119C5+c129C5+c139C5;
assign A19C5=(C19C5>=0)?1:0;

ninexnine_unit ninexnine_unit_4476(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c109D5)
);

ninexnine_unit ninexnine_unit_4477(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c119D5)
);

ninexnine_unit ninexnine_unit_4478(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c129D5)
);

ninexnine_unit ninexnine_unit_4479(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c139D5)
);

assign C19D5=c109D5+c119D5+c129D5+c139D5;
assign A19D5=(C19D5>=0)?1:0;

ninexnine_unit ninexnine_unit_4480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A05)
);

ninexnine_unit ninexnine_unit_4481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A05)
);

ninexnine_unit ninexnine_unit_4482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A05)
);

ninexnine_unit ninexnine_unit_4483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A05)
);

assign C1A05=c10A05+c11A05+c12A05+c13A05;
assign A1A05=(C1A05>=0)?1:0;

ninexnine_unit ninexnine_unit_4484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A15)
);

ninexnine_unit ninexnine_unit_4485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A15)
);

ninexnine_unit ninexnine_unit_4486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A15)
);

ninexnine_unit ninexnine_unit_4487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A15)
);

assign C1A15=c10A15+c11A15+c12A15+c13A15;
assign A1A15=(C1A15>=0)?1:0;

ninexnine_unit ninexnine_unit_4488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A25)
);

ninexnine_unit ninexnine_unit_4489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A25)
);

ninexnine_unit ninexnine_unit_4490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A25)
);

ninexnine_unit ninexnine_unit_4491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A25)
);

assign C1A25=c10A25+c11A25+c12A25+c13A25;
assign A1A25=(C1A25>=0)?1:0;

ninexnine_unit ninexnine_unit_4492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A35)
);

ninexnine_unit ninexnine_unit_4493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A35)
);

ninexnine_unit ninexnine_unit_4494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A35)
);

ninexnine_unit ninexnine_unit_4495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A35)
);

assign C1A35=c10A35+c11A35+c12A35+c13A35;
assign A1A35=(C1A35>=0)?1:0;

ninexnine_unit ninexnine_unit_4496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A45)
);

ninexnine_unit ninexnine_unit_4497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A45)
);

ninexnine_unit ninexnine_unit_4498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A45)
);

ninexnine_unit ninexnine_unit_4499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A45)
);

assign C1A45=c10A45+c11A45+c12A45+c13A45;
assign A1A45=(C1A45>=0)?1:0;

ninexnine_unit ninexnine_unit_4500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A55)
);

ninexnine_unit ninexnine_unit_4501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A55)
);

ninexnine_unit ninexnine_unit_4502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A55)
);

ninexnine_unit ninexnine_unit_4503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A55)
);

assign C1A55=c10A55+c11A55+c12A55+c13A55;
assign A1A55=(C1A55>=0)?1:0;

ninexnine_unit ninexnine_unit_4504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A65)
);

ninexnine_unit ninexnine_unit_4505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A65)
);

ninexnine_unit ninexnine_unit_4506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A65)
);

ninexnine_unit ninexnine_unit_4507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A65)
);

assign C1A65=c10A65+c11A65+c12A65+c13A65;
assign A1A65=(C1A65>=0)?1:0;

ninexnine_unit ninexnine_unit_4508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A75)
);

ninexnine_unit ninexnine_unit_4509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A75)
);

ninexnine_unit ninexnine_unit_4510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A75)
);

ninexnine_unit ninexnine_unit_4511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A75)
);

assign C1A75=c10A75+c11A75+c12A75+c13A75;
assign A1A75=(C1A75>=0)?1:0;

ninexnine_unit ninexnine_unit_4512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A85)
);

ninexnine_unit ninexnine_unit_4513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A85)
);

ninexnine_unit ninexnine_unit_4514(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A85)
);

ninexnine_unit ninexnine_unit_4515(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A85)
);

assign C1A85=c10A85+c11A85+c12A85+c13A85;
assign A1A85=(C1A85>=0)?1:0;

ninexnine_unit ninexnine_unit_4516(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10A95)
);

ninexnine_unit ninexnine_unit_4517(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11A95)
);

ninexnine_unit ninexnine_unit_4518(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12A95)
);

ninexnine_unit ninexnine_unit_4519(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13A95)
);

assign C1A95=c10A95+c11A95+c12A95+c13A95;
assign A1A95=(C1A95>=0)?1:0;

ninexnine_unit ninexnine_unit_4520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10AA5)
);

ninexnine_unit ninexnine_unit_4521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11AA5)
);

ninexnine_unit ninexnine_unit_4522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12AA5)
);

ninexnine_unit ninexnine_unit_4523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13AA5)
);

assign C1AA5=c10AA5+c11AA5+c12AA5+c13AA5;
assign A1AA5=(C1AA5>=0)?1:0;

ninexnine_unit ninexnine_unit_4524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10AB5)
);

ninexnine_unit ninexnine_unit_4525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11AB5)
);

ninexnine_unit ninexnine_unit_4526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12AB5)
);

ninexnine_unit ninexnine_unit_4527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13AB5)
);

assign C1AB5=c10AB5+c11AB5+c12AB5+c13AB5;
assign A1AB5=(C1AB5>=0)?1:0;

ninexnine_unit ninexnine_unit_4528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10AC5)
);

ninexnine_unit ninexnine_unit_4529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11AC5)
);

ninexnine_unit ninexnine_unit_4530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12AC5)
);

ninexnine_unit ninexnine_unit_4531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13AC5)
);

assign C1AC5=c10AC5+c11AC5+c12AC5+c13AC5;
assign A1AC5=(C1AC5>=0)?1:0;

ninexnine_unit ninexnine_unit_4532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10AD5)
);

ninexnine_unit ninexnine_unit_4533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11AD5)
);

ninexnine_unit ninexnine_unit_4534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12AD5)
);

ninexnine_unit ninexnine_unit_4535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13AD5)
);

assign C1AD5=c10AD5+c11AD5+c12AD5+c13AD5;
assign A1AD5=(C1AD5>=0)?1:0;

ninexnine_unit ninexnine_unit_4536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B05)
);

ninexnine_unit ninexnine_unit_4537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B05)
);

ninexnine_unit ninexnine_unit_4538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B05)
);

ninexnine_unit ninexnine_unit_4539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B05)
);

assign C1B05=c10B05+c11B05+c12B05+c13B05;
assign A1B05=(C1B05>=0)?1:0;

ninexnine_unit ninexnine_unit_4540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B15)
);

ninexnine_unit ninexnine_unit_4541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B15)
);

ninexnine_unit ninexnine_unit_4542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B15)
);

ninexnine_unit ninexnine_unit_4543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B15)
);

assign C1B15=c10B15+c11B15+c12B15+c13B15;
assign A1B15=(C1B15>=0)?1:0;

ninexnine_unit ninexnine_unit_4544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B25)
);

ninexnine_unit ninexnine_unit_4545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B25)
);

ninexnine_unit ninexnine_unit_4546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B25)
);

ninexnine_unit ninexnine_unit_4547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B25)
);

assign C1B25=c10B25+c11B25+c12B25+c13B25;
assign A1B25=(C1B25>=0)?1:0;

ninexnine_unit ninexnine_unit_4548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B35)
);

ninexnine_unit ninexnine_unit_4549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B35)
);

ninexnine_unit ninexnine_unit_4550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B35)
);

ninexnine_unit ninexnine_unit_4551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B35)
);

assign C1B35=c10B35+c11B35+c12B35+c13B35;
assign A1B35=(C1B35>=0)?1:0;

ninexnine_unit ninexnine_unit_4552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B45)
);

ninexnine_unit ninexnine_unit_4553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B45)
);

ninexnine_unit ninexnine_unit_4554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B45)
);

ninexnine_unit ninexnine_unit_4555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B45)
);

assign C1B45=c10B45+c11B45+c12B45+c13B45;
assign A1B45=(C1B45>=0)?1:0;

ninexnine_unit ninexnine_unit_4556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B55)
);

ninexnine_unit ninexnine_unit_4557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B55)
);

ninexnine_unit ninexnine_unit_4558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B55)
);

ninexnine_unit ninexnine_unit_4559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B55)
);

assign C1B55=c10B55+c11B55+c12B55+c13B55;
assign A1B55=(C1B55>=0)?1:0;

ninexnine_unit ninexnine_unit_4560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B65)
);

ninexnine_unit ninexnine_unit_4561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B65)
);

ninexnine_unit ninexnine_unit_4562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B65)
);

ninexnine_unit ninexnine_unit_4563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B65)
);

assign C1B65=c10B65+c11B65+c12B65+c13B65;
assign A1B65=(C1B65>=0)?1:0;

ninexnine_unit ninexnine_unit_4564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B75)
);

ninexnine_unit ninexnine_unit_4565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B75)
);

ninexnine_unit ninexnine_unit_4566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B75)
);

ninexnine_unit ninexnine_unit_4567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B75)
);

assign C1B75=c10B75+c11B75+c12B75+c13B75;
assign A1B75=(C1B75>=0)?1:0;

ninexnine_unit ninexnine_unit_4568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B85)
);

ninexnine_unit ninexnine_unit_4569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B85)
);

ninexnine_unit ninexnine_unit_4570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B85)
);

ninexnine_unit ninexnine_unit_4571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B85)
);

assign C1B85=c10B85+c11B85+c12B85+c13B85;
assign A1B85=(C1B85>=0)?1:0;

ninexnine_unit ninexnine_unit_4572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10B95)
);

ninexnine_unit ninexnine_unit_4573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11B95)
);

ninexnine_unit ninexnine_unit_4574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12B95)
);

ninexnine_unit ninexnine_unit_4575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13B95)
);

assign C1B95=c10B95+c11B95+c12B95+c13B95;
assign A1B95=(C1B95>=0)?1:0;

ninexnine_unit ninexnine_unit_4576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10BA5)
);

ninexnine_unit ninexnine_unit_4577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11BA5)
);

ninexnine_unit ninexnine_unit_4578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12BA5)
);

ninexnine_unit ninexnine_unit_4579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13BA5)
);

assign C1BA5=c10BA5+c11BA5+c12BA5+c13BA5;
assign A1BA5=(C1BA5>=0)?1:0;

ninexnine_unit ninexnine_unit_4580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10BB5)
);

ninexnine_unit ninexnine_unit_4581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11BB5)
);

ninexnine_unit ninexnine_unit_4582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12BB5)
);

ninexnine_unit ninexnine_unit_4583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13BB5)
);

assign C1BB5=c10BB5+c11BB5+c12BB5+c13BB5;
assign A1BB5=(C1BB5>=0)?1:0;

ninexnine_unit ninexnine_unit_4584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10BC5)
);

ninexnine_unit ninexnine_unit_4585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11BC5)
);

ninexnine_unit ninexnine_unit_4586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12BC5)
);

ninexnine_unit ninexnine_unit_4587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13BC5)
);

assign C1BC5=c10BC5+c11BC5+c12BC5+c13BC5;
assign A1BC5=(C1BC5>=0)?1:0;

ninexnine_unit ninexnine_unit_4588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10BD5)
);

ninexnine_unit ninexnine_unit_4589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11BD5)
);

ninexnine_unit ninexnine_unit_4590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12BD5)
);

ninexnine_unit ninexnine_unit_4591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13BD5)
);

assign C1BD5=c10BD5+c11BD5+c12BD5+c13BD5;
assign A1BD5=(C1BD5>=0)?1:0;

ninexnine_unit ninexnine_unit_4592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C05)
);

ninexnine_unit ninexnine_unit_4593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C05)
);

ninexnine_unit ninexnine_unit_4594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C05)
);

ninexnine_unit ninexnine_unit_4595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C05)
);

assign C1C05=c10C05+c11C05+c12C05+c13C05;
assign A1C05=(C1C05>=0)?1:0;

ninexnine_unit ninexnine_unit_4596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C15)
);

ninexnine_unit ninexnine_unit_4597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C15)
);

ninexnine_unit ninexnine_unit_4598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C15)
);

ninexnine_unit ninexnine_unit_4599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C15)
);

assign C1C15=c10C15+c11C15+c12C15+c13C15;
assign A1C15=(C1C15>=0)?1:0;

ninexnine_unit ninexnine_unit_4600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C25)
);

ninexnine_unit ninexnine_unit_4601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C25)
);

ninexnine_unit ninexnine_unit_4602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C25)
);

ninexnine_unit ninexnine_unit_4603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C25)
);

assign C1C25=c10C25+c11C25+c12C25+c13C25;
assign A1C25=(C1C25>=0)?1:0;

ninexnine_unit ninexnine_unit_4604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C35)
);

ninexnine_unit ninexnine_unit_4605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C35)
);

ninexnine_unit ninexnine_unit_4606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C35)
);

ninexnine_unit ninexnine_unit_4607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C35)
);

assign C1C35=c10C35+c11C35+c12C35+c13C35;
assign A1C35=(C1C35>=0)?1:0;

ninexnine_unit ninexnine_unit_4608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C45)
);

ninexnine_unit ninexnine_unit_4609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C45)
);

ninexnine_unit ninexnine_unit_4610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C45)
);

ninexnine_unit ninexnine_unit_4611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C45)
);

assign C1C45=c10C45+c11C45+c12C45+c13C45;
assign A1C45=(C1C45>=0)?1:0;

ninexnine_unit ninexnine_unit_4612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C55)
);

ninexnine_unit ninexnine_unit_4613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C55)
);

ninexnine_unit ninexnine_unit_4614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C55)
);

ninexnine_unit ninexnine_unit_4615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C55)
);

assign C1C55=c10C55+c11C55+c12C55+c13C55;
assign A1C55=(C1C55>=0)?1:0;

ninexnine_unit ninexnine_unit_4616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C65)
);

ninexnine_unit ninexnine_unit_4617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C65)
);

ninexnine_unit ninexnine_unit_4618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C65)
);

ninexnine_unit ninexnine_unit_4619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C65)
);

assign C1C65=c10C65+c11C65+c12C65+c13C65;
assign A1C65=(C1C65>=0)?1:0;

ninexnine_unit ninexnine_unit_4620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C75)
);

ninexnine_unit ninexnine_unit_4621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C75)
);

ninexnine_unit ninexnine_unit_4622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C75)
);

ninexnine_unit ninexnine_unit_4623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C75)
);

assign C1C75=c10C75+c11C75+c12C75+c13C75;
assign A1C75=(C1C75>=0)?1:0;

ninexnine_unit ninexnine_unit_4624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C85)
);

ninexnine_unit ninexnine_unit_4625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C85)
);

ninexnine_unit ninexnine_unit_4626(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C85)
);

ninexnine_unit ninexnine_unit_4627(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C85)
);

assign C1C85=c10C85+c11C85+c12C85+c13C85;
assign A1C85=(C1C85>=0)?1:0;

ninexnine_unit ninexnine_unit_4628(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10C95)
);

ninexnine_unit ninexnine_unit_4629(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11C95)
);

ninexnine_unit ninexnine_unit_4630(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12C95)
);

ninexnine_unit ninexnine_unit_4631(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13C95)
);

assign C1C95=c10C95+c11C95+c12C95+c13C95;
assign A1C95=(C1C95>=0)?1:0;

ninexnine_unit ninexnine_unit_4632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10CA5)
);

ninexnine_unit ninexnine_unit_4633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11CA5)
);

ninexnine_unit ninexnine_unit_4634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12CA5)
);

ninexnine_unit ninexnine_unit_4635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13CA5)
);

assign C1CA5=c10CA5+c11CA5+c12CA5+c13CA5;
assign A1CA5=(C1CA5>=0)?1:0;

ninexnine_unit ninexnine_unit_4636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10CB5)
);

ninexnine_unit ninexnine_unit_4637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11CB5)
);

ninexnine_unit ninexnine_unit_4638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12CB5)
);

ninexnine_unit ninexnine_unit_4639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13CB5)
);

assign C1CB5=c10CB5+c11CB5+c12CB5+c13CB5;
assign A1CB5=(C1CB5>=0)?1:0;

ninexnine_unit ninexnine_unit_4640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10CC5)
);

ninexnine_unit ninexnine_unit_4641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11CC5)
);

ninexnine_unit ninexnine_unit_4642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12CC5)
);

ninexnine_unit ninexnine_unit_4643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13CC5)
);

assign C1CC5=c10CC5+c11CC5+c12CC5+c13CC5;
assign A1CC5=(C1CC5>=0)?1:0;

ninexnine_unit ninexnine_unit_4644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10CD5)
);

ninexnine_unit ninexnine_unit_4645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11CD5)
);

ninexnine_unit ninexnine_unit_4646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12CD5)
);

ninexnine_unit ninexnine_unit_4647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13CD5)
);

assign C1CD5=c10CD5+c11CD5+c12CD5+c13CD5;
assign A1CD5=(C1CD5>=0)?1:0;

ninexnine_unit ninexnine_unit_4648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D05)
);

ninexnine_unit ninexnine_unit_4649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D05)
);

ninexnine_unit ninexnine_unit_4650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D05)
);

ninexnine_unit ninexnine_unit_4651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D05)
);

assign C1D05=c10D05+c11D05+c12D05+c13D05;
assign A1D05=(C1D05>=0)?1:0;

ninexnine_unit ninexnine_unit_4652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D15)
);

ninexnine_unit ninexnine_unit_4653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D15)
);

ninexnine_unit ninexnine_unit_4654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D15)
);

ninexnine_unit ninexnine_unit_4655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D15)
);

assign C1D15=c10D15+c11D15+c12D15+c13D15;
assign A1D15=(C1D15>=0)?1:0;

ninexnine_unit ninexnine_unit_4656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D25)
);

ninexnine_unit ninexnine_unit_4657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D25)
);

ninexnine_unit ninexnine_unit_4658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D25)
);

ninexnine_unit ninexnine_unit_4659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D25)
);

assign C1D25=c10D25+c11D25+c12D25+c13D25;
assign A1D25=(C1D25>=0)?1:0;

ninexnine_unit ninexnine_unit_4660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D35)
);

ninexnine_unit ninexnine_unit_4661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D35)
);

ninexnine_unit ninexnine_unit_4662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D35)
);

ninexnine_unit ninexnine_unit_4663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D35)
);

assign C1D35=c10D35+c11D35+c12D35+c13D35;
assign A1D35=(C1D35>=0)?1:0;

ninexnine_unit ninexnine_unit_4664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D45)
);

ninexnine_unit ninexnine_unit_4665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D45)
);

ninexnine_unit ninexnine_unit_4666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D45)
);

ninexnine_unit ninexnine_unit_4667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D45)
);

assign C1D45=c10D45+c11D45+c12D45+c13D45;
assign A1D45=(C1D45>=0)?1:0;

ninexnine_unit ninexnine_unit_4668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D55)
);

ninexnine_unit ninexnine_unit_4669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D55)
);

ninexnine_unit ninexnine_unit_4670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D55)
);

ninexnine_unit ninexnine_unit_4671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D55)
);

assign C1D55=c10D55+c11D55+c12D55+c13D55;
assign A1D55=(C1D55>=0)?1:0;

ninexnine_unit ninexnine_unit_4672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D65)
);

ninexnine_unit ninexnine_unit_4673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D65)
);

ninexnine_unit ninexnine_unit_4674(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D65)
);

ninexnine_unit ninexnine_unit_4675(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D65)
);

assign C1D65=c10D65+c11D65+c12D65+c13D65;
assign A1D65=(C1D65>=0)?1:0;

ninexnine_unit ninexnine_unit_4676(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D75)
);

ninexnine_unit ninexnine_unit_4677(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D75)
);

ninexnine_unit ninexnine_unit_4678(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D75)
);

ninexnine_unit ninexnine_unit_4679(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D75)
);

assign C1D75=c10D75+c11D75+c12D75+c13D75;
assign A1D75=(C1D75>=0)?1:0;

ninexnine_unit ninexnine_unit_4680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D85)
);

ninexnine_unit ninexnine_unit_4681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D85)
);

ninexnine_unit ninexnine_unit_4682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D85)
);

ninexnine_unit ninexnine_unit_4683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D85)
);

assign C1D85=c10D85+c11D85+c12D85+c13D85;
assign A1D85=(C1D85>=0)?1:0;

ninexnine_unit ninexnine_unit_4684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10D95)
);

ninexnine_unit ninexnine_unit_4685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11D95)
);

ninexnine_unit ninexnine_unit_4686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12D95)
);

ninexnine_unit ninexnine_unit_4687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13D95)
);

assign C1D95=c10D95+c11D95+c12D95+c13D95;
assign A1D95=(C1D95>=0)?1:0;

ninexnine_unit ninexnine_unit_4688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10DA5)
);

ninexnine_unit ninexnine_unit_4689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11DA5)
);

ninexnine_unit ninexnine_unit_4690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12DA5)
);

ninexnine_unit ninexnine_unit_4691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13DA5)
);

assign C1DA5=c10DA5+c11DA5+c12DA5+c13DA5;
assign A1DA5=(C1DA5>=0)?1:0;

ninexnine_unit ninexnine_unit_4692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10DB5)
);

ninexnine_unit ninexnine_unit_4693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11DB5)
);

ninexnine_unit ninexnine_unit_4694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12DB5)
);

ninexnine_unit ninexnine_unit_4695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13DB5)
);

assign C1DB5=c10DB5+c11DB5+c12DB5+c13DB5;
assign A1DB5=(C1DB5>=0)?1:0;

ninexnine_unit ninexnine_unit_4696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10DC5)
);

ninexnine_unit ninexnine_unit_4697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11DC5)
);

ninexnine_unit ninexnine_unit_4698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12DC5)
);

ninexnine_unit ninexnine_unit_4699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13DC5)
);

assign C1DC5=c10DC5+c11DC5+c12DC5+c13DC5;
assign A1DC5=(C1DC5>=0)?1:0;

ninexnine_unit ninexnine_unit_4700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10DD5)
);

ninexnine_unit ninexnine_unit_4701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11DD5)
);

ninexnine_unit ninexnine_unit_4702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12DD5)
);

ninexnine_unit ninexnine_unit_4703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13DD5)
);

assign C1DD5=c10DD5+c11DD5+c12DD5+c13DD5;
assign A1DD5=(C1DD5>=0)?1:0;

ninexnine_unit ninexnine_unit_4704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10006)
);

ninexnine_unit ninexnine_unit_4705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11006)
);

ninexnine_unit ninexnine_unit_4706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12006)
);

ninexnine_unit ninexnine_unit_4707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13006)
);

assign C1006=c10006+c11006+c12006+c13006;
assign A1006=(C1006>=0)?1:0;

ninexnine_unit ninexnine_unit_4708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10016)
);

ninexnine_unit ninexnine_unit_4709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11016)
);

ninexnine_unit ninexnine_unit_4710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12016)
);

ninexnine_unit ninexnine_unit_4711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13016)
);

assign C1016=c10016+c11016+c12016+c13016;
assign A1016=(C1016>=0)?1:0;

ninexnine_unit ninexnine_unit_4712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10026)
);

ninexnine_unit ninexnine_unit_4713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11026)
);

ninexnine_unit ninexnine_unit_4714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12026)
);

ninexnine_unit ninexnine_unit_4715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13026)
);

assign C1026=c10026+c11026+c12026+c13026;
assign A1026=(C1026>=0)?1:0;

ninexnine_unit ninexnine_unit_4716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10036)
);

ninexnine_unit ninexnine_unit_4717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11036)
);

ninexnine_unit ninexnine_unit_4718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12036)
);

ninexnine_unit ninexnine_unit_4719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13036)
);

assign C1036=c10036+c11036+c12036+c13036;
assign A1036=(C1036>=0)?1:0;

ninexnine_unit ninexnine_unit_4720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10046)
);

ninexnine_unit ninexnine_unit_4721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11046)
);

ninexnine_unit ninexnine_unit_4722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12046)
);

ninexnine_unit ninexnine_unit_4723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13046)
);

assign C1046=c10046+c11046+c12046+c13046;
assign A1046=(C1046>=0)?1:0;

ninexnine_unit ninexnine_unit_4724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10056)
);

ninexnine_unit ninexnine_unit_4725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11056)
);

ninexnine_unit ninexnine_unit_4726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12056)
);

ninexnine_unit ninexnine_unit_4727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13056)
);

assign C1056=c10056+c11056+c12056+c13056;
assign A1056=(C1056>=0)?1:0;

ninexnine_unit ninexnine_unit_4728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10066)
);

ninexnine_unit ninexnine_unit_4729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11066)
);

ninexnine_unit ninexnine_unit_4730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12066)
);

ninexnine_unit ninexnine_unit_4731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13066)
);

assign C1066=c10066+c11066+c12066+c13066;
assign A1066=(C1066>=0)?1:0;

ninexnine_unit ninexnine_unit_4732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10076)
);

ninexnine_unit ninexnine_unit_4733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11076)
);

ninexnine_unit ninexnine_unit_4734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12076)
);

ninexnine_unit ninexnine_unit_4735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13076)
);

assign C1076=c10076+c11076+c12076+c13076;
assign A1076=(C1076>=0)?1:0;

ninexnine_unit ninexnine_unit_4736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10086)
);

ninexnine_unit ninexnine_unit_4737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11086)
);

ninexnine_unit ninexnine_unit_4738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12086)
);

ninexnine_unit ninexnine_unit_4739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13086)
);

assign C1086=c10086+c11086+c12086+c13086;
assign A1086=(C1086>=0)?1:0;

ninexnine_unit ninexnine_unit_4740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10096)
);

ninexnine_unit ninexnine_unit_4741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11096)
);

ninexnine_unit ninexnine_unit_4742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12096)
);

ninexnine_unit ninexnine_unit_4743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13096)
);

assign C1096=c10096+c11096+c12096+c13096;
assign A1096=(C1096>=0)?1:0;

ninexnine_unit ninexnine_unit_4744(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c100A6)
);

ninexnine_unit ninexnine_unit_4745(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c110A6)
);

ninexnine_unit ninexnine_unit_4746(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c120A6)
);

ninexnine_unit ninexnine_unit_4747(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c130A6)
);

assign C10A6=c100A6+c110A6+c120A6+c130A6;
assign A10A6=(C10A6>=0)?1:0;

ninexnine_unit ninexnine_unit_4748(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c100B6)
);

ninexnine_unit ninexnine_unit_4749(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c110B6)
);

ninexnine_unit ninexnine_unit_4750(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c120B6)
);

ninexnine_unit ninexnine_unit_4751(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c130B6)
);

assign C10B6=c100B6+c110B6+c120B6+c130B6;
assign A10B6=(C10B6>=0)?1:0;

ninexnine_unit ninexnine_unit_4752(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c100C6)
);

ninexnine_unit ninexnine_unit_4753(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c110C6)
);

ninexnine_unit ninexnine_unit_4754(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c120C6)
);

ninexnine_unit ninexnine_unit_4755(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c130C6)
);

assign C10C6=c100C6+c110C6+c120C6+c130C6;
assign A10C6=(C10C6>=0)?1:0;

ninexnine_unit ninexnine_unit_4756(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c100D6)
);

ninexnine_unit ninexnine_unit_4757(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c110D6)
);

ninexnine_unit ninexnine_unit_4758(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c120D6)
);

ninexnine_unit ninexnine_unit_4759(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c130D6)
);

assign C10D6=c100D6+c110D6+c120D6+c130D6;
assign A10D6=(C10D6>=0)?1:0;

ninexnine_unit ninexnine_unit_4760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10106)
);

ninexnine_unit ninexnine_unit_4761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11106)
);

ninexnine_unit ninexnine_unit_4762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12106)
);

ninexnine_unit ninexnine_unit_4763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13106)
);

assign C1106=c10106+c11106+c12106+c13106;
assign A1106=(C1106>=0)?1:0;

ninexnine_unit ninexnine_unit_4764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10116)
);

ninexnine_unit ninexnine_unit_4765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11116)
);

ninexnine_unit ninexnine_unit_4766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12116)
);

ninexnine_unit ninexnine_unit_4767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13116)
);

assign C1116=c10116+c11116+c12116+c13116;
assign A1116=(C1116>=0)?1:0;

ninexnine_unit ninexnine_unit_4768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10126)
);

ninexnine_unit ninexnine_unit_4769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11126)
);

ninexnine_unit ninexnine_unit_4770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12126)
);

ninexnine_unit ninexnine_unit_4771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13126)
);

assign C1126=c10126+c11126+c12126+c13126;
assign A1126=(C1126>=0)?1:0;

ninexnine_unit ninexnine_unit_4772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10136)
);

ninexnine_unit ninexnine_unit_4773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11136)
);

ninexnine_unit ninexnine_unit_4774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12136)
);

ninexnine_unit ninexnine_unit_4775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13136)
);

assign C1136=c10136+c11136+c12136+c13136;
assign A1136=(C1136>=0)?1:0;

ninexnine_unit ninexnine_unit_4776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10146)
);

ninexnine_unit ninexnine_unit_4777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11146)
);

ninexnine_unit ninexnine_unit_4778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12146)
);

ninexnine_unit ninexnine_unit_4779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13146)
);

assign C1146=c10146+c11146+c12146+c13146;
assign A1146=(C1146>=0)?1:0;

ninexnine_unit ninexnine_unit_4780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10156)
);

ninexnine_unit ninexnine_unit_4781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11156)
);

ninexnine_unit ninexnine_unit_4782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12156)
);

ninexnine_unit ninexnine_unit_4783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13156)
);

assign C1156=c10156+c11156+c12156+c13156;
assign A1156=(C1156>=0)?1:0;

ninexnine_unit ninexnine_unit_4784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10166)
);

ninexnine_unit ninexnine_unit_4785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11166)
);

ninexnine_unit ninexnine_unit_4786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12166)
);

ninexnine_unit ninexnine_unit_4787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13166)
);

assign C1166=c10166+c11166+c12166+c13166;
assign A1166=(C1166>=0)?1:0;

ninexnine_unit ninexnine_unit_4788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10176)
);

ninexnine_unit ninexnine_unit_4789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11176)
);

ninexnine_unit ninexnine_unit_4790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12176)
);

ninexnine_unit ninexnine_unit_4791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13176)
);

assign C1176=c10176+c11176+c12176+c13176;
assign A1176=(C1176>=0)?1:0;

ninexnine_unit ninexnine_unit_4792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10186)
);

ninexnine_unit ninexnine_unit_4793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11186)
);

ninexnine_unit ninexnine_unit_4794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12186)
);

ninexnine_unit ninexnine_unit_4795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13186)
);

assign C1186=c10186+c11186+c12186+c13186;
assign A1186=(C1186>=0)?1:0;

ninexnine_unit ninexnine_unit_4796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10196)
);

ninexnine_unit ninexnine_unit_4797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11196)
);

ninexnine_unit ninexnine_unit_4798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12196)
);

ninexnine_unit ninexnine_unit_4799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13196)
);

assign C1196=c10196+c11196+c12196+c13196;
assign A1196=(C1196>=0)?1:0;

ninexnine_unit ninexnine_unit_4800(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c101A6)
);

ninexnine_unit ninexnine_unit_4801(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c111A6)
);

ninexnine_unit ninexnine_unit_4802(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c121A6)
);

ninexnine_unit ninexnine_unit_4803(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c131A6)
);

assign C11A6=c101A6+c111A6+c121A6+c131A6;
assign A11A6=(C11A6>=0)?1:0;

ninexnine_unit ninexnine_unit_4804(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c101B6)
);

ninexnine_unit ninexnine_unit_4805(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c111B6)
);

ninexnine_unit ninexnine_unit_4806(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c121B6)
);

ninexnine_unit ninexnine_unit_4807(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c131B6)
);

assign C11B6=c101B6+c111B6+c121B6+c131B6;
assign A11B6=(C11B6>=0)?1:0;

ninexnine_unit ninexnine_unit_4808(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c101C6)
);

ninexnine_unit ninexnine_unit_4809(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c111C6)
);

ninexnine_unit ninexnine_unit_4810(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c121C6)
);

ninexnine_unit ninexnine_unit_4811(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c131C6)
);

assign C11C6=c101C6+c111C6+c121C6+c131C6;
assign A11C6=(C11C6>=0)?1:0;

ninexnine_unit ninexnine_unit_4812(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c101D6)
);

ninexnine_unit ninexnine_unit_4813(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c111D6)
);

ninexnine_unit ninexnine_unit_4814(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c121D6)
);

ninexnine_unit ninexnine_unit_4815(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c131D6)
);

assign C11D6=c101D6+c111D6+c121D6+c131D6;
assign A11D6=(C11D6>=0)?1:0;

ninexnine_unit ninexnine_unit_4816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10206)
);

ninexnine_unit ninexnine_unit_4817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11206)
);

ninexnine_unit ninexnine_unit_4818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12206)
);

ninexnine_unit ninexnine_unit_4819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13206)
);

assign C1206=c10206+c11206+c12206+c13206;
assign A1206=(C1206>=0)?1:0;

ninexnine_unit ninexnine_unit_4820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10216)
);

ninexnine_unit ninexnine_unit_4821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11216)
);

ninexnine_unit ninexnine_unit_4822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12216)
);

ninexnine_unit ninexnine_unit_4823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13216)
);

assign C1216=c10216+c11216+c12216+c13216;
assign A1216=(C1216>=0)?1:0;

ninexnine_unit ninexnine_unit_4824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10226)
);

ninexnine_unit ninexnine_unit_4825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11226)
);

ninexnine_unit ninexnine_unit_4826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12226)
);

ninexnine_unit ninexnine_unit_4827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13226)
);

assign C1226=c10226+c11226+c12226+c13226;
assign A1226=(C1226>=0)?1:0;

ninexnine_unit ninexnine_unit_4828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10236)
);

ninexnine_unit ninexnine_unit_4829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11236)
);

ninexnine_unit ninexnine_unit_4830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12236)
);

ninexnine_unit ninexnine_unit_4831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13236)
);

assign C1236=c10236+c11236+c12236+c13236;
assign A1236=(C1236>=0)?1:0;

ninexnine_unit ninexnine_unit_4832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10246)
);

ninexnine_unit ninexnine_unit_4833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11246)
);

ninexnine_unit ninexnine_unit_4834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12246)
);

ninexnine_unit ninexnine_unit_4835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13246)
);

assign C1246=c10246+c11246+c12246+c13246;
assign A1246=(C1246>=0)?1:0;

ninexnine_unit ninexnine_unit_4836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10256)
);

ninexnine_unit ninexnine_unit_4837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11256)
);

ninexnine_unit ninexnine_unit_4838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12256)
);

ninexnine_unit ninexnine_unit_4839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13256)
);

assign C1256=c10256+c11256+c12256+c13256;
assign A1256=(C1256>=0)?1:0;

ninexnine_unit ninexnine_unit_4840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10266)
);

ninexnine_unit ninexnine_unit_4841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11266)
);

ninexnine_unit ninexnine_unit_4842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12266)
);

ninexnine_unit ninexnine_unit_4843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13266)
);

assign C1266=c10266+c11266+c12266+c13266;
assign A1266=(C1266>=0)?1:0;

ninexnine_unit ninexnine_unit_4844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10276)
);

ninexnine_unit ninexnine_unit_4845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11276)
);

ninexnine_unit ninexnine_unit_4846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12276)
);

ninexnine_unit ninexnine_unit_4847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13276)
);

assign C1276=c10276+c11276+c12276+c13276;
assign A1276=(C1276>=0)?1:0;

ninexnine_unit ninexnine_unit_4848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10286)
);

ninexnine_unit ninexnine_unit_4849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11286)
);

ninexnine_unit ninexnine_unit_4850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12286)
);

ninexnine_unit ninexnine_unit_4851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13286)
);

assign C1286=c10286+c11286+c12286+c13286;
assign A1286=(C1286>=0)?1:0;

ninexnine_unit ninexnine_unit_4852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10296)
);

ninexnine_unit ninexnine_unit_4853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11296)
);

ninexnine_unit ninexnine_unit_4854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12296)
);

ninexnine_unit ninexnine_unit_4855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13296)
);

assign C1296=c10296+c11296+c12296+c13296;
assign A1296=(C1296>=0)?1:0;

ninexnine_unit ninexnine_unit_4856(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c102A6)
);

ninexnine_unit ninexnine_unit_4857(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c112A6)
);

ninexnine_unit ninexnine_unit_4858(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c122A6)
);

ninexnine_unit ninexnine_unit_4859(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c132A6)
);

assign C12A6=c102A6+c112A6+c122A6+c132A6;
assign A12A6=(C12A6>=0)?1:0;

ninexnine_unit ninexnine_unit_4860(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c102B6)
);

ninexnine_unit ninexnine_unit_4861(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c112B6)
);

ninexnine_unit ninexnine_unit_4862(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c122B6)
);

ninexnine_unit ninexnine_unit_4863(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c132B6)
);

assign C12B6=c102B6+c112B6+c122B6+c132B6;
assign A12B6=(C12B6>=0)?1:0;

ninexnine_unit ninexnine_unit_4864(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c102C6)
);

ninexnine_unit ninexnine_unit_4865(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c112C6)
);

ninexnine_unit ninexnine_unit_4866(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c122C6)
);

ninexnine_unit ninexnine_unit_4867(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c132C6)
);

assign C12C6=c102C6+c112C6+c122C6+c132C6;
assign A12C6=(C12C6>=0)?1:0;

ninexnine_unit ninexnine_unit_4868(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c102D6)
);

ninexnine_unit ninexnine_unit_4869(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c112D6)
);

ninexnine_unit ninexnine_unit_4870(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c122D6)
);

ninexnine_unit ninexnine_unit_4871(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c132D6)
);

assign C12D6=c102D6+c112D6+c122D6+c132D6;
assign A12D6=(C12D6>=0)?1:0;

ninexnine_unit ninexnine_unit_4872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10306)
);

ninexnine_unit ninexnine_unit_4873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11306)
);

ninexnine_unit ninexnine_unit_4874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12306)
);

ninexnine_unit ninexnine_unit_4875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13306)
);

assign C1306=c10306+c11306+c12306+c13306;
assign A1306=(C1306>=0)?1:0;

ninexnine_unit ninexnine_unit_4876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10316)
);

ninexnine_unit ninexnine_unit_4877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11316)
);

ninexnine_unit ninexnine_unit_4878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12316)
);

ninexnine_unit ninexnine_unit_4879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13316)
);

assign C1316=c10316+c11316+c12316+c13316;
assign A1316=(C1316>=0)?1:0;

ninexnine_unit ninexnine_unit_4880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10326)
);

ninexnine_unit ninexnine_unit_4881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11326)
);

ninexnine_unit ninexnine_unit_4882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12326)
);

ninexnine_unit ninexnine_unit_4883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13326)
);

assign C1326=c10326+c11326+c12326+c13326;
assign A1326=(C1326>=0)?1:0;

ninexnine_unit ninexnine_unit_4884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10336)
);

ninexnine_unit ninexnine_unit_4885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11336)
);

ninexnine_unit ninexnine_unit_4886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12336)
);

ninexnine_unit ninexnine_unit_4887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13336)
);

assign C1336=c10336+c11336+c12336+c13336;
assign A1336=(C1336>=0)?1:0;

ninexnine_unit ninexnine_unit_4888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10346)
);

ninexnine_unit ninexnine_unit_4889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11346)
);

ninexnine_unit ninexnine_unit_4890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12346)
);

ninexnine_unit ninexnine_unit_4891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13346)
);

assign C1346=c10346+c11346+c12346+c13346;
assign A1346=(C1346>=0)?1:0;

ninexnine_unit ninexnine_unit_4892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10356)
);

ninexnine_unit ninexnine_unit_4893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11356)
);

ninexnine_unit ninexnine_unit_4894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12356)
);

ninexnine_unit ninexnine_unit_4895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13356)
);

assign C1356=c10356+c11356+c12356+c13356;
assign A1356=(C1356>=0)?1:0;

ninexnine_unit ninexnine_unit_4896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10366)
);

ninexnine_unit ninexnine_unit_4897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11366)
);

ninexnine_unit ninexnine_unit_4898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12366)
);

ninexnine_unit ninexnine_unit_4899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13366)
);

assign C1366=c10366+c11366+c12366+c13366;
assign A1366=(C1366>=0)?1:0;

ninexnine_unit ninexnine_unit_4900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10376)
);

ninexnine_unit ninexnine_unit_4901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11376)
);

ninexnine_unit ninexnine_unit_4902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12376)
);

ninexnine_unit ninexnine_unit_4903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13376)
);

assign C1376=c10376+c11376+c12376+c13376;
assign A1376=(C1376>=0)?1:0;

ninexnine_unit ninexnine_unit_4904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10386)
);

ninexnine_unit ninexnine_unit_4905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11386)
);

ninexnine_unit ninexnine_unit_4906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12386)
);

ninexnine_unit ninexnine_unit_4907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13386)
);

assign C1386=c10386+c11386+c12386+c13386;
assign A1386=(C1386>=0)?1:0;

ninexnine_unit ninexnine_unit_4908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10396)
);

ninexnine_unit ninexnine_unit_4909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11396)
);

ninexnine_unit ninexnine_unit_4910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12396)
);

ninexnine_unit ninexnine_unit_4911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13396)
);

assign C1396=c10396+c11396+c12396+c13396;
assign A1396=(C1396>=0)?1:0;

ninexnine_unit ninexnine_unit_4912(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c103A6)
);

ninexnine_unit ninexnine_unit_4913(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c113A6)
);

ninexnine_unit ninexnine_unit_4914(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c123A6)
);

ninexnine_unit ninexnine_unit_4915(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c133A6)
);

assign C13A6=c103A6+c113A6+c123A6+c133A6;
assign A13A6=(C13A6>=0)?1:0;

ninexnine_unit ninexnine_unit_4916(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c103B6)
);

ninexnine_unit ninexnine_unit_4917(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c113B6)
);

ninexnine_unit ninexnine_unit_4918(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c123B6)
);

ninexnine_unit ninexnine_unit_4919(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c133B6)
);

assign C13B6=c103B6+c113B6+c123B6+c133B6;
assign A13B6=(C13B6>=0)?1:0;

ninexnine_unit ninexnine_unit_4920(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c103C6)
);

ninexnine_unit ninexnine_unit_4921(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c113C6)
);

ninexnine_unit ninexnine_unit_4922(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c123C6)
);

ninexnine_unit ninexnine_unit_4923(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c133C6)
);

assign C13C6=c103C6+c113C6+c123C6+c133C6;
assign A13C6=(C13C6>=0)?1:0;

ninexnine_unit ninexnine_unit_4924(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c103D6)
);

ninexnine_unit ninexnine_unit_4925(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c113D6)
);

ninexnine_unit ninexnine_unit_4926(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c123D6)
);

ninexnine_unit ninexnine_unit_4927(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c133D6)
);

assign C13D6=c103D6+c113D6+c123D6+c133D6;
assign A13D6=(C13D6>=0)?1:0;

ninexnine_unit ninexnine_unit_4928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10406)
);

ninexnine_unit ninexnine_unit_4929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11406)
);

ninexnine_unit ninexnine_unit_4930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12406)
);

ninexnine_unit ninexnine_unit_4931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13406)
);

assign C1406=c10406+c11406+c12406+c13406;
assign A1406=(C1406>=0)?1:0;

ninexnine_unit ninexnine_unit_4932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10416)
);

ninexnine_unit ninexnine_unit_4933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11416)
);

ninexnine_unit ninexnine_unit_4934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12416)
);

ninexnine_unit ninexnine_unit_4935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13416)
);

assign C1416=c10416+c11416+c12416+c13416;
assign A1416=(C1416>=0)?1:0;

ninexnine_unit ninexnine_unit_4936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10426)
);

ninexnine_unit ninexnine_unit_4937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11426)
);

ninexnine_unit ninexnine_unit_4938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12426)
);

ninexnine_unit ninexnine_unit_4939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13426)
);

assign C1426=c10426+c11426+c12426+c13426;
assign A1426=(C1426>=0)?1:0;

ninexnine_unit ninexnine_unit_4940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10436)
);

ninexnine_unit ninexnine_unit_4941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11436)
);

ninexnine_unit ninexnine_unit_4942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12436)
);

ninexnine_unit ninexnine_unit_4943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13436)
);

assign C1436=c10436+c11436+c12436+c13436;
assign A1436=(C1436>=0)?1:0;

ninexnine_unit ninexnine_unit_4944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10446)
);

ninexnine_unit ninexnine_unit_4945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11446)
);

ninexnine_unit ninexnine_unit_4946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12446)
);

ninexnine_unit ninexnine_unit_4947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13446)
);

assign C1446=c10446+c11446+c12446+c13446;
assign A1446=(C1446>=0)?1:0;

ninexnine_unit ninexnine_unit_4948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10456)
);

ninexnine_unit ninexnine_unit_4949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11456)
);

ninexnine_unit ninexnine_unit_4950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12456)
);

ninexnine_unit ninexnine_unit_4951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13456)
);

assign C1456=c10456+c11456+c12456+c13456;
assign A1456=(C1456>=0)?1:0;

ninexnine_unit ninexnine_unit_4952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10466)
);

ninexnine_unit ninexnine_unit_4953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11466)
);

ninexnine_unit ninexnine_unit_4954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12466)
);

ninexnine_unit ninexnine_unit_4955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13466)
);

assign C1466=c10466+c11466+c12466+c13466;
assign A1466=(C1466>=0)?1:0;

ninexnine_unit ninexnine_unit_4956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10476)
);

ninexnine_unit ninexnine_unit_4957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11476)
);

ninexnine_unit ninexnine_unit_4958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12476)
);

ninexnine_unit ninexnine_unit_4959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13476)
);

assign C1476=c10476+c11476+c12476+c13476;
assign A1476=(C1476>=0)?1:0;

ninexnine_unit ninexnine_unit_4960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10486)
);

ninexnine_unit ninexnine_unit_4961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11486)
);

ninexnine_unit ninexnine_unit_4962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12486)
);

ninexnine_unit ninexnine_unit_4963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13486)
);

assign C1486=c10486+c11486+c12486+c13486;
assign A1486=(C1486>=0)?1:0;

ninexnine_unit ninexnine_unit_4964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10496)
);

ninexnine_unit ninexnine_unit_4965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11496)
);

ninexnine_unit ninexnine_unit_4966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12496)
);

ninexnine_unit ninexnine_unit_4967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13496)
);

assign C1496=c10496+c11496+c12496+c13496;
assign A1496=(C1496>=0)?1:0;

ninexnine_unit ninexnine_unit_4968(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c104A6)
);

ninexnine_unit ninexnine_unit_4969(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c114A6)
);

ninexnine_unit ninexnine_unit_4970(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c124A6)
);

ninexnine_unit ninexnine_unit_4971(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c134A6)
);

assign C14A6=c104A6+c114A6+c124A6+c134A6;
assign A14A6=(C14A6>=0)?1:0;

ninexnine_unit ninexnine_unit_4972(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c104B6)
);

ninexnine_unit ninexnine_unit_4973(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c114B6)
);

ninexnine_unit ninexnine_unit_4974(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c124B6)
);

ninexnine_unit ninexnine_unit_4975(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c134B6)
);

assign C14B6=c104B6+c114B6+c124B6+c134B6;
assign A14B6=(C14B6>=0)?1:0;

ninexnine_unit ninexnine_unit_4976(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c104C6)
);

ninexnine_unit ninexnine_unit_4977(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c114C6)
);

ninexnine_unit ninexnine_unit_4978(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c124C6)
);

ninexnine_unit ninexnine_unit_4979(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c134C6)
);

assign C14C6=c104C6+c114C6+c124C6+c134C6;
assign A14C6=(C14C6>=0)?1:0;

ninexnine_unit ninexnine_unit_4980(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c104D6)
);

ninexnine_unit ninexnine_unit_4981(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c114D6)
);

ninexnine_unit ninexnine_unit_4982(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c124D6)
);

ninexnine_unit ninexnine_unit_4983(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c134D6)
);

assign C14D6=c104D6+c114D6+c124D6+c134D6;
assign A14D6=(C14D6>=0)?1:0;

ninexnine_unit ninexnine_unit_4984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10506)
);

ninexnine_unit ninexnine_unit_4985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11506)
);

ninexnine_unit ninexnine_unit_4986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12506)
);

ninexnine_unit ninexnine_unit_4987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13506)
);

assign C1506=c10506+c11506+c12506+c13506;
assign A1506=(C1506>=0)?1:0;

ninexnine_unit ninexnine_unit_4988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10516)
);

ninexnine_unit ninexnine_unit_4989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11516)
);

ninexnine_unit ninexnine_unit_4990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12516)
);

ninexnine_unit ninexnine_unit_4991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13516)
);

assign C1516=c10516+c11516+c12516+c13516;
assign A1516=(C1516>=0)?1:0;

ninexnine_unit ninexnine_unit_4992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10526)
);

ninexnine_unit ninexnine_unit_4993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11526)
);

ninexnine_unit ninexnine_unit_4994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12526)
);

ninexnine_unit ninexnine_unit_4995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13526)
);

assign C1526=c10526+c11526+c12526+c13526;
assign A1526=(C1526>=0)?1:0;

ninexnine_unit ninexnine_unit_4996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10536)
);

ninexnine_unit ninexnine_unit_4997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11536)
);

ninexnine_unit ninexnine_unit_4998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12536)
);

ninexnine_unit ninexnine_unit_4999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13536)
);

assign C1536=c10536+c11536+c12536+c13536;
assign A1536=(C1536>=0)?1:0;

ninexnine_unit ninexnine_unit_5000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10546)
);

ninexnine_unit ninexnine_unit_5001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11546)
);

ninexnine_unit ninexnine_unit_5002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12546)
);

ninexnine_unit ninexnine_unit_5003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13546)
);

assign C1546=c10546+c11546+c12546+c13546;
assign A1546=(C1546>=0)?1:0;

ninexnine_unit ninexnine_unit_5004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10556)
);

ninexnine_unit ninexnine_unit_5005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11556)
);

ninexnine_unit ninexnine_unit_5006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12556)
);

ninexnine_unit ninexnine_unit_5007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13556)
);

assign C1556=c10556+c11556+c12556+c13556;
assign A1556=(C1556>=0)?1:0;

ninexnine_unit ninexnine_unit_5008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10566)
);

ninexnine_unit ninexnine_unit_5009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11566)
);

ninexnine_unit ninexnine_unit_5010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12566)
);

ninexnine_unit ninexnine_unit_5011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13566)
);

assign C1566=c10566+c11566+c12566+c13566;
assign A1566=(C1566>=0)?1:0;

ninexnine_unit ninexnine_unit_5012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10576)
);

ninexnine_unit ninexnine_unit_5013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11576)
);

ninexnine_unit ninexnine_unit_5014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12576)
);

ninexnine_unit ninexnine_unit_5015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13576)
);

assign C1576=c10576+c11576+c12576+c13576;
assign A1576=(C1576>=0)?1:0;

ninexnine_unit ninexnine_unit_5016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10586)
);

ninexnine_unit ninexnine_unit_5017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11586)
);

ninexnine_unit ninexnine_unit_5018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12586)
);

ninexnine_unit ninexnine_unit_5019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13586)
);

assign C1586=c10586+c11586+c12586+c13586;
assign A1586=(C1586>=0)?1:0;

ninexnine_unit ninexnine_unit_5020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10596)
);

ninexnine_unit ninexnine_unit_5021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11596)
);

ninexnine_unit ninexnine_unit_5022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12596)
);

ninexnine_unit ninexnine_unit_5023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13596)
);

assign C1596=c10596+c11596+c12596+c13596;
assign A1596=(C1596>=0)?1:0;

ninexnine_unit ninexnine_unit_5024(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c105A6)
);

ninexnine_unit ninexnine_unit_5025(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c115A6)
);

ninexnine_unit ninexnine_unit_5026(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c125A6)
);

ninexnine_unit ninexnine_unit_5027(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c135A6)
);

assign C15A6=c105A6+c115A6+c125A6+c135A6;
assign A15A6=(C15A6>=0)?1:0;

ninexnine_unit ninexnine_unit_5028(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c105B6)
);

ninexnine_unit ninexnine_unit_5029(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c115B6)
);

ninexnine_unit ninexnine_unit_5030(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c125B6)
);

ninexnine_unit ninexnine_unit_5031(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c135B6)
);

assign C15B6=c105B6+c115B6+c125B6+c135B6;
assign A15B6=(C15B6>=0)?1:0;

ninexnine_unit ninexnine_unit_5032(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c105C6)
);

ninexnine_unit ninexnine_unit_5033(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c115C6)
);

ninexnine_unit ninexnine_unit_5034(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c125C6)
);

ninexnine_unit ninexnine_unit_5035(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c135C6)
);

assign C15C6=c105C6+c115C6+c125C6+c135C6;
assign A15C6=(C15C6>=0)?1:0;

ninexnine_unit ninexnine_unit_5036(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c105D6)
);

ninexnine_unit ninexnine_unit_5037(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c115D6)
);

ninexnine_unit ninexnine_unit_5038(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c125D6)
);

ninexnine_unit ninexnine_unit_5039(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c135D6)
);

assign C15D6=c105D6+c115D6+c125D6+c135D6;
assign A15D6=(C15D6>=0)?1:0;

ninexnine_unit ninexnine_unit_5040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10606)
);

ninexnine_unit ninexnine_unit_5041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11606)
);

ninexnine_unit ninexnine_unit_5042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12606)
);

ninexnine_unit ninexnine_unit_5043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13606)
);

assign C1606=c10606+c11606+c12606+c13606;
assign A1606=(C1606>=0)?1:0;

ninexnine_unit ninexnine_unit_5044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10616)
);

ninexnine_unit ninexnine_unit_5045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11616)
);

ninexnine_unit ninexnine_unit_5046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12616)
);

ninexnine_unit ninexnine_unit_5047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13616)
);

assign C1616=c10616+c11616+c12616+c13616;
assign A1616=(C1616>=0)?1:0;

ninexnine_unit ninexnine_unit_5048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10626)
);

ninexnine_unit ninexnine_unit_5049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11626)
);

ninexnine_unit ninexnine_unit_5050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12626)
);

ninexnine_unit ninexnine_unit_5051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13626)
);

assign C1626=c10626+c11626+c12626+c13626;
assign A1626=(C1626>=0)?1:0;

ninexnine_unit ninexnine_unit_5052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10636)
);

ninexnine_unit ninexnine_unit_5053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11636)
);

ninexnine_unit ninexnine_unit_5054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12636)
);

ninexnine_unit ninexnine_unit_5055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13636)
);

assign C1636=c10636+c11636+c12636+c13636;
assign A1636=(C1636>=0)?1:0;

ninexnine_unit ninexnine_unit_5056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10646)
);

ninexnine_unit ninexnine_unit_5057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11646)
);

ninexnine_unit ninexnine_unit_5058(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12646)
);

ninexnine_unit ninexnine_unit_5059(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13646)
);

assign C1646=c10646+c11646+c12646+c13646;
assign A1646=(C1646>=0)?1:0;

ninexnine_unit ninexnine_unit_5060(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10656)
);

ninexnine_unit ninexnine_unit_5061(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11656)
);

ninexnine_unit ninexnine_unit_5062(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12656)
);

ninexnine_unit ninexnine_unit_5063(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13656)
);

assign C1656=c10656+c11656+c12656+c13656;
assign A1656=(C1656>=0)?1:0;

ninexnine_unit ninexnine_unit_5064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10666)
);

ninexnine_unit ninexnine_unit_5065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11666)
);

ninexnine_unit ninexnine_unit_5066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12666)
);

ninexnine_unit ninexnine_unit_5067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13666)
);

assign C1666=c10666+c11666+c12666+c13666;
assign A1666=(C1666>=0)?1:0;

ninexnine_unit ninexnine_unit_5068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10676)
);

ninexnine_unit ninexnine_unit_5069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11676)
);

ninexnine_unit ninexnine_unit_5070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12676)
);

ninexnine_unit ninexnine_unit_5071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13676)
);

assign C1676=c10676+c11676+c12676+c13676;
assign A1676=(C1676>=0)?1:0;

ninexnine_unit ninexnine_unit_5072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10686)
);

ninexnine_unit ninexnine_unit_5073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11686)
);

ninexnine_unit ninexnine_unit_5074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12686)
);

ninexnine_unit ninexnine_unit_5075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13686)
);

assign C1686=c10686+c11686+c12686+c13686;
assign A1686=(C1686>=0)?1:0;

ninexnine_unit ninexnine_unit_5076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10696)
);

ninexnine_unit ninexnine_unit_5077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11696)
);

ninexnine_unit ninexnine_unit_5078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12696)
);

ninexnine_unit ninexnine_unit_5079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13696)
);

assign C1696=c10696+c11696+c12696+c13696;
assign A1696=(C1696>=0)?1:0;

ninexnine_unit ninexnine_unit_5080(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c106A6)
);

ninexnine_unit ninexnine_unit_5081(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c116A6)
);

ninexnine_unit ninexnine_unit_5082(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c126A6)
);

ninexnine_unit ninexnine_unit_5083(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c136A6)
);

assign C16A6=c106A6+c116A6+c126A6+c136A6;
assign A16A6=(C16A6>=0)?1:0;

ninexnine_unit ninexnine_unit_5084(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c106B6)
);

ninexnine_unit ninexnine_unit_5085(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c116B6)
);

ninexnine_unit ninexnine_unit_5086(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c126B6)
);

ninexnine_unit ninexnine_unit_5087(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c136B6)
);

assign C16B6=c106B6+c116B6+c126B6+c136B6;
assign A16B6=(C16B6>=0)?1:0;

ninexnine_unit ninexnine_unit_5088(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c106C6)
);

ninexnine_unit ninexnine_unit_5089(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c116C6)
);

ninexnine_unit ninexnine_unit_5090(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c126C6)
);

ninexnine_unit ninexnine_unit_5091(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c136C6)
);

assign C16C6=c106C6+c116C6+c126C6+c136C6;
assign A16C6=(C16C6>=0)?1:0;

ninexnine_unit ninexnine_unit_5092(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c106D6)
);

ninexnine_unit ninexnine_unit_5093(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c116D6)
);

ninexnine_unit ninexnine_unit_5094(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c126D6)
);

ninexnine_unit ninexnine_unit_5095(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c136D6)
);

assign C16D6=c106D6+c116D6+c126D6+c136D6;
assign A16D6=(C16D6>=0)?1:0;

ninexnine_unit ninexnine_unit_5096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10706)
);

ninexnine_unit ninexnine_unit_5097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11706)
);

ninexnine_unit ninexnine_unit_5098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12706)
);

ninexnine_unit ninexnine_unit_5099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13706)
);

assign C1706=c10706+c11706+c12706+c13706;
assign A1706=(C1706>=0)?1:0;

ninexnine_unit ninexnine_unit_5100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10716)
);

ninexnine_unit ninexnine_unit_5101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11716)
);

ninexnine_unit ninexnine_unit_5102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12716)
);

ninexnine_unit ninexnine_unit_5103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13716)
);

assign C1716=c10716+c11716+c12716+c13716;
assign A1716=(C1716>=0)?1:0;

ninexnine_unit ninexnine_unit_5104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10726)
);

ninexnine_unit ninexnine_unit_5105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11726)
);

ninexnine_unit ninexnine_unit_5106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12726)
);

ninexnine_unit ninexnine_unit_5107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13726)
);

assign C1726=c10726+c11726+c12726+c13726;
assign A1726=(C1726>=0)?1:0;

ninexnine_unit ninexnine_unit_5108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10736)
);

ninexnine_unit ninexnine_unit_5109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11736)
);

ninexnine_unit ninexnine_unit_5110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12736)
);

ninexnine_unit ninexnine_unit_5111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13736)
);

assign C1736=c10736+c11736+c12736+c13736;
assign A1736=(C1736>=0)?1:0;

ninexnine_unit ninexnine_unit_5112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10746)
);

ninexnine_unit ninexnine_unit_5113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11746)
);

ninexnine_unit ninexnine_unit_5114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12746)
);

ninexnine_unit ninexnine_unit_5115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13746)
);

assign C1746=c10746+c11746+c12746+c13746;
assign A1746=(C1746>=0)?1:0;

ninexnine_unit ninexnine_unit_5116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10756)
);

ninexnine_unit ninexnine_unit_5117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11756)
);

ninexnine_unit ninexnine_unit_5118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12756)
);

ninexnine_unit ninexnine_unit_5119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13756)
);

assign C1756=c10756+c11756+c12756+c13756;
assign A1756=(C1756>=0)?1:0;

ninexnine_unit ninexnine_unit_5120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10766)
);

ninexnine_unit ninexnine_unit_5121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11766)
);

ninexnine_unit ninexnine_unit_5122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12766)
);

ninexnine_unit ninexnine_unit_5123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13766)
);

assign C1766=c10766+c11766+c12766+c13766;
assign A1766=(C1766>=0)?1:0;

ninexnine_unit ninexnine_unit_5124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10776)
);

ninexnine_unit ninexnine_unit_5125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11776)
);

ninexnine_unit ninexnine_unit_5126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12776)
);

ninexnine_unit ninexnine_unit_5127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13776)
);

assign C1776=c10776+c11776+c12776+c13776;
assign A1776=(C1776>=0)?1:0;

ninexnine_unit ninexnine_unit_5128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10786)
);

ninexnine_unit ninexnine_unit_5129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11786)
);

ninexnine_unit ninexnine_unit_5130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12786)
);

ninexnine_unit ninexnine_unit_5131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13786)
);

assign C1786=c10786+c11786+c12786+c13786;
assign A1786=(C1786>=0)?1:0;

ninexnine_unit ninexnine_unit_5132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10796)
);

ninexnine_unit ninexnine_unit_5133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11796)
);

ninexnine_unit ninexnine_unit_5134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12796)
);

ninexnine_unit ninexnine_unit_5135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13796)
);

assign C1796=c10796+c11796+c12796+c13796;
assign A1796=(C1796>=0)?1:0;

ninexnine_unit ninexnine_unit_5136(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c107A6)
);

ninexnine_unit ninexnine_unit_5137(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c117A6)
);

ninexnine_unit ninexnine_unit_5138(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c127A6)
);

ninexnine_unit ninexnine_unit_5139(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c137A6)
);

assign C17A6=c107A6+c117A6+c127A6+c137A6;
assign A17A6=(C17A6>=0)?1:0;

ninexnine_unit ninexnine_unit_5140(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c107B6)
);

ninexnine_unit ninexnine_unit_5141(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c117B6)
);

ninexnine_unit ninexnine_unit_5142(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c127B6)
);

ninexnine_unit ninexnine_unit_5143(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c137B6)
);

assign C17B6=c107B6+c117B6+c127B6+c137B6;
assign A17B6=(C17B6>=0)?1:0;

ninexnine_unit ninexnine_unit_5144(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c107C6)
);

ninexnine_unit ninexnine_unit_5145(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c117C6)
);

ninexnine_unit ninexnine_unit_5146(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c127C6)
);

ninexnine_unit ninexnine_unit_5147(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c137C6)
);

assign C17C6=c107C6+c117C6+c127C6+c137C6;
assign A17C6=(C17C6>=0)?1:0;

ninexnine_unit ninexnine_unit_5148(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c107D6)
);

ninexnine_unit ninexnine_unit_5149(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c117D6)
);

ninexnine_unit ninexnine_unit_5150(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c127D6)
);

ninexnine_unit ninexnine_unit_5151(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c137D6)
);

assign C17D6=c107D6+c117D6+c127D6+c137D6;
assign A17D6=(C17D6>=0)?1:0;

ninexnine_unit ninexnine_unit_5152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10806)
);

ninexnine_unit ninexnine_unit_5153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11806)
);

ninexnine_unit ninexnine_unit_5154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12806)
);

ninexnine_unit ninexnine_unit_5155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13806)
);

assign C1806=c10806+c11806+c12806+c13806;
assign A1806=(C1806>=0)?1:0;

ninexnine_unit ninexnine_unit_5156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10816)
);

ninexnine_unit ninexnine_unit_5157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11816)
);

ninexnine_unit ninexnine_unit_5158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12816)
);

ninexnine_unit ninexnine_unit_5159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13816)
);

assign C1816=c10816+c11816+c12816+c13816;
assign A1816=(C1816>=0)?1:0;

ninexnine_unit ninexnine_unit_5160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10826)
);

ninexnine_unit ninexnine_unit_5161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11826)
);

ninexnine_unit ninexnine_unit_5162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12826)
);

ninexnine_unit ninexnine_unit_5163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13826)
);

assign C1826=c10826+c11826+c12826+c13826;
assign A1826=(C1826>=0)?1:0;

ninexnine_unit ninexnine_unit_5164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10836)
);

ninexnine_unit ninexnine_unit_5165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11836)
);

ninexnine_unit ninexnine_unit_5166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12836)
);

ninexnine_unit ninexnine_unit_5167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13836)
);

assign C1836=c10836+c11836+c12836+c13836;
assign A1836=(C1836>=0)?1:0;

ninexnine_unit ninexnine_unit_5168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10846)
);

ninexnine_unit ninexnine_unit_5169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11846)
);

ninexnine_unit ninexnine_unit_5170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12846)
);

ninexnine_unit ninexnine_unit_5171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13846)
);

assign C1846=c10846+c11846+c12846+c13846;
assign A1846=(C1846>=0)?1:0;

ninexnine_unit ninexnine_unit_5172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10856)
);

ninexnine_unit ninexnine_unit_5173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11856)
);

ninexnine_unit ninexnine_unit_5174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12856)
);

ninexnine_unit ninexnine_unit_5175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13856)
);

assign C1856=c10856+c11856+c12856+c13856;
assign A1856=(C1856>=0)?1:0;

ninexnine_unit ninexnine_unit_5176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10866)
);

ninexnine_unit ninexnine_unit_5177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11866)
);

ninexnine_unit ninexnine_unit_5178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12866)
);

ninexnine_unit ninexnine_unit_5179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13866)
);

assign C1866=c10866+c11866+c12866+c13866;
assign A1866=(C1866>=0)?1:0;

ninexnine_unit ninexnine_unit_5180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10876)
);

ninexnine_unit ninexnine_unit_5181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11876)
);

ninexnine_unit ninexnine_unit_5182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12876)
);

ninexnine_unit ninexnine_unit_5183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13876)
);

assign C1876=c10876+c11876+c12876+c13876;
assign A1876=(C1876>=0)?1:0;

ninexnine_unit ninexnine_unit_5184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10886)
);

ninexnine_unit ninexnine_unit_5185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11886)
);

ninexnine_unit ninexnine_unit_5186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12886)
);

ninexnine_unit ninexnine_unit_5187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13886)
);

assign C1886=c10886+c11886+c12886+c13886;
assign A1886=(C1886>=0)?1:0;

ninexnine_unit ninexnine_unit_5188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10896)
);

ninexnine_unit ninexnine_unit_5189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11896)
);

ninexnine_unit ninexnine_unit_5190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12896)
);

ninexnine_unit ninexnine_unit_5191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13896)
);

assign C1896=c10896+c11896+c12896+c13896;
assign A1896=(C1896>=0)?1:0;

ninexnine_unit ninexnine_unit_5192(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c108A6)
);

ninexnine_unit ninexnine_unit_5193(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c118A6)
);

ninexnine_unit ninexnine_unit_5194(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c128A6)
);

ninexnine_unit ninexnine_unit_5195(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c138A6)
);

assign C18A6=c108A6+c118A6+c128A6+c138A6;
assign A18A6=(C18A6>=0)?1:0;

ninexnine_unit ninexnine_unit_5196(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c108B6)
);

ninexnine_unit ninexnine_unit_5197(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c118B6)
);

ninexnine_unit ninexnine_unit_5198(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c128B6)
);

ninexnine_unit ninexnine_unit_5199(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c138B6)
);

assign C18B6=c108B6+c118B6+c128B6+c138B6;
assign A18B6=(C18B6>=0)?1:0;

ninexnine_unit ninexnine_unit_5200(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c108C6)
);

ninexnine_unit ninexnine_unit_5201(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c118C6)
);

ninexnine_unit ninexnine_unit_5202(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c128C6)
);

ninexnine_unit ninexnine_unit_5203(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c138C6)
);

assign C18C6=c108C6+c118C6+c128C6+c138C6;
assign A18C6=(C18C6>=0)?1:0;

ninexnine_unit ninexnine_unit_5204(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c108D6)
);

ninexnine_unit ninexnine_unit_5205(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c118D6)
);

ninexnine_unit ninexnine_unit_5206(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c128D6)
);

ninexnine_unit ninexnine_unit_5207(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c138D6)
);

assign C18D6=c108D6+c118D6+c128D6+c138D6;
assign A18D6=(C18D6>=0)?1:0;

ninexnine_unit ninexnine_unit_5208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10906)
);

ninexnine_unit ninexnine_unit_5209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11906)
);

ninexnine_unit ninexnine_unit_5210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12906)
);

ninexnine_unit ninexnine_unit_5211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13906)
);

assign C1906=c10906+c11906+c12906+c13906;
assign A1906=(C1906>=0)?1:0;

ninexnine_unit ninexnine_unit_5212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10916)
);

ninexnine_unit ninexnine_unit_5213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11916)
);

ninexnine_unit ninexnine_unit_5214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12916)
);

ninexnine_unit ninexnine_unit_5215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13916)
);

assign C1916=c10916+c11916+c12916+c13916;
assign A1916=(C1916>=0)?1:0;

ninexnine_unit ninexnine_unit_5216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10926)
);

ninexnine_unit ninexnine_unit_5217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11926)
);

ninexnine_unit ninexnine_unit_5218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12926)
);

ninexnine_unit ninexnine_unit_5219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13926)
);

assign C1926=c10926+c11926+c12926+c13926;
assign A1926=(C1926>=0)?1:0;

ninexnine_unit ninexnine_unit_5220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10936)
);

ninexnine_unit ninexnine_unit_5221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11936)
);

ninexnine_unit ninexnine_unit_5222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12936)
);

ninexnine_unit ninexnine_unit_5223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13936)
);

assign C1936=c10936+c11936+c12936+c13936;
assign A1936=(C1936>=0)?1:0;

ninexnine_unit ninexnine_unit_5224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10946)
);

ninexnine_unit ninexnine_unit_5225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11946)
);

ninexnine_unit ninexnine_unit_5226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12946)
);

ninexnine_unit ninexnine_unit_5227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13946)
);

assign C1946=c10946+c11946+c12946+c13946;
assign A1946=(C1946>=0)?1:0;

ninexnine_unit ninexnine_unit_5228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10956)
);

ninexnine_unit ninexnine_unit_5229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11956)
);

ninexnine_unit ninexnine_unit_5230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12956)
);

ninexnine_unit ninexnine_unit_5231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13956)
);

assign C1956=c10956+c11956+c12956+c13956;
assign A1956=(C1956>=0)?1:0;

ninexnine_unit ninexnine_unit_5232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10966)
);

ninexnine_unit ninexnine_unit_5233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11966)
);

ninexnine_unit ninexnine_unit_5234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12966)
);

ninexnine_unit ninexnine_unit_5235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13966)
);

assign C1966=c10966+c11966+c12966+c13966;
assign A1966=(C1966>=0)?1:0;

ninexnine_unit ninexnine_unit_5236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10976)
);

ninexnine_unit ninexnine_unit_5237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11976)
);

ninexnine_unit ninexnine_unit_5238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12976)
);

ninexnine_unit ninexnine_unit_5239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13976)
);

assign C1976=c10976+c11976+c12976+c13976;
assign A1976=(C1976>=0)?1:0;

ninexnine_unit ninexnine_unit_5240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10986)
);

ninexnine_unit ninexnine_unit_5241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11986)
);

ninexnine_unit ninexnine_unit_5242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12986)
);

ninexnine_unit ninexnine_unit_5243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13986)
);

assign C1986=c10986+c11986+c12986+c13986;
assign A1986=(C1986>=0)?1:0;

ninexnine_unit ninexnine_unit_5244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10996)
);

ninexnine_unit ninexnine_unit_5245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11996)
);

ninexnine_unit ninexnine_unit_5246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12996)
);

ninexnine_unit ninexnine_unit_5247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13996)
);

assign C1996=c10996+c11996+c12996+c13996;
assign A1996=(C1996>=0)?1:0;

ninexnine_unit ninexnine_unit_5248(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c109A6)
);

ninexnine_unit ninexnine_unit_5249(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c119A6)
);

ninexnine_unit ninexnine_unit_5250(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c129A6)
);

ninexnine_unit ninexnine_unit_5251(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c139A6)
);

assign C19A6=c109A6+c119A6+c129A6+c139A6;
assign A19A6=(C19A6>=0)?1:0;

ninexnine_unit ninexnine_unit_5252(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c109B6)
);

ninexnine_unit ninexnine_unit_5253(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c119B6)
);

ninexnine_unit ninexnine_unit_5254(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c129B6)
);

ninexnine_unit ninexnine_unit_5255(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c139B6)
);

assign C19B6=c109B6+c119B6+c129B6+c139B6;
assign A19B6=(C19B6>=0)?1:0;

ninexnine_unit ninexnine_unit_5256(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c109C6)
);

ninexnine_unit ninexnine_unit_5257(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c119C6)
);

ninexnine_unit ninexnine_unit_5258(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c129C6)
);

ninexnine_unit ninexnine_unit_5259(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c139C6)
);

assign C19C6=c109C6+c119C6+c129C6+c139C6;
assign A19C6=(C19C6>=0)?1:0;

ninexnine_unit ninexnine_unit_5260(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c109D6)
);

ninexnine_unit ninexnine_unit_5261(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c119D6)
);

ninexnine_unit ninexnine_unit_5262(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c129D6)
);

ninexnine_unit ninexnine_unit_5263(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c139D6)
);

assign C19D6=c109D6+c119D6+c129D6+c139D6;
assign A19D6=(C19D6>=0)?1:0;

ninexnine_unit ninexnine_unit_5264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A06)
);

ninexnine_unit ninexnine_unit_5265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A06)
);

ninexnine_unit ninexnine_unit_5266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A06)
);

ninexnine_unit ninexnine_unit_5267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A06)
);

assign C1A06=c10A06+c11A06+c12A06+c13A06;
assign A1A06=(C1A06>=0)?1:0;

ninexnine_unit ninexnine_unit_5268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A16)
);

ninexnine_unit ninexnine_unit_5269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A16)
);

ninexnine_unit ninexnine_unit_5270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A16)
);

ninexnine_unit ninexnine_unit_5271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A16)
);

assign C1A16=c10A16+c11A16+c12A16+c13A16;
assign A1A16=(C1A16>=0)?1:0;

ninexnine_unit ninexnine_unit_5272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A26)
);

ninexnine_unit ninexnine_unit_5273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A26)
);

ninexnine_unit ninexnine_unit_5274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A26)
);

ninexnine_unit ninexnine_unit_5275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A26)
);

assign C1A26=c10A26+c11A26+c12A26+c13A26;
assign A1A26=(C1A26>=0)?1:0;

ninexnine_unit ninexnine_unit_5276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A36)
);

ninexnine_unit ninexnine_unit_5277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A36)
);

ninexnine_unit ninexnine_unit_5278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A36)
);

ninexnine_unit ninexnine_unit_5279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A36)
);

assign C1A36=c10A36+c11A36+c12A36+c13A36;
assign A1A36=(C1A36>=0)?1:0;

ninexnine_unit ninexnine_unit_5280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A46)
);

ninexnine_unit ninexnine_unit_5281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A46)
);

ninexnine_unit ninexnine_unit_5282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A46)
);

ninexnine_unit ninexnine_unit_5283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A46)
);

assign C1A46=c10A46+c11A46+c12A46+c13A46;
assign A1A46=(C1A46>=0)?1:0;

ninexnine_unit ninexnine_unit_5284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A56)
);

ninexnine_unit ninexnine_unit_5285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A56)
);

ninexnine_unit ninexnine_unit_5286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A56)
);

ninexnine_unit ninexnine_unit_5287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A56)
);

assign C1A56=c10A56+c11A56+c12A56+c13A56;
assign A1A56=(C1A56>=0)?1:0;

ninexnine_unit ninexnine_unit_5288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A66)
);

ninexnine_unit ninexnine_unit_5289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A66)
);

ninexnine_unit ninexnine_unit_5290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A66)
);

ninexnine_unit ninexnine_unit_5291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A66)
);

assign C1A66=c10A66+c11A66+c12A66+c13A66;
assign A1A66=(C1A66>=0)?1:0;

ninexnine_unit ninexnine_unit_5292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A76)
);

ninexnine_unit ninexnine_unit_5293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A76)
);

ninexnine_unit ninexnine_unit_5294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A76)
);

ninexnine_unit ninexnine_unit_5295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A76)
);

assign C1A76=c10A76+c11A76+c12A76+c13A76;
assign A1A76=(C1A76>=0)?1:0;

ninexnine_unit ninexnine_unit_5296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A86)
);

ninexnine_unit ninexnine_unit_5297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A86)
);

ninexnine_unit ninexnine_unit_5298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A86)
);

ninexnine_unit ninexnine_unit_5299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A86)
);

assign C1A86=c10A86+c11A86+c12A86+c13A86;
assign A1A86=(C1A86>=0)?1:0;

ninexnine_unit ninexnine_unit_5300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10A96)
);

ninexnine_unit ninexnine_unit_5301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11A96)
);

ninexnine_unit ninexnine_unit_5302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12A96)
);

ninexnine_unit ninexnine_unit_5303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13A96)
);

assign C1A96=c10A96+c11A96+c12A96+c13A96;
assign A1A96=(C1A96>=0)?1:0;

ninexnine_unit ninexnine_unit_5304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10AA6)
);

ninexnine_unit ninexnine_unit_5305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11AA6)
);

ninexnine_unit ninexnine_unit_5306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12AA6)
);

ninexnine_unit ninexnine_unit_5307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13AA6)
);

assign C1AA6=c10AA6+c11AA6+c12AA6+c13AA6;
assign A1AA6=(C1AA6>=0)?1:0;

ninexnine_unit ninexnine_unit_5308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10AB6)
);

ninexnine_unit ninexnine_unit_5309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11AB6)
);

ninexnine_unit ninexnine_unit_5310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12AB6)
);

ninexnine_unit ninexnine_unit_5311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13AB6)
);

assign C1AB6=c10AB6+c11AB6+c12AB6+c13AB6;
assign A1AB6=(C1AB6>=0)?1:0;

ninexnine_unit ninexnine_unit_5312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10AC6)
);

ninexnine_unit ninexnine_unit_5313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11AC6)
);

ninexnine_unit ninexnine_unit_5314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12AC6)
);

ninexnine_unit ninexnine_unit_5315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13AC6)
);

assign C1AC6=c10AC6+c11AC6+c12AC6+c13AC6;
assign A1AC6=(C1AC6>=0)?1:0;

ninexnine_unit ninexnine_unit_5316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10AD6)
);

ninexnine_unit ninexnine_unit_5317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11AD6)
);

ninexnine_unit ninexnine_unit_5318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12AD6)
);

ninexnine_unit ninexnine_unit_5319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13AD6)
);

assign C1AD6=c10AD6+c11AD6+c12AD6+c13AD6;
assign A1AD6=(C1AD6>=0)?1:0;

ninexnine_unit ninexnine_unit_5320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B06)
);

ninexnine_unit ninexnine_unit_5321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B06)
);

ninexnine_unit ninexnine_unit_5322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B06)
);

ninexnine_unit ninexnine_unit_5323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B06)
);

assign C1B06=c10B06+c11B06+c12B06+c13B06;
assign A1B06=(C1B06>=0)?1:0;

ninexnine_unit ninexnine_unit_5324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B16)
);

ninexnine_unit ninexnine_unit_5325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B16)
);

ninexnine_unit ninexnine_unit_5326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B16)
);

ninexnine_unit ninexnine_unit_5327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B16)
);

assign C1B16=c10B16+c11B16+c12B16+c13B16;
assign A1B16=(C1B16>=0)?1:0;

ninexnine_unit ninexnine_unit_5328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B26)
);

ninexnine_unit ninexnine_unit_5329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B26)
);

ninexnine_unit ninexnine_unit_5330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B26)
);

ninexnine_unit ninexnine_unit_5331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B26)
);

assign C1B26=c10B26+c11B26+c12B26+c13B26;
assign A1B26=(C1B26>=0)?1:0;

ninexnine_unit ninexnine_unit_5332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B36)
);

ninexnine_unit ninexnine_unit_5333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B36)
);

ninexnine_unit ninexnine_unit_5334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B36)
);

ninexnine_unit ninexnine_unit_5335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B36)
);

assign C1B36=c10B36+c11B36+c12B36+c13B36;
assign A1B36=(C1B36>=0)?1:0;

ninexnine_unit ninexnine_unit_5336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B46)
);

ninexnine_unit ninexnine_unit_5337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B46)
);

ninexnine_unit ninexnine_unit_5338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B46)
);

ninexnine_unit ninexnine_unit_5339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B46)
);

assign C1B46=c10B46+c11B46+c12B46+c13B46;
assign A1B46=(C1B46>=0)?1:0;

ninexnine_unit ninexnine_unit_5340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B56)
);

ninexnine_unit ninexnine_unit_5341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B56)
);

ninexnine_unit ninexnine_unit_5342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B56)
);

ninexnine_unit ninexnine_unit_5343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B56)
);

assign C1B56=c10B56+c11B56+c12B56+c13B56;
assign A1B56=(C1B56>=0)?1:0;

ninexnine_unit ninexnine_unit_5344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B66)
);

ninexnine_unit ninexnine_unit_5345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B66)
);

ninexnine_unit ninexnine_unit_5346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B66)
);

ninexnine_unit ninexnine_unit_5347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B66)
);

assign C1B66=c10B66+c11B66+c12B66+c13B66;
assign A1B66=(C1B66>=0)?1:0;

ninexnine_unit ninexnine_unit_5348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B76)
);

ninexnine_unit ninexnine_unit_5349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B76)
);

ninexnine_unit ninexnine_unit_5350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B76)
);

ninexnine_unit ninexnine_unit_5351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B76)
);

assign C1B76=c10B76+c11B76+c12B76+c13B76;
assign A1B76=(C1B76>=0)?1:0;

ninexnine_unit ninexnine_unit_5352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B86)
);

ninexnine_unit ninexnine_unit_5353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B86)
);

ninexnine_unit ninexnine_unit_5354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B86)
);

ninexnine_unit ninexnine_unit_5355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B86)
);

assign C1B86=c10B86+c11B86+c12B86+c13B86;
assign A1B86=(C1B86>=0)?1:0;

ninexnine_unit ninexnine_unit_5356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10B96)
);

ninexnine_unit ninexnine_unit_5357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11B96)
);

ninexnine_unit ninexnine_unit_5358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12B96)
);

ninexnine_unit ninexnine_unit_5359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13B96)
);

assign C1B96=c10B96+c11B96+c12B96+c13B96;
assign A1B96=(C1B96>=0)?1:0;

ninexnine_unit ninexnine_unit_5360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10BA6)
);

ninexnine_unit ninexnine_unit_5361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11BA6)
);

ninexnine_unit ninexnine_unit_5362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12BA6)
);

ninexnine_unit ninexnine_unit_5363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13BA6)
);

assign C1BA6=c10BA6+c11BA6+c12BA6+c13BA6;
assign A1BA6=(C1BA6>=0)?1:0;

ninexnine_unit ninexnine_unit_5364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10BB6)
);

ninexnine_unit ninexnine_unit_5365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11BB6)
);

ninexnine_unit ninexnine_unit_5366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12BB6)
);

ninexnine_unit ninexnine_unit_5367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13BB6)
);

assign C1BB6=c10BB6+c11BB6+c12BB6+c13BB6;
assign A1BB6=(C1BB6>=0)?1:0;

ninexnine_unit ninexnine_unit_5368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10BC6)
);

ninexnine_unit ninexnine_unit_5369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11BC6)
);

ninexnine_unit ninexnine_unit_5370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12BC6)
);

ninexnine_unit ninexnine_unit_5371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13BC6)
);

assign C1BC6=c10BC6+c11BC6+c12BC6+c13BC6;
assign A1BC6=(C1BC6>=0)?1:0;

ninexnine_unit ninexnine_unit_5372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10BD6)
);

ninexnine_unit ninexnine_unit_5373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11BD6)
);

ninexnine_unit ninexnine_unit_5374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12BD6)
);

ninexnine_unit ninexnine_unit_5375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13BD6)
);

assign C1BD6=c10BD6+c11BD6+c12BD6+c13BD6;
assign A1BD6=(C1BD6>=0)?1:0;

ninexnine_unit ninexnine_unit_5376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C06)
);

ninexnine_unit ninexnine_unit_5377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C06)
);

ninexnine_unit ninexnine_unit_5378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C06)
);

ninexnine_unit ninexnine_unit_5379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C06)
);

assign C1C06=c10C06+c11C06+c12C06+c13C06;
assign A1C06=(C1C06>=0)?1:0;

ninexnine_unit ninexnine_unit_5380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C16)
);

ninexnine_unit ninexnine_unit_5381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C16)
);

ninexnine_unit ninexnine_unit_5382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C16)
);

ninexnine_unit ninexnine_unit_5383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C16)
);

assign C1C16=c10C16+c11C16+c12C16+c13C16;
assign A1C16=(C1C16>=0)?1:0;

ninexnine_unit ninexnine_unit_5384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C26)
);

ninexnine_unit ninexnine_unit_5385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C26)
);

ninexnine_unit ninexnine_unit_5386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C26)
);

ninexnine_unit ninexnine_unit_5387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C26)
);

assign C1C26=c10C26+c11C26+c12C26+c13C26;
assign A1C26=(C1C26>=0)?1:0;

ninexnine_unit ninexnine_unit_5388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C36)
);

ninexnine_unit ninexnine_unit_5389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C36)
);

ninexnine_unit ninexnine_unit_5390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C36)
);

ninexnine_unit ninexnine_unit_5391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C36)
);

assign C1C36=c10C36+c11C36+c12C36+c13C36;
assign A1C36=(C1C36>=0)?1:0;

ninexnine_unit ninexnine_unit_5392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C46)
);

ninexnine_unit ninexnine_unit_5393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C46)
);

ninexnine_unit ninexnine_unit_5394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C46)
);

ninexnine_unit ninexnine_unit_5395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C46)
);

assign C1C46=c10C46+c11C46+c12C46+c13C46;
assign A1C46=(C1C46>=0)?1:0;

ninexnine_unit ninexnine_unit_5396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C56)
);

ninexnine_unit ninexnine_unit_5397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C56)
);

ninexnine_unit ninexnine_unit_5398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C56)
);

ninexnine_unit ninexnine_unit_5399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C56)
);

assign C1C56=c10C56+c11C56+c12C56+c13C56;
assign A1C56=(C1C56>=0)?1:0;

ninexnine_unit ninexnine_unit_5400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C66)
);

ninexnine_unit ninexnine_unit_5401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C66)
);

ninexnine_unit ninexnine_unit_5402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C66)
);

ninexnine_unit ninexnine_unit_5403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C66)
);

assign C1C66=c10C66+c11C66+c12C66+c13C66;
assign A1C66=(C1C66>=0)?1:0;

ninexnine_unit ninexnine_unit_5404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C76)
);

ninexnine_unit ninexnine_unit_5405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C76)
);

ninexnine_unit ninexnine_unit_5406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C76)
);

ninexnine_unit ninexnine_unit_5407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C76)
);

assign C1C76=c10C76+c11C76+c12C76+c13C76;
assign A1C76=(C1C76>=0)?1:0;

ninexnine_unit ninexnine_unit_5408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C86)
);

ninexnine_unit ninexnine_unit_5409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C86)
);

ninexnine_unit ninexnine_unit_5410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C86)
);

ninexnine_unit ninexnine_unit_5411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C86)
);

assign C1C86=c10C86+c11C86+c12C86+c13C86;
assign A1C86=(C1C86>=0)?1:0;

ninexnine_unit ninexnine_unit_5412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10C96)
);

ninexnine_unit ninexnine_unit_5413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11C96)
);

ninexnine_unit ninexnine_unit_5414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12C96)
);

ninexnine_unit ninexnine_unit_5415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13C96)
);

assign C1C96=c10C96+c11C96+c12C96+c13C96;
assign A1C96=(C1C96>=0)?1:0;

ninexnine_unit ninexnine_unit_5416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10CA6)
);

ninexnine_unit ninexnine_unit_5417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11CA6)
);

ninexnine_unit ninexnine_unit_5418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12CA6)
);

ninexnine_unit ninexnine_unit_5419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13CA6)
);

assign C1CA6=c10CA6+c11CA6+c12CA6+c13CA6;
assign A1CA6=(C1CA6>=0)?1:0;

ninexnine_unit ninexnine_unit_5420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10CB6)
);

ninexnine_unit ninexnine_unit_5421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11CB6)
);

ninexnine_unit ninexnine_unit_5422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12CB6)
);

ninexnine_unit ninexnine_unit_5423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13CB6)
);

assign C1CB6=c10CB6+c11CB6+c12CB6+c13CB6;
assign A1CB6=(C1CB6>=0)?1:0;

ninexnine_unit ninexnine_unit_5424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10CC6)
);

ninexnine_unit ninexnine_unit_5425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11CC6)
);

ninexnine_unit ninexnine_unit_5426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12CC6)
);

ninexnine_unit ninexnine_unit_5427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13CC6)
);

assign C1CC6=c10CC6+c11CC6+c12CC6+c13CC6;
assign A1CC6=(C1CC6>=0)?1:0;

ninexnine_unit ninexnine_unit_5428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10CD6)
);

ninexnine_unit ninexnine_unit_5429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11CD6)
);

ninexnine_unit ninexnine_unit_5430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12CD6)
);

ninexnine_unit ninexnine_unit_5431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13CD6)
);

assign C1CD6=c10CD6+c11CD6+c12CD6+c13CD6;
assign A1CD6=(C1CD6>=0)?1:0;

ninexnine_unit ninexnine_unit_5432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D06)
);

ninexnine_unit ninexnine_unit_5433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D06)
);

ninexnine_unit ninexnine_unit_5434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D06)
);

ninexnine_unit ninexnine_unit_5435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D06)
);

assign C1D06=c10D06+c11D06+c12D06+c13D06;
assign A1D06=(C1D06>=0)?1:0;

ninexnine_unit ninexnine_unit_5436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D16)
);

ninexnine_unit ninexnine_unit_5437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D16)
);

ninexnine_unit ninexnine_unit_5438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D16)
);

ninexnine_unit ninexnine_unit_5439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D16)
);

assign C1D16=c10D16+c11D16+c12D16+c13D16;
assign A1D16=(C1D16>=0)?1:0;

ninexnine_unit ninexnine_unit_5440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D26)
);

ninexnine_unit ninexnine_unit_5441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D26)
);

ninexnine_unit ninexnine_unit_5442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D26)
);

ninexnine_unit ninexnine_unit_5443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D26)
);

assign C1D26=c10D26+c11D26+c12D26+c13D26;
assign A1D26=(C1D26>=0)?1:0;

ninexnine_unit ninexnine_unit_5444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D36)
);

ninexnine_unit ninexnine_unit_5445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D36)
);

ninexnine_unit ninexnine_unit_5446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D36)
);

ninexnine_unit ninexnine_unit_5447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D36)
);

assign C1D36=c10D36+c11D36+c12D36+c13D36;
assign A1D36=(C1D36>=0)?1:0;

ninexnine_unit ninexnine_unit_5448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D46)
);

ninexnine_unit ninexnine_unit_5449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D46)
);

ninexnine_unit ninexnine_unit_5450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D46)
);

ninexnine_unit ninexnine_unit_5451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D46)
);

assign C1D46=c10D46+c11D46+c12D46+c13D46;
assign A1D46=(C1D46>=0)?1:0;

ninexnine_unit ninexnine_unit_5452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D56)
);

ninexnine_unit ninexnine_unit_5453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D56)
);

ninexnine_unit ninexnine_unit_5454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D56)
);

ninexnine_unit ninexnine_unit_5455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D56)
);

assign C1D56=c10D56+c11D56+c12D56+c13D56;
assign A1D56=(C1D56>=0)?1:0;

ninexnine_unit ninexnine_unit_5456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D66)
);

ninexnine_unit ninexnine_unit_5457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D66)
);

ninexnine_unit ninexnine_unit_5458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D66)
);

ninexnine_unit ninexnine_unit_5459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D66)
);

assign C1D66=c10D66+c11D66+c12D66+c13D66;
assign A1D66=(C1D66>=0)?1:0;

ninexnine_unit ninexnine_unit_5460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D76)
);

ninexnine_unit ninexnine_unit_5461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D76)
);

ninexnine_unit ninexnine_unit_5462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D76)
);

ninexnine_unit ninexnine_unit_5463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D76)
);

assign C1D76=c10D76+c11D76+c12D76+c13D76;
assign A1D76=(C1D76>=0)?1:0;

ninexnine_unit ninexnine_unit_5464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D86)
);

ninexnine_unit ninexnine_unit_5465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D86)
);

ninexnine_unit ninexnine_unit_5466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D86)
);

ninexnine_unit ninexnine_unit_5467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D86)
);

assign C1D86=c10D86+c11D86+c12D86+c13D86;
assign A1D86=(C1D86>=0)?1:0;

ninexnine_unit ninexnine_unit_5468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10D96)
);

ninexnine_unit ninexnine_unit_5469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11D96)
);

ninexnine_unit ninexnine_unit_5470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12D96)
);

ninexnine_unit ninexnine_unit_5471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13D96)
);

assign C1D96=c10D96+c11D96+c12D96+c13D96;
assign A1D96=(C1D96>=0)?1:0;

ninexnine_unit ninexnine_unit_5472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10DA6)
);

ninexnine_unit ninexnine_unit_5473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11DA6)
);

ninexnine_unit ninexnine_unit_5474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12DA6)
);

ninexnine_unit ninexnine_unit_5475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13DA6)
);

assign C1DA6=c10DA6+c11DA6+c12DA6+c13DA6;
assign A1DA6=(C1DA6>=0)?1:0;

ninexnine_unit ninexnine_unit_5476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10DB6)
);

ninexnine_unit ninexnine_unit_5477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11DB6)
);

ninexnine_unit ninexnine_unit_5478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12DB6)
);

ninexnine_unit ninexnine_unit_5479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13DB6)
);

assign C1DB6=c10DB6+c11DB6+c12DB6+c13DB6;
assign A1DB6=(C1DB6>=0)?1:0;

ninexnine_unit ninexnine_unit_5480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10DC6)
);

ninexnine_unit ninexnine_unit_5481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11DC6)
);

ninexnine_unit ninexnine_unit_5482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12DC6)
);

ninexnine_unit ninexnine_unit_5483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13DC6)
);

assign C1DC6=c10DC6+c11DC6+c12DC6+c13DC6;
assign A1DC6=(C1DC6>=0)?1:0;

ninexnine_unit ninexnine_unit_5484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10DD6)
);

ninexnine_unit ninexnine_unit_5485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11DD6)
);

ninexnine_unit ninexnine_unit_5486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12DD6)
);

ninexnine_unit ninexnine_unit_5487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13DD6)
);

assign C1DD6=c10DD6+c11DD6+c12DD6+c13DD6;
assign A1DD6=(C1DD6>=0)?1:0;

ninexnine_unit ninexnine_unit_5488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10007)
);

ninexnine_unit ninexnine_unit_5489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11007)
);

ninexnine_unit ninexnine_unit_5490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12007)
);

ninexnine_unit ninexnine_unit_5491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13007)
);

assign C1007=c10007+c11007+c12007+c13007;
assign A1007=(C1007>=0)?1:0;

ninexnine_unit ninexnine_unit_5492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10017)
);

ninexnine_unit ninexnine_unit_5493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11017)
);

ninexnine_unit ninexnine_unit_5494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12017)
);

ninexnine_unit ninexnine_unit_5495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13017)
);

assign C1017=c10017+c11017+c12017+c13017;
assign A1017=(C1017>=0)?1:0;

ninexnine_unit ninexnine_unit_5496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10027)
);

ninexnine_unit ninexnine_unit_5497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11027)
);

ninexnine_unit ninexnine_unit_5498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12027)
);

ninexnine_unit ninexnine_unit_5499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13027)
);

assign C1027=c10027+c11027+c12027+c13027;
assign A1027=(C1027>=0)?1:0;

ninexnine_unit ninexnine_unit_5500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10037)
);

ninexnine_unit ninexnine_unit_5501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11037)
);

ninexnine_unit ninexnine_unit_5502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12037)
);

ninexnine_unit ninexnine_unit_5503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1033),
				.a1(P1043),
				.a2(P1053),
				.a3(P1133),
				.a4(P1143),
				.a5(P1153),
				.a6(P1233),
				.a7(P1243),
				.a8(P1253),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13037)
);

assign C1037=c10037+c11037+c12037+c13037;
assign A1037=(C1037>=0)?1:0;

ninexnine_unit ninexnine_unit_5504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10047)
);

ninexnine_unit ninexnine_unit_5505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11047)
);

ninexnine_unit ninexnine_unit_5506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12047)
);

ninexnine_unit ninexnine_unit_5507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1043),
				.a1(P1053),
				.a2(P1063),
				.a3(P1143),
				.a4(P1153),
				.a5(P1163),
				.a6(P1243),
				.a7(P1253),
				.a8(P1263),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13047)
);

assign C1047=c10047+c11047+c12047+c13047;
assign A1047=(C1047>=0)?1:0;

ninexnine_unit ninexnine_unit_5508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1050),
				.a1(P1060),
				.a2(P1070),
				.a3(P1150),
				.a4(P1160),
				.a5(P1170),
				.a6(P1250),
				.a7(P1260),
				.a8(P1270),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10057)
);

ninexnine_unit ninexnine_unit_5509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1051),
				.a1(P1061),
				.a2(P1071),
				.a3(P1151),
				.a4(P1161),
				.a5(P1171),
				.a6(P1251),
				.a7(P1261),
				.a8(P1271),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11057)
);

ninexnine_unit ninexnine_unit_5510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1052),
				.a1(P1062),
				.a2(P1072),
				.a3(P1152),
				.a4(P1162),
				.a5(P1172),
				.a6(P1252),
				.a7(P1262),
				.a8(P1272),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12057)
);

ninexnine_unit ninexnine_unit_5511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1053),
				.a1(P1063),
				.a2(P1073),
				.a3(P1153),
				.a4(P1163),
				.a5(P1173),
				.a6(P1253),
				.a7(P1263),
				.a8(P1273),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13057)
);

assign C1057=c10057+c11057+c12057+c13057;
assign A1057=(C1057>=0)?1:0;

ninexnine_unit ninexnine_unit_5512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1060),
				.a1(P1070),
				.a2(P1080),
				.a3(P1160),
				.a4(P1170),
				.a5(P1180),
				.a6(P1260),
				.a7(P1270),
				.a8(P1280),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10067)
);

ninexnine_unit ninexnine_unit_5513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1061),
				.a1(P1071),
				.a2(P1081),
				.a3(P1161),
				.a4(P1171),
				.a5(P1181),
				.a6(P1261),
				.a7(P1271),
				.a8(P1281),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11067)
);

ninexnine_unit ninexnine_unit_5514(
				.clk(clk),
				.rstn(rstn),
				.a0(P1062),
				.a1(P1072),
				.a2(P1082),
				.a3(P1162),
				.a4(P1172),
				.a5(P1182),
				.a6(P1262),
				.a7(P1272),
				.a8(P1282),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12067)
);

ninexnine_unit ninexnine_unit_5515(
				.clk(clk),
				.rstn(rstn),
				.a0(P1063),
				.a1(P1073),
				.a2(P1083),
				.a3(P1163),
				.a4(P1173),
				.a5(P1183),
				.a6(P1263),
				.a7(P1273),
				.a8(P1283),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13067)
);

assign C1067=c10067+c11067+c12067+c13067;
assign A1067=(C1067>=0)?1:0;

ninexnine_unit ninexnine_unit_5516(
				.clk(clk),
				.rstn(rstn),
				.a0(P1070),
				.a1(P1080),
				.a2(P1090),
				.a3(P1170),
				.a4(P1180),
				.a5(P1190),
				.a6(P1270),
				.a7(P1280),
				.a8(P1290),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10077)
);

ninexnine_unit ninexnine_unit_5517(
				.clk(clk),
				.rstn(rstn),
				.a0(P1071),
				.a1(P1081),
				.a2(P1091),
				.a3(P1171),
				.a4(P1181),
				.a5(P1191),
				.a6(P1271),
				.a7(P1281),
				.a8(P1291),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11077)
);

ninexnine_unit ninexnine_unit_5518(
				.clk(clk),
				.rstn(rstn),
				.a0(P1072),
				.a1(P1082),
				.a2(P1092),
				.a3(P1172),
				.a4(P1182),
				.a5(P1192),
				.a6(P1272),
				.a7(P1282),
				.a8(P1292),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12077)
);

ninexnine_unit ninexnine_unit_5519(
				.clk(clk),
				.rstn(rstn),
				.a0(P1073),
				.a1(P1083),
				.a2(P1093),
				.a3(P1173),
				.a4(P1183),
				.a5(P1193),
				.a6(P1273),
				.a7(P1283),
				.a8(P1293),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13077)
);

assign C1077=c10077+c11077+c12077+c13077;
assign A1077=(C1077>=0)?1:0;

ninexnine_unit ninexnine_unit_5520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1080),
				.a1(P1090),
				.a2(P10A0),
				.a3(P1180),
				.a4(P1190),
				.a5(P11A0),
				.a6(P1280),
				.a7(P1290),
				.a8(P12A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10087)
);

ninexnine_unit ninexnine_unit_5521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1081),
				.a1(P1091),
				.a2(P10A1),
				.a3(P1181),
				.a4(P1191),
				.a5(P11A1),
				.a6(P1281),
				.a7(P1291),
				.a8(P12A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11087)
);

ninexnine_unit ninexnine_unit_5522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1082),
				.a1(P1092),
				.a2(P10A2),
				.a3(P1182),
				.a4(P1192),
				.a5(P11A2),
				.a6(P1282),
				.a7(P1292),
				.a8(P12A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12087)
);

ninexnine_unit ninexnine_unit_5523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1083),
				.a1(P1093),
				.a2(P10A3),
				.a3(P1183),
				.a4(P1193),
				.a5(P11A3),
				.a6(P1283),
				.a7(P1293),
				.a8(P12A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13087)
);

assign C1087=c10087+c11087+c12087+c13087;
assign A1087=(C1087>=0)?1:0;

ninexnine_unit ninexnine_unit_5524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1090),
				.a1(P10A0),
				.a2(P10B0),
				.a3(P1190),
				.a4(P11A0),
				.a5(P11B0),
				.a6(P1290),
				.a7(P12A0),
				.a8(P12B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10097)
);

ninexnine_unit ninexnine_unit_5525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1091),
				.a1(P10A1),
				.a2(P10B1),
				.a3(P1191),
				.a4(P11A1),
				.a5(P11B1),
				.a6(P1291),
				.a7(P12A1),
				.a8(P12B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11097)
);

ninexnine_unit ninexnine_unit_5526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1092),
				.a1(P10A2),
				.a2(P10B2),
				.a3(P1192),
				.a4(P11A2),
				.a5(P11B2),
				.a6(P1292),
				.a7(P12A2),
				.a8(P12B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12097)
);

ninexnine_unit ninexnine_unit_5527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1093),
				.a1(P10A3),
				.a2(P10B3),
				.a3(P1193),
				.a4(P11A3),
				.a5(P11B3),
				.a6(P1293),
				.a7(P12A3),
				.a8(P12B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13097)
);

assign C1097=c10097+c11097+c12097+c13097;
assign A1097=(C1097>=0)?1:0;

ninexnine_unit ninexnine_unit_5528(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A0),
				.a1(P10B0),
				.a2(P10C0),
				.a3(P11A0),
				.a4(P11B0),
				.a5(P11C0),
				.a6(P12A0),
				.a7(P12B0),
				.a8(P12C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c100A7)
);

ninexnine_unit ninexnine_unit_5529(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A1),
				.a1(P10B1),
				.a2(P10C1),
				.a3(P11A1),
				.a4(P11B1),
				.a5(P11C1),
				.a6(P12A1),
				.a7(P12B1),
				.a8(P12C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c110A7)
);

ninexnine_unit ninexnine_unit_5530(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A2),
				.a1(P10B2),
				.a2(P10C2),
				.a3(P11A2),
				.a4(P11B2),
				.a5(P11C2),
				.a6(P12A2),
				.a7(P12B2),
				.a8(P12C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c120A7)
);

ninexnine_unit ninexnine_unit_5531(
				.clk(clk),
				.rstn(rstn),
				.a0(P10A3),
				.a1(P10B3),
				.a2(P10C3),
				.a3(P11A3),
				.a4(P11B3),
				.a5(P11C3),
				.a6(P12A3),
				.a7(P12B3),
				.a8(P12C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c130A7)
);

assign C10A7=c100A7+c110A7+c120A7+c130A7;
assign A10A7=(C10A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5532(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B0),
				.a1(P10C0),
				.a2(P10D0),
				.a3(P11B0),
				.a4(P11C0),
				.a5(P11D0),
				.a6(P12B0),
				.a7(P12C0),
				.a8(P12D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c100B7)
);

ninexnine_unit ninexnine_unit_5533(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B1),
				.a1(P10C1),
				.a2(P10D1),
				.a3(P11B1),
				.a4(P11C1),
				.a5(P11D1),
				.a6(P12B1),
				.a7(P12C1),
				.a8(P12D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c110B7)
);

ninexnine_unit ninexnine_unit_5534(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B2),
				.a1(P10C2),
				.a2(P10D2),
				.a3(P11B2),
				.a4(P11C2),
				.a5(P11D2),
				.a6(P12B2),
				.a7(P12C2),
				.a8(P12D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c120B7)
);

ninexnine_unit ninexnine_unit_5535(
				.clk(clk),
				.rstn(rstn),
				.a0(P10B3),
				.a1(P10C3),
				.a2(P10D3),
				.a3(P11B3),
				.a4(P11C3),
				.a5(P11D3),
				.a6(P12B3),
				.a7(P12C3),
				.a8(P12D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c130B7)
);

assign C10B7=c100B7+c110B7+c120B7+c130B7;
assign A10B7=(C10B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5536(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C0),
				.a1(P10D0),
				.a2(P10E0),
				.a3(P11C0),
				.a4(P11D0),
				.a5(P11E0),
				.a6(P12C0),
				.a7(P12D0),
				.a8(P12E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c100C7)
);

ninexnine_unit ninexnine_unit_5537(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C1),
				.a1(P10D1),
				.a2(P10E1),
				.a3(P11C1),
				.a4(P11D1),
				.a5(P11E1),
				.a6(P12C1),
				.a7(P12D1),
				.a8(P12E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c110C7)
);

ninexnine_unit ninexnine_unit_5538(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C2),
				.a1(P10D2),
				.a2(P10E2),
				.a3(P11C2),
				.a4(P11D2),
				.a5(P11E2),
				.a6(P12C2),
				.a7(P12D2),
				.a8(P12E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c120C7)
);

ninexnine_unit ninexnine_unit_5539(
				.clk(clk),
				.rstn(rstn),
				.a0(P10C3),
				.a1(P10D3),
				.a2(P10E3),
				.a3(P11C3),
				.a4(P11D3),
				.a5(P11E3),
				.a6(P12C3),
				.a7(P12D3),
				.a8(P12E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c130C7)
);

assign C10C7=c100C7+c110C7+c120C7+c130C7;
assign A10C7=(C10C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5540(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D0),
				.a1(P10E0),
				.a2(P10F0),
				.a3(P11D0),
				.a4(P11E0),
				.a5(P11F0),
				.a6(P12D0),
				.a7(P12E0),
				.a8(P12F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c100D7)
);

ninexnine_unit ninexnine_unit_5541(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D1),
				.a1(P10E1),
				.a2(P10F1),
				.a3(P11D1),
				.a4(P11E1),
				.a5(P11F1),
				.a6(P12D1),
				.a7(P12E1),
				.a8(P12F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c110D7)
);

ninexnine_unit ninexnine_unit_5542(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D2),
				.a1(P10E2),
				.a2(P10F2),
				.a3(P11D2),
				.a4(P11E2),
				.a5(P11F2),
				.a6(P12D2),
				.a7(P12E2),
				.a8(P12F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c120D7)
);

ninexnine_unit ninexnine_unit_5543(
				.clk(clk),
				.rstn(rstn),
				.a0(P10D3),
				.a1(P10E3),
				.a2(P10F3),
				.a3(P11D3),
				.a4(P11E3),
				.a5(P11F3),
				.a6(P12D3),
				.a7(P12E3),
				.a8(P12F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c130D7)
);

assign C10D7=c100D7+c110D7+c120D7+c130D7;
assign A10D7=(C10D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10107)
);

ninexnine_unit ninexnine_unit_5545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11107)
);

ninexnine_unit ninexnine_unit_5546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12107)
);

ninexnine_unit ninexnine_unit_5547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13107)
);

assign C1107=c10107+c11107+c12107+c13107;
assign A1107=(C1107>=0)?1:0;

ninexnine_unit ninexnine_unit_5548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10117)
);

ninexnine_unit ninexnine_unit_5549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11117)
);

ninexnine_unit ninexnine_unit_5550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12117)
);

ninexnine_unit ninexnine_unit_5551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13117)
);

assign C1117=c10117+c11117+c12117+c13117;
assign A1117=(C1117>=0)?1:0;

ninexnine_unit ninexnine_unit_5552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10127)
);

ninexnine_unit ninexnine_unit_5553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11127)
);

ninexnine_unit ninexnine_unit_5554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12127)
);

ninexnine_unit ninexnine_unit_5555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13127)
);

assign C1127=c10127+c11127+c12127+c13127;
assign A1127=(C1127>=0)?1:0;

ninexnine_unit ninexnine_unit_5556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10137)
);

ninexnine_unit ninexnine_unit_5557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11137)
);

ninexnine_unit ninexnine_unit_5558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12137)
);

ninexnine_unit ninexnine_unit_5559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1133),
				.a1(P1143),
				.a2(P1153),
				.a3(P1233),
				.a4(P1243),
				.a5(P1253),
				.a6(P1333),
				.a7(P1343),
				.a8(P1353),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13137)
);

assign C1137=c10137+c11137+c12137+c13137;
assign A1137=(C1137>=0)?1:0;

ninexnine_unit ninexnine_unit_5560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10147)
);

ninexnine_unit ninexnine_unit_5561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11147)
);

ninexnine_unit ninexnine_unit_5562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12147)
);

ninexnine_unit ninexnine_unit_5563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1143),
				.a1(P1153),
				.a2(P1163),
				.a3(P1243),
				.a4(P1253),
				.a5(P1263),
				.a6(P1343),
				.a7(P1353),
				.a8(P1363),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13147)
);

assign C1147=c10147+c11147+c12147+c13147;
assign A1147=(C1147>=0)?1:0;

ninexnine_unit ninexnine_unit_5564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1150),
				.a1(P1160),
				.a2(P1170),
				.a3(P1250),
				.a4(P1260),
				.a5(P1270),
				.a6(P1350),
				.a7(P1360),
				.a8(P1370),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10157)
);

ninexnine_unit ninexnine_unit_5565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1151),
				.a1(P1161),
				.a2(P1171),
				.a3(P1251),
				.a4(P1261),
				.a5(P1271),
				.a6(P1351),
				.a7(P1361),
				.a8(P1371),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11157)
);

ninexnine_unit ninexnine_unit_5566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1152),
				.a1(P1162),
				.a2(P1172),
				.a3(P1252),
				.a4(P1262),
				.a5(P1272),
				.a6(P1352),
				.a7(P1362),
				.a8(P1372),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12157)
);

ninexnine_unit ninexnine_unit_5567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1153),
				.a1(P1163),
				.a2(P1173),
				.a3(P1253),
				.a4(P1263),
				.a5(P1273),
				.a6(P1353),
				.a7(P1363),
				.a8(P1373),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13157)
);

assign C1157=c10157+c11157+c12157+c13157;
assign A1157=(C1157>=0)?1:0;

ninexnine_unit ninexnine_unit_5568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1160),
				.a1(P1170),
				.a2(P1180),
				.a3(P1260),
				.a4(P1270),
				.a5(P1280),
				.a6(P1360),
				.a7(P1370),
				.a8(P1380),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10167)
);

ninexnine_unit ninexnine_unit_5569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1161),
				.a1(P1171),
				.a2(P1181),
				.a3(P1261),
				.a4(P1271),
				.a5(P1281),
				.a6(P1361),
				.a7(P1371),
				.a8(P1381),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11167)
);

ninexnine_unit ninexnine_unit_5570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1162),
				.a1(P1172),
				.a2(P1182),
				.a3(P1262),
				.a4(P1272),
				.a5(P1282),
				.a6(P1362),
				.a7(P1372),
				.a8(P1382),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12167)
);

ninexnine_unit ninexnine_unit_5571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1163),
				.a1(P1173),
				.a2(P1183),
				.a3(P1263),
				.a4(P1273),
				.a5(P1283),
				.a6(P1363),
				.a7(P1373),
				.a8(P1383),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13167)
);

assign C1167=c10167+c11167+c12167+c13167;
assign A1167=(C1167>=0)?1:0;

ninexnine_unit ninexnine_unit_5572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1170),
				.a1(P1180),
				.a2(P1190),
				.a3(P1270),
				.a4(P1280),
				.a5(P1290),
				.a6(P1370),
				.a7(P1380),
				.a8(P1390),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10177)
);

ninexnine_unit ninexnine_unit_5573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1171),
				.a1(P1181),
				.a2(P1191),
				.a3(P1271),
				.a4(P1281),
				.a5(P1291),
				.a6(P1371),
				.a7(P1381),
				.a8(P1391),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11177)
);

ninexnine_unit ninexnine_unit_5574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1172),
				.a1(P1182),
				.a2(P1192),
				.a3(P1272),
				.a4(P1282),
				.a5(P1292),
				.a6(P1372),
				.a7(P1382),
				.a8(P1392),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12177)
);

ninexnine_unit ninexnine_unit_5575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1173),
				.a1(P1183),
				.a2(P1193),
				.a3(P1273),
				.a4(P1283),
				.a5(P1293),
				.a6(P1373),
				.a7(P1383),
				.a8(P1393),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13177)
);

assign C1177=c10177+c11177+c12177+c13177;
assign A1177=(C1177>=0)?1:0;

ninexnine_unit ninexnine_unit_5576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1180),
				.a1(P1190),
				.a2(P11A0),
				.a3(P1280),
				.a4(P1290),
				.a5(P12A0),
				.a6(P1380),
				.a7(P1390),
				.a8(P13A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10187)
);

ninexnine_unit ninexnine_unit_5577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1181),
				.a1(P1191),
				.a2(P11A1),
				.a3(P1281),
				.a4(P1291),
				.a5(P12A1),
				.a6(P1381),
				.a7(P1391),
				.a8(P13A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11187)
);

ninexnine_unit ninexnine_unit_5578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1182),
				.a1(P1192),
				.a2(P11A2),
				.a3(P1282),
				.a4(P1292),
				.a5(P12A2),
				.a6(P1382),
				.a7(P1392),
				.a8(P13A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12187)
);

ninexnine_unit ninexnine_unit_5579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1183),
				.a1(P1193),
				.a2(P11A3),
				.a3(P1283),
				.a4(P1293),
				.a5(P12A3),
				.a6(P1383),
				.a7(P1393),
				.a8(P13A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13187)
);

assign C1187=c10187+c11187+c12187+c13187;
assign A1187=(C1187>=0)?1:0;

ninexnine_unit ninexnine_unit_5580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1190),
				.a1(P11A0),
				.a2(P11B0),
				.a3(P1290),
				.a4(P12A0),
				.a5(P12B0),
				.a6(P1390),
				.a7(P13A0),
				.a8(P13B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10197)
);

ninexnine_unit ninexnine_unit_5581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1191),
				.a1(P11A1),
				.a2(P11B1),
				.a3(P1291),
				.a4(P12A1),
				.a5(P12B1),
				.a6(P1391),
				.a7(P13A1),
				.a8(P13B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11197)
);

ninexnine_unit ninexnine_unit_5582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1192),
				.a1(P11A2),
				.a2(P11B2),
				.a3(P1292),
				.a4(P12A2),
				.a5(P12B2),
				.a6(P1392),
				.a7(P13A2),
				.a8(P13B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12197)
);

ninexnine_unit ninexnine_unit_5583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1193),
				.a1(P11A3),
				.a2(P11B3),
				.a3(P1293),
				.a4(P12A3),
				.a5(P12B3),
				.a6(P1393),
				.a7(P13A3),
				.a8(P13B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13197)
);

assign C1197=c10197+c11197+c12197+c13197;
assign A1197=(C1197>=0)?1:0;

ninexnine_unit ninexnine_unit_5584(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A0),
				.a1(P11B0),
				.a2(P11C0),
				.a3(P12A0),
				.a4(P12B0),
				.a5(P12C0),
				.a6(P13A0),
				.a7(P13B0),
				.a8(P13C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c101A7)
);

ninexnine_unit ninexnine_unit_5585(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A1),
				.a1(P11B1),
				.a2(P11C1),
				.a3(P12A1),
				.a4(P12B1),
				.a5(P12C1),
				.a6(P13A1),
				.a7(P13B1),
				.a8(P13C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c111A7)
);

ninexnine_unit ninexnine_unit_5586(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A2),
				.a1(P11B2),
				.a2(P11C2),
				.a3(P12A2),
				.a4(P12B2),
				.a5(P12C2),
				.a6(P13A2),
				.a7(P13B2),
				.a8(P13C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c121A7)
);

ninexnine_unit ninexnine_unit_5587(
				.clk(clk),
				.rstn(rstn),
				.a0(P11A3),
				.a1(P11B3),
				.a2(P11C3),
				.a3(P12A3),
				.a4(P12B3),
				.a5(P12C3),
				.a6(P13A3),
				.a7(P13B3),
				.a8(P13C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c131A7)
);

assign C11A7=c101A7+c111A7+c121A7+c131A7;
assign A11A7=(C11A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5588(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B0),
				.a1(P11C0),
				.a2(P11D0),
				.a3(P12B0),
				.a4(P12C0),
				.a5(P12D0),
				.a6(P13B0),
				.a7(P13C0),
				.a8(P13D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c101B7)
);

ninexnine_unit ninexnine_unit_5589(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B1),
				.a1(P11C1),
				.a2(P11D1),
				.a3(P12B1),
				.a4(P12C1),
				.a5(P12D1),
				.a6(P13B1),
				.a7(P13C1),
				.a8(P13D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c111B7)
);

ninexnine_unit ninexnine_unit_5590(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B2),
				.a1(P11C2),
				.a2(P11D2),
				.a3(P12B2),
				.a4(P12C2),
				.a5(P12D2),
				.a6(P13B2),
				.a7(P13C2),
				.a8(P13D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c121B7)
);

ninexnine_unit ninexnine_unit_5591(
				.clk(clk),
				.rstn(rstn),
				.a0(P11B3),
				.a1(P11C3),
				.a2(P11D3),
				.a3(P12B3),
				.a4(P12C3),
				.a5(P12D3),
				.a6(P13B3),
				.a7(P13C3),
				.a8(P13D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c131B7)
);

assign C11B7=c101B7+c111B7+c121B7+c131B7;
assign A11B7=(C11B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5592(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C0),
				.a1(P11D0),
				.a2(P11E0),
				.a3(P12C0),
				.a4(P12D0),
				.a5(P12E0),
				.a6(P13C0),
				.a7(P13D0),
				.a8(P13E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c101C7)
);

ninexnine_unit ninexnine_unit_5593(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C1),
				.a1(P11D1),
				.a2(P11E1),
				.a3(P12C1),
				.a4(P12D1),
				.a5(P12E1),
				.a6(P13C1),
				.a7(P13D1),
				.a8(P13E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c111C7)
);

ninexnine_unit ninexnine_unit_5594(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C2),
				.a1(P11D2),
				.a2(P11E2),
				.a3(P12C2),
				.a4(P12D2),
				.a5(P12E2),
				.a6(P13C2),
				.a7(P13D2),
				.a8(P13E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c121C7)
);

ninexnine_unit ninexnine_unit_5595(
				.clk(clk),
				.rstn(rstn),
				.a0(P11C3),
				.a1(P11D3),
				.a2(P11E3),
				.a3(P12C3),
				.a4(P12D3),
				.a5(P12E3),
				.a6(P13C3),
				.a7(P13D3),
				.a8(P13E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c131C7)
);

assign C11C7=c101C7+c111C7+c121C7+c131C7;
assign A11C7=(C11C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5596(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D0),
				.a1(P11E0),
				.a2(P11F0),
				.a3(P12D0),
				.a4(P12E0),
				.a5(P12F0),
				.a6(P13D0),
				.a7(P13E0),
				.a8(P13F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c101D7)
);

ninexnine_unit ninexnine_unit_5597(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D1),
				.a1(P11E1),
				.a2(P11F1),
				.a3(P12D1),
				.a4(P12E1),
				.a5(P12F1),
				.a6(P13D1),
				.a7(P13E1),
				.a8(P13F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c111D7)
);

ninexnine_unit ninexnine_unit_5598(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D2),
				.a1(P11E2),
				.a2(P11F2),
				.a3(P12D2),
				.a4(P12E2),
				.a5(P12F2),
				.a6(P13D2),
				.a7(P13E2),
				.a8(P13F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c121D7)
);

ninexnine_unit ninexnine_unit_5599(
				.clk(clk),
				.rstn(rstn),
				.a0(P11D3),
				.a1(P11E3),
				.a2(P11F3),
				.a3(P12D3),
				.a4(P12E3),
				.a5(P12F3),
				.a6(P13D3),
				.a7(P13E3),
				.a8(P13F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c131D7)
);

assign C11D7=c101D7+c111D7+c121D7+c131D7;
assign A11D7=(C11D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10207)
);

ninexnine_unit ninexnine_unit_5601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11207)
);

ninexnine_unit ninexnine_unit_5602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12207)
);

ninexnine_unit ninexnine_unit_5603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13207)
);

assign C1207=c10207+c11207+c12207+c13207;
assign A1207=(C1207>=0)?1:0;

ninexnine_unit ninexnine_unit_5604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10217)
);

ninexnine_unit ninexnine_unit_5605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11217)
);

ninexnine_unit ninexnine_unit_5606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12217)
);

ninexnine_unit ninexnine_unit_5607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13217)
);

assign C1217=c10217+c11217+c12217+c13217;
assign A1217=(C1217>=0)?1:0;

ninexnine_unit ninexnine_unit_5608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10227)
);

ninexnine_unit ninexnine_unit_5609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11227)
);

ninexnine_unit ninexnine_unit_5610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12227)
);

ninexnine_unit ninexnine_unit_5611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13227)
);

assign C1227=c10227+c11227+c12227+c13227;
assign A1227=(C1227>=0)?1:0;

ninexnine_unit ninexnine_unit_5612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10237)
);

ninexnine_unit ninexnine_unit_5613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11237)
);

ninexnine_unit ninexnine_unit_5614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12237)
);

ninexnine_unit ninexnine_unit_5615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1233),
				.a1(P1243),
				.a2(P1253),
				.a3(P1333),
				.a4(P1343),
				.a5(P1353),
				.a6(P1433),
				.a7(P1443),
				.a8(P1453),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13237)
);

assign C1237=c10237+c11237+c12237+c13237;
assign A1237=(C1237>=0)?1:0;

ninexnine_unit ninexnine_unit_5616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10247)
);

ninexnine_unit ninexnine_unit_5617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11247)
);

ninexnine_unit ninexnine_unit_5618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12247)
);

ninexnine_unit ninexnine_unit_5619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1243),
				.a1(P1253),
				.a2(P1263),
				.a3(P1343),
				.a4(P1353),
				.a5(P1363),
				.a6(P1443),
				.a7(P1453),
				.a8(P1463),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13247)
);

assign C1247=c10247+c11247+c12247+c13247;
assign A1247=(C1247>=0)?1:0;

ninexnine_unit ninexnine_unit_5620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1250),
				.a1(P1260),
				.a2(P1270),
				.a3(P1350),
				.a4(P1360),
				.a5(P1370),
				.a6(P1450),
				.a7(P1460),
				.a8(P1470),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10257)
);

ninexnine_unit ninexnine_unit_5621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1251),
				.a1(P1261),
				.a2(P1271),
				.a3(P1351),
				.a4(P1361),
				.a5(P1371),
				.a6(P1451),
				.a7(P1461),
				.a8(P1471),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11257)
);

ninexnine_unit ninexnine_unit_5622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1252),
				.a1(P1262),
				.a2(P1272),
				.a3(P1352),
				.a4(P1362),
				.a5(P1372),
				.a6(P1452),
				.a7(P1462),
				.a8(P1472),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12257)
);

ninexnine_unit ninexnine_unit_5623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1253),
				.a1(P1263),
				.a2(P1273),
				.a3(P1353),
				.a4(P1363),
				.a5(P1373),
				.a6(P1453),
				.a7(P1463),
				.a8(P1473),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13257)
);

assign C1257=c10257+c11257+c12257+c13257;
assign A1257=(C1257>=0)?1:0;

ninexnine_unit ninexnine_unit_5624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1260),
				.a1(P1270),
				.a2(P1280),
				.a3(P1360),
				.a4(P1370),
				.a5(P1380),
				.a6(P1460),
				.a7(P1470),
				.a8(P1480),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10267)
);

ninexnine_unit ninexnine_unit_5625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1261),
				.a1(P1271),
				.a2(P1281),
				.a3(P1361),
				.a4(P1371),
				.a5(P1381),
				.a6(P1461),
				.a7(P1471),
				.a8(P1481),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11267)
);

ninexnine_unit ninexnine_unit_5626(
				.clk(clk),
				.rstn(rstn),
				.a0(P1262),
				.a1(P1272),
				.a2(P1282),
				.a3(P1362),
				.a4(P1372),
				.a5(P1382),
				.a6(P1462),
				.a7(P1472),
				.a8(P1482),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12267)
);

ninexnine_unit ninexnine_unit_5627(
				.clk(clk),
				.rstn(rstn),
				.a0(P1263),
				.a1(P1273),
				.a2(P1283),
				.a3(P1363),
				.a4(P1373),
				.a5(P1383),
				.a6(P1463),
				.a7(P1473),
				.a8(P1483),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13267)
);

assign C1267=c10267+c11267+c12267+c13267;
assign A1267=(C1267>=0)?1:0;

ninexnine_unit ninexnine_unit_5628(
				.clk(clk),
				.rstn(rstn),
				.a0(P1270),
				.a1(P1280),
				.a2(P1290),
				.a3(P1370),
				.a4(P1380),
				.a5(P1390),
				.a6(P1470),
				.a7(P1480),
				.a8(P1490),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10277)
);

ninexnine_unit ninexnine_unit_5629(
				.clk(clk),
				.rstn(rstn),
				.a0(P1271),
				.a1(P1281),
				.a2(P1291),
				.a3(P1371),
				.a4(P1381),
				.a5(P1391),
				.a6(P1471),
				.a7(P1481),
				.a8(P1491),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11277)
);

ninexnine_unit ninexnine_unit_5630(
				.clk(clk),
				.rstn(rstn),
				.a0(P1272),
				.a1(P1282),
				.a2(P1292),
				.a3(P1372),
				.a4(P1382),
				.a5(P1392),
				.a6(P1472),
				.a7(P1482),
				.a8(P1492),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12277)
);

ninexnine_unit ninexnine_unit_5631(
				.clk(clk),
				.rstn(rstn),
				.a0(P1273),
				.a1(P1283),
				.a2(P1293),
				.a3(P1373),
				.a4(P1383),
				.a5(P1393),
				.a6(P1473),
				.a7(P1483),
				.a8(P1493),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13277)
);

assign C1277=c10277+c11277+c12277+c13277;
assign A1277=(C1277>=0)?1:0;

ninexnine_unit ninexnine_unit_5632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1280),
				.a1(P1290),
				.a2(P12A0),
				.a3(P1380),
				.a4(P1390),
				.a5(P13A0),
				.a6(P1480),
				.a7(P1490),
				.a8(P14A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10287)
);

ninexnine_unit ninexnine_unit_5633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1281),
				.a1(P1291),
				.a2(P12A1),
				.a3(P1381),
				.a4(P1391),
				.a5(P13A1),
				.a6(P1481),
				.a7(P1491),
				.a8(P14A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11287)
);

ninexnine_unit ninexnine_unit_5634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1282),
				.a1(P1292),
				.a2(P12A2),
				.a3(P1382),
				.a4(P1392),
				.a5(P13A2),
				.a6(P1482),
				.a7(P1492),
				.a8(P14A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12287)
);

ninexnine_unit ninexnine_unit_5635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1283),
				.a1(P1293),
				.a2(P12A3),
				.a3(P1383),
				.a4(P1393),
				.a5(P13A3),
				.a6(P1483),
				.a7(P1493),
				.a8(P14A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13287)
);

assign C1287=c10287+c11287+c12287+c13287;
assign A1287=(C1287>=0)?1:0;

ninexnine_unit ninexnine_unit_5636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1290),
				.a1(P12A0),
				.a2(P12B0),
				.a3(P1390),
				.a4(P13A0),
				.a5(P13B0),
				.a6(P1490),
				.a7(P14A0),
				.a8(P14B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10297)
);

ninexnine_unit ninexnine_unit_5637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1291),
				.a1(P12A1),
				.a2(P12B1),
				.a3(P1391),
				.a4(P13A1),
				.a5(P13B1),
				.a6(P1491),
				.a7(P14A1),
				.a8(P14B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11297)
);

ninexnine_unit ninexnine_unit_5638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1292),
				.a1(P12A2),
				.a2(P12B2),
				.a3(P1392),
				.a4(P13A2),
				.a5(P13B2),
				.a6(P1492),
				.a7(P14A2),
				.a8(P14B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12297)
);

ninexnine_unit ninexnine_unit_5639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1293),
				.a1(P12A3),
				.a2(P12B3),
				.a3(P1393),
				.a4(P13A3),
				.a5(P13B3),
				.a6(P1493),
				.a7(P14A3),
				.a8(P14B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13297)
);

assign C1297=c10297+c11297+c12297+c13297;
assign A1297=(C1297>=0)?1:0;

ninexnine_unit ninexnine_unit_5640(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A0),
				.a1(P12B0),
				.a2(P12C0),
				.a3(P13A0),
				.a4(P13B0),
				.a5(P13C0),
				.a6(P14A0),
				.a7(P14B0),
				.a8(P14C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c102A7)
);

ninexnine_unit ninexnine_unit_5641(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A1),
				.a1(P12B1),
				.a2(P12C1),
				.a3(P13A1),
				.a4(P13B1),
				.a5(P13C1),
				.a6(P14A1),
				.a7(P14B1),
				.a8(P14C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c112A7)
);

ninexnine_unit ninexnine_unit_5642(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A2),
				.a1(P12B2),
				.a2(P12C2),
				.a3(P13A2),
				.a4(P13B2),
				.a5(P13C2),
				.a6(P14A2),
				.a7(P14B2),
				.a8(P14C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c122A7)
);

ninexnine_unit ninexnine_unit_5643(
				.clk(clk),
				.rstn(rstn),
				.a0(P12A3),
				.a1(P12B3),
				.a2(P12C3),
				.a3(P13A3),
				.a4(P13B3),
				.a5(P13C3),
				.a6(P14A3),
				.a7(P14B3),
				.a8(P14C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c132A7)
);

assign C12A7=c102A7+c112A7+c122A7+c132A7;
assign A12A7=(C12A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5644(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B0),
				.a1(P12C0),
				.a2(P12D0),
				.a3(P13B0),
				.a4(P13C0),
				.a5(P13D0),
				.a6(P14B0),
				.a7(P14C0),
				.a8(P14D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c102B7)
);

ninexnine_unit ninexnine_unit_5645(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B1),
				.a1(P12C1),
				.a2(P12D1),
				.a3(P13B1),
				.a4(P13C1),
				.a5(P13D1),
				.a6(P14B1),
				.a7(P14C1),
				.a8(P14D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c112B7)
);

ninexnine_unit ninexnine_unit_5646(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B2),
				.a1(P12C2),
				.a2(P12D2),
				.a3(P13B2),
				.a4(P13C2),
				.a5(P13D2),
				.a6(P14B2),
				.a7(P14C2),
				.a8(P14D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c122B7)
);

ninexnine_unit ninexnine_unit_5647(
				.clk(clk),
				.rstn(rstn),
				.a0(P12B3),
				.a1(P12C3),
				.a2(P12D3),
				.a3(P13B3),
				.a4(P13C3),
				.a5(P13D3),
				.a6(P14B3),
				.a7(P14C3),
				.a8(P14D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c132B7)
);

assign C12B7=c102B7+c112B7+c122B7+c132B7;
assign A12B7=(C12B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5648(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C0),
				.a1(P12D0),
				.a2(P12E0),
				.a3(P13C0),
				.a4(P13D0),
				.a5(P13E0),
				.a6(P14C0),
				.a7(P14D0),
				.a8(P14E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c102C7)
);

ninexnine_unit ninexnine_unit_5649(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C1),
				.a1(P12D1),
				.a2(P12E1),
				.a3(P13C1),
				.a4(P13D1),
				.a5(P13E1),
				.a6(P14C1),
				.a7(P14D1),
				.a8(P14E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c112C7)
);

ninexnine_unit ninexnine_unit_5650(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C2),
				.a1(P12D2),
				.a2(P12E2),
				.a3(P13C2),
				.a4(P13D2),
				.a5(P13E2),
				.a6(P14C2),
				.a7(P14D2),
				.a8(P14E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c122C7)
);

ninexnine_unit ninexnine_unit_5651(
				.clk(clk),
				.rstn(rstn),
				.a0(P12C3),
				.a1(P12D3),
				.a2(P12E3),
				.a3(P13C3),
				.a4(P13D3),
				.a5(P13E3),
				.a6(P14C3),
				.a7(P14D3),
				.a8(P14E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c132C7)
);

assign C12C7=c102C7+c112C7+c122C7+c132C7;
assign A12C7=(C12C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5652(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D0),
				.a1(P12E0),
				.a2(P12F0),
				.a3(P13D0),
				.a4(P13E0),
				.a5(P13F0),
				.a6(P14D0),
				.a7(P14E0),
				.a8(P14F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c102D7)
);

ninexnine_unit ninexnine_unit_5653(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D1),
				.a1(P12E1),
				.a2(P12F1),
				.a3(P13D1),
				.a4(P13E1),
				.a5(P13F1),
				.a6(P14D1),
				.a7(P14E1),
				.a8(P14F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c112D7)
);

ninexnine_unit ninexnine_unit_5654(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D2),
				.a1(P12E2),
				.a2(P12F2),
				.a3(P13D2),
				.a4(P13E2),
				.a5(P13F2),
				.a6(P14D2),
				.a7(P14E2),
				.a8(P14F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c122D7)
);

ninexnine_unit ninexnine_unit_5655(
				.clk(clk),
				.rstn(rstn),
				.a0(P12D3),
				.a1(P12E3),
				.a2(P12F3),
				.a3(P13D3),
				.a4(P13E3),
				.a5(P13F3),
				.a6(P14D3),
				.a7(P14E3),
				.a8(P14F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c132D7)
);

assign C12D7=c102D7+c112D7+c122D7+c132D7;
assign A12D7=(C12D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10307)
);

ninexnine_unit ninexnine_unit_5657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11307)
);

ninexnine_unit ninexnine_unit_5658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12307)
);

ninexnine_unit ninexnine_unit_5659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1303),
				.a1(P1313),
				.a2(P1323),
				.a3(P1403),
				.a4(P1413),
				.a5(P1423),
				.a6(P1503),
				.a7(P1513),
				.a8(P1523),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13307)
);

assign C1307=c10307+c11307+c12307+c13307;
assign A1307=(C1307>=0)?1:0;

ninexnine_unit ninexnine_unit_5660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10317)
);

ninexnine_unit ninexnine_unit_5661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11317)
);

ninexnine_unit ninexnine_unit_5662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12317)
);

ninexnine_unit ninexnine_unit_5663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1313),
				.a1(P1323),
				.a2(P1333),
				.a3(P1413),
				.a4(P1423),
				.a5(P1433),
				.a6(P1513),
				.a7(P1523),
				.a8(P1533),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13317)
);

assign C1317=c10317+c11317+c12317+c13317;
assign A1317=(C1317>=0)?1:0;

ninexnine_unit ninexnine_unit_5664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10327)
);

ninexnine_unit ninexnine_unit_5665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11327)
);

ninexnine_unit ninexnine_unit_5666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12327)
);

ninexnine_unit ninexnine_unit_5667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1323),
				.a1(P1333),
				.a2(P1343),
				.a3(P1423),
				.a4(P1433),
				.a5(P1443),
				.a6(P1523),
				.a7(P1533),
				.a8(P1543),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13327)
);

assign C1327=c10327+c11327+c12327+c13327;
assign A1327=(C1327>=0)?1:0;

ninexnine_unit ninexnine_unit_5668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10337)
);

ninexnine_unit ninexnine_unit_5669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11337)
);

ninexnine_unit ninexnine_unit_5670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12337)
);

ninexnine_unit ninexnine_unit_5671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1333),
				.a1(P1343),
				.a2(P1353),
				.a3(P1433),
				.a4(P1443),
				.a5(P1453),
				.a6(P1533),
				.a7(P1543),
				.a8(P1553),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13337)
);

assign C1337=c10337+c11337+c12337+c13337;
assign A1337=(C1337>=0)?1:0;

ninexnine_unit ninexnine_unit_5672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10347)
);

ninexnine_unit ninexnine_unit_5673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11347)
);

ninexnine_unit ninexnine_unit_5674(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12347)
);

ninexnine_unit ninexnine_unit_5675(
				.clk(clk),
				.rstn(rstn),
				.a0(P1343),
				.a1(P1353),
				.a2(P1363),
				.a3(P1443),
				.a4(P1453),
				.a5(P1463),
				.a6(P1543),
				.a7(P1553),
				.a8(P1563),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13347)
);

assign C1347=c10347+c11347+c12347+c13347;
assign A1347=(C1347>=0)?1:0;

ninexnine_unit ninexnine_unit_5676(
				.clk(clk),
				.rstn(rstn),
				.a0(P1350),
				.a1(P1360),
				.a2(P1370),
				.a3(P1450),
				.a4(P1460),
				.a5(P1470),
				.a6(P1550),
				.a7(P1560),
				.a8(P1570),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10357)
);

ninexnine_unit ninexnine_unit_5677(
				.clk(clk),
				.rstn(rstn),
				.a0(P1351),
				.a1(P1361),
				.a2(P1371),
				.a3(P1451),
				.a4(P1461),
				.a5(P1471),
				.a6(P1551),
				.a7(P1561),
				.a8(P1571),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11357)
);

ninexnine_unit ninexnine_unit_5678(
				.clk(clk),
				.rstn(rstn),
				.a0(P1352),
				.a1(P1362),
				.a2(P1372),
				.a3(P1452),
				.a4(P1462),
				.a5(P1472),
				.a6(P1552),
				.a7(P1562),
				.a8(P1572),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12357)
);

ninexnine_unit ninexnine_unit_5679(
				.clk(clk),
				.rstn(rstn),
				.a0(P1353),
				.a1(P1363),
				.a2(P1373),
				.a3(P1453),
				.a4(P1463),
				.a5(P1473),
				.a6(P1553),
				.a7(P1563),
				.a8(P1573),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13357)
);

assign C1357=c10357+c11357+c12357+c13357;
assign A1357=(C1357>=0)?1:0;

ninexnine_unit ninexnine_unit_5680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1360),
				.a1(P1370),
				.a2(P1380),
				.a3(P1460),
				.a4(P1470),
				.a5(P1480),
				.a6(P1560),
				.a7(P1570),
				.a8(P1580),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10367)
);

ninexnine_unit ninexnine_unit_5681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1361),
				.a1(P1371),
				.a2(P1381),
				.a3(P1461),
				.a4(P1471),
				.a5(P1481),
				.a6(P1561),
				.a7(P1571),
				.a8(P1581),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11367)
);

ninexnine_unit ninexnine_unit_5682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1362),
				.a1(P1372),
				.a2(P1382),
				.a3(P1462),
				.a4(P1472),
				.a5(P1482),
				.a6(P1562),
				.a7(P1572),
				.a8(P1582),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12367)
);

ninexnine_unit ninexnine_unit_5683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1363),
				.a1(P1373),
				.a2(P1383),
				.a3(P1463),
				.a4(P1473),
				.a5(P1483),
				.a6(P1563),
				.a7(P1573),
				.a8(P1583),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13367)
);

assign C1367=c10367+c11367+c12367+c13367;
assign A1367=(C1367>=0)?1:0;

ninexnine_unit ninexnine_unit_5684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1370),
				.a1(P1380),
				.a2(P1390),
				.a3(P1470),
				.a4(P1480),
				.a5(P1490),
				.a6(P1570),
				.a7(P1580),
				.a8(P1590),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10377)
);

ninexnine_unit ninexnine_unit_5685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1371),
				.a1(P1381),
				.a2(P1391),
				.a3(P1471),
				.a4(P1481),
				.a5(P1491),
				.a6(P1571),
				.a7(P1581),
				.a8(P1591),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11377)
);

ninexnine_unit ninexnine_unit_5686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1372),
				.a1(P1382),
				.a2(P1392),
				.a3(P1472),
				.a4(P1482),
				.a5(P1492),
				.a6(P1572),
				.a7(P1582),
				.a8(P1592),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12377)
);

ninexnine_unit ninexnine_unit_5687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1373),
				.a1(P1383),
				.a2(P1393),
				.a3(P1473),
				.a4(P1483),
				.a5(P1493),
				.a6(P1573),
				.a7(P1583),
				.a8(P1593),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13377)
);

assign C1377=c10377+c11377+c12377+c13377;
assign A1377=(C1377>=0)?1:0;

ninexnine_unit ninexnine_unit_5688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1380),
				.a1(P1390),
				.a2(P13A0),
				.a3(P1480),
				.a4(P1490),
				.a5(P14A0),
				.a6(P1580),
				.a7(P1590),
				.a8(P15A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10387)
);

ninexnine_unit ninexnine_unit_5689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1381),
				.a1(P1391),
				.a2(P13A1),
				.a3(P1481),
				.a4(P1491),
				.a5(P14A1),
				.a6(P1581),
				.a7(P1591),
				.a8(P15A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11387)
);

ninexnine_unit ninexnine_unit_5690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1382),
				.a1(P1392),
				.a2(P13A2),
				.a3(P1482),
				.a4(P1492),
				.a5(P14A2),
				.a6(P1582),
				.a7(P1592),
				.a8(P15A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12387)
);

ninexnine_unit ninexnine_unit_5691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1383),
				.a1(P1393),
				.a2(P13A3),
				.a3(P1483),
				.a4(P1493),
				.a5(P14A3),
				.a6(P1583),
				.a7(P1593),
				.a8(P15A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13387)
);

assign C1387=c10387+c11387+c12387+c13387;
assign A1387=(C1387>=0)?1:0;

ninexnine_unit ninexnine_unit_5692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1390),
				.a1(P13A0),
				.a2(P13B0),
				.a3(P1490),
				.a4(P14A0),
				.a5(P14B0),
				.a6(P1590),
				.a7(P15A0),
				.a8(P15B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10397)
);

ninexnine_unit ninexnine_unit_5693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1391),
				.a1(P13A1),
				.a2(P13B1),
				.a3(P1491),
				.a4(P14A1),
				.a5(P14B1),
				.a6(P1591),
				.a7(P15A1),
				.a8(P15B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11397)
);

ninexnine_unit ninexnine_unit_5694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1392),
				.a1(P13A2),
				.a2(P13B2),
				.a3(P1492),
				.a4(P14A2),
				.a5(P14B2),
				.a6(P1592),
				.a7(P15A2),
				.a8(P15B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12397)
);

ninexnine_unit ninexnine_unit_5695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1393),
				.a1(P13A3),
				.a2(P13B3),
				.a3(P1493),
				.a4(P14A3),
				.a5(P14B3),
				.a6(P1593),
				.a7(P15A3),
				.a8(P15B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13397)
);

assign C1397=c10397+c11397+c12397+c13397;
assign A1397=(C1397>=0)?1:0;

ninexnine_unit ninexnine_unit_5696(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A0),
				.a1(P13B0),
				.a2(P13C0),
				.a3(P14A0),
				.a4(P14B0),
				.a5(P14C0),
				.a6(P15A0),
				.a7(P15B0),
				.a8(P15C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c103A7)
);

ninexnine_unit ninexnine_unit_5697(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A1),
				.a1(P13B1),
				.a2(P13C1),
				.a3(P14A1),
				.a4(P14B1),
				.a5(P14C1),
				.a6(P15A1),
				.a7(P15B1),
				.a8(P15C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c113A7)
);

ninexnine_unit ninexnine_unit_5698(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A2),
				.a1(P13B2),
				.a2(P13C2),
				.a3(P14A2),
				.a4(P14B2),
				.a5(P14C2),
				.a6(P15A2),
				.a7(P15B2),
				.a8(P15C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c123A7)
);

ninexnine_unit ninexnine_unit_5699(
				.clk(clk),
				.rstn(rstn),
				.a0(P13A3),
				.a1(P13B3),
				.a2(P13C3),
				.a3(P14A3),
				.a4(P14B3),
				.a5(P14C3),
				.a6(P15A3),
				.a7(P15B3),
				.a8(P15C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c133A7)
);

assign C13A7=c103A7+c113A7+c123A7+c133A7;
assign A13A7=(C13A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5700(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B0),
				.a1(P13C0),
				.a2(P13D0),
				.a3(P14B0),
				.a4(P14C0),
				.a5(P14D0),
				.a6(P15B0),
				.a7(P15C0),
				.a8(P15D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c103B7)
);

ninexnine_unit ninexnine_unit_5701(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B1),
				.a1(P13C1),
				.a2(P13D1),
				.a3(P14B1),
				.a4(P14C1),
				.a5(P14D1),
				.a6(P15B1),
				.a7(P15C1),
				.a8(P15D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c113B7)
);

ninexnine_unit ninexnine_unit_5702(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B2),
				.a1(P13C2),
				.a2(P13D2),
				.a3(P14B2),
				.a4(P14C2),
				.a5(P14D2),
				.a6(P15B2),
				.a7(P15C2),
				.a8(P15D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c123B7)
);

ninexnine_unit ninexnine_unit_5703(
				.clk(clk),
				.rstn(rstn),
				.a0(P13B3),
				.a1(P13C3),
				.a2(P13D3),
				.a3(P14B3),
				.a4(P14C3),
				.a5(P14D3),
				.a6(P15B3),
				.a7(P15C3),
				.a8(P15D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c133B7)
);

assign C13B7=c103B7+c113B7+c123B7+c133B7;
assign A13B7=(C13B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5704(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C0),
				.a1(P13D0),
				.a2(P13E0),
				.a3(P14C0),
				.a4(P14D0),
				.a5(P14E0),
				.a6(P15C0),
				.a7(P15D0),
				.a8(P15E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c103C7)
);

ninexnine_unit ninexnine_unit_5705(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C1),
				.a1(P13D1),
				.a2(P13E1),
				.a3(P14C1),
				.a4(P14D1),
				.a5(P14E1),
				.a6(P15C1),
				.a7(P15D1),
				.a8(P15E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c113C7)
);

ninexnine_unit ninexnine_unit_5706(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C2),
				.a1(P13D2),
				.a2(P13E2),
				.a3(P14C2),
				.a4(P14D2),
				.a5(P14E2),
				.a6(P15C2),
				.a7(P15D2),
				.a8(P15E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c123C7)
);

ninexnine_unit ninexnine_unit_5707(
				.clk(clk),
				.rstn(rstn),
				.a0(P13C3),
				.a1(P13D3),
				.a2(P13E3),
				.a3(P14C3),
				.a4(P14D3),
				.a5(P14E3),
				.a6(P15C3),
				.a7(P15D3),
				.a8(P15E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c133C7)
);

assign C13C7=c103C7+c113C7+c123C7+c133C7;
assign A13C7=(C13C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5708(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D0),
				.a1(P13E0),
				.a2(P13F0),
				.a3(P14D0),
				.a4(P14E0),
				.a5(P14F0),
				.a6(P15D0),
				.a7(P15E0),
				.a8(P15F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c103D7)
);

ninexnine_unit ninexnine_unit_5709(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D1),
				.a1(P13E1),
				.a2(P13F1),
				.a3(P14D1),
				.a4(P14E1),
				.a5(P14F1),
				.a6(P15D1),
				.a7(P15E1),
				.a8(P15F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c113D7)
);

ninexnine_unit ninexnine_unit_5710(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D2),
				.a1(P13E2),
				.a2(P13F2),
				.a3(P14D2),
				.a4(P14E2),
				.a5(P14F2),
				.a6(P15D2),
				.a7(P15E2),
				.a8(P15F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c123D7)
);

ninexnine_unit ninexnine_unit_5711(
				.clk(clk),
				.rstn(rstn),
				.a0(P13D3),
				.a1(P13E3),
				.a2(P13F3),
				.a3(P14D3),
				.a4(P14E3),
				.a5(P14F3),
				.a6(P15D3),
				.a7(P15E3),
				.a8(P15F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c133D7)
);

assign C13D7=c103D7+c113D7+c123D7+c133D7;
assign A13D7=(C13D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10407)
);

ninexnine_unit ninexnine_unit_5713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11407)
);

ninexnine_unit ninexnine_unit_5714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12407)
);

ninexnine_unit ninexnine_unit_5715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1403),
				.a1(P1413),
				.a2(P1423),
				.a3(P1503),
				.a4(P1513),
				.a5(P1523),
				.a6(P1603),
				.a7(P1613),
				.a8(P1623),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13407)
);

assign C1407=c10407+c11407+c12407+c13407;
assign A1407=(C1407>=0)?1:0;

ninexnine_unit ninexnine_unit_5716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10417)
);

ninexnine_unit ninexnine_unit_5717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11417)
);

ninexnine_unit ninexnine_unit_5718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12417)
);

ninexnine_unit ninexnine_unit_5719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1413),
				.a1(P1423),
				.a2(P1433),
				.a3(P1513),
				.a4(P1523),
				.a5(P1533),
				.a6(P1613),
				.a7(P1623),
				.a8(P1633),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13417)
);

assign C1417=c10417+c11417+c12417+c13417;
assign A1417=(C1417>=0)?1:0;

ninexnine_unit ninexnine_unit_5720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10427)
);

ninexnine_unit ninexnine_unit_5721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11427)
);

ninexnine_unit ninexnine_unit_5722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12427)
);

ninexnine_unit ninexnine_unit_5723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1423),
				.a1(P1433),
				.a2(P1443),
				.a3(P1523),
				.a4(P1533),
				.a5(P1543),
				.a6(P1623),
				.a7(P1633),
				.a8(P1643),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13427)
);

assign C1427=c10427+c11427+c12427+c13427;
assign A1427=(C1427>=0)?1:0;

ninexnine_unit ninexnine_unit_5724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10437)
);

ninexnine_unit ninexnine_unit_5725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11437)
);

ninexnine_unit ninexnine_unit_5726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12437)
);

ninexnine_unit ninexnine_unit_5727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1433),
				.a1(P1443),
				.a2(P1453),
				.a3(P1533),
				.a4(P1543),
				.a5(P1553),
				.a6(P1633),
				.a7(P1643),
				.a8(P1653),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13437)
);

assign C1437=c10437+c11437+c12437+c13437;
assign A1437=(C1437>=0)?1:0;

ninexnine_unit ninexnine_unit_5728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10447)
);

ninexnine_unit ninexnine_unit_5729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11447)
);

ninexnine_unit ninexnine_unit_5730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12447)
);

ninexnine_unit ninexnine_unit_5731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1443),
				.a1(P1453),
				.a2(P1463),
				.a3(P1543),
				.a4(P1553),
				.a5(P1563),
				.a6(P1643),
				.a7(P1653),
				.a8(P1663),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13447)
);

assign C1447=c10447+c11447+c12447+c13447;
assign A1447=(C1447>=0)?1:0;

ninexnine_unit ninexnine_unit_5732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1450),
				.a1(P1460),
				.a2(P1470),
				.a3(P1550),
				.a4(P1560),
				.a5(P1570),
				.a6(P1650),
				.a7(P1660),
				.a8(P1670),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10457)
);

ninexnine_unit ninexnine_unit_5733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1451),
				.a1(P1461),
				.a2(P1471),
				.a3(P1551),
				.a4(P1561),
				.a5(P1571),
				.a6(P1651),
				.a7(P1661),
				.a8(P1671),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11457)
);

ninexnine_unit ninexnine_unit_5734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1452),
				.a1(P1462),
				.a2(P1472),
				.a3(P1552),
				.a4(P1562),
				.a5(P1572),
				.a6(P1652),
				.a7(P1662),
				.a8(P1672),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12457)
);

ninexnine_unit ninexnine_unit_5735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1453),
				.a1(P1463),
				.a2(P1473),
				.a3(P1553),
				.a4(P1563),
				.a5(P1573),
				.a6(P1653),
				.a7(P1663),
				.a8(P1673),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13457)
);

assign C1457=c10457+c11457+c12457+c13457;
assign A1457=(C1457>=0)?1:0;

ninexnine_unit ninexnine_unit_5736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1460),
				.a1(P1470),
				.a2(P1480),
				.a3(P1560),
				.a4(P1570),
				.a5(P1580),
				.a6(P1660),
				.a7(P1670),
				.a8(P1680),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10467)
);

ninexnine_unit ninexnine_unit_5737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1461),
				.a1(P1471),
				.a2(P1481),
				.a3(P1561),
				.a4(P1571),
				.a5(P1581),
				.a6(P1661),
				.a7(P1671),
				.a8(P1681),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11467)
);

ninexnine_unit ninexnine_unit_5738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1462),
				.a1(P1472),
				.a2(P1482),
				.a3(P1562),
				.a4(P1572),
				.a5(P1582),
				.a6(P1662),
				.a7(P1672),
				.a8(P1682),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12467)
);

ninexnine_unit ninexnine_unit_5739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1463),
				.a1(P1473),
				.a2(P1483),
				.a3(P1563),
				.a4(P1573),
				.a5(P1583),
				.a6(P1663),
				.a7(P1673),
				.a8(P1683),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13467)
);

assign C1467=c10467+c11467+c12467+c13467;
assign A1467=(C1467>=0)?1:0;

ninexnine_unit ninexnine_unit_5740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1470),
				.a1(P1480),
				.a2(P1490),
				.a3(P1570),
				.a4(P1580),
				.a5(P1590),
				.a6(P1670),
				.a7(P1680),
				.a8(P1690),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10477)
);

ninexnine_unit ninexnine_unit_5741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1471),
				.a1(P1481),
				.a2(P1491),
				.a3(P1571),
				.a4(P1581),
				.a5(P1591),
				.a6(P1671),
				.a7(P1681),
				.a8(P1691),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11477)
);

ninexnine_unit ninexnine_unit_5742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1472),
				.a1(P1482),
				.a2(P1492),
				.a3(P1572),
				.a4(P1582),
				.a5(P1592),
				.a6(P1672),
				.a7(P1682),
				.a8(P1692),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12477)
);

ninexnine_unit ninexnine_unit_5743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1473),
				.a1(P1483),
				.a2(P1493),
				.a3(P1573),
				.a4(P1583),
				.a5(P1593),
				.a6(P1673),
				.a7(P1683),
				.a8(P1693),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13477)
);

assign C1477=c10477+c11477+c12477+c13477;
assign A1477=(C1477>=0)?1:0;

ninexnine_unit ninexnine_unit_5744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1480),
				.a1(P1490),
				.a2(P14A0),
				.a3(P1580),
				.a4(P1590),
				.a5(P15A0),
				.a6(P1680),
				.a7(P1690),
				.a8(P16A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10487)
);

ninexnine_unit ninexnine_unit_5745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1481),
				.a1(P1491),
				.a2(P14A1),
				.a3(P1581),
				.a4(P1591),
				.a5(P15A1),
				.a6(P1681),
				.a7(P1691),
				.a8(P16A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11487)
);

ninexnine_unit ninexnine_unit_5746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1482),
				.a1(P1492),
				.a2(P14A2),
				.a3(P1582),
				.a4(P1592),
				.a5(P15A2),
				.a6(P1682),
				.a7(P1692),
				.a8(P16A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12487)
);

ninexnine_unit ninexnine_unit_5747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1483),
				.a1(P1493),
				.a2(P14A3),
				.a3(P1583),
				.a4(P1593),
				.a5(P15A3),
				.a6(P1683),
				.a7(P1693),
				.a8(P16A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13487)
);

assign C1487=c10487+c11487+c12487+c13487;
assign A1487=(C1487>=0)?1:0;

ninexnine_unit ninexnine_unit_5748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1490),
				.a1(P14A0),
				.a2(P14B0),
				.a3(P1590),
				.a4(P15A0),
				.a5(P15B0),
				.a6(P1690),
				.a7(P16A0),
				.a8(P16B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10497)
);

ninexnine_unit ninexnine_unit_5749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1491),
				.a1(P14A1),
				.a2(P14B1),
				.a3(P1591),
				.a4(P15A1),
				.a5(P15B1),
				.a6(P1691),
				.a7(P16A1),
				.a8(P16B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11497)
);

ninexnine_unit ninexnine_unit_5750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1492),
				.a1(P14A2),
				.a2(P14B2),
				.a3(P1592),
				.a4(P15A2),
				.a5(P15B2),
				.a6(P1692),
				.a7(P16A2),
				.a8(P16B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12497)
);

ninexnine_unit ninexnine_unit_5751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1493),
				.a1(P14A3),
				.a2(P14B3),
				.a3(P1593),
				.a4(P15A3),
				.a5(P15B3),
				.a6(P1693),
				.a7(P16A3),
				.a8(P16B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13497)
);

assign C1497=c10497+c11497+c12497+c13497;
assign A1497=(C1497>=0)?1:0;

ninexnine_unit ninexnine_unit_5752(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A0),
				.a1(P14B0),
				.a2(P14C0),
				.a3(P15A0),
				.a4(P15B0),
				.a5(P15C0),
				.a6(P16A0),
				.a7(P16B0),
				.a8(P16C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c104A7)
);

ninexnine_unit ninexnine_unit_5753(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A1),
				.a1(P14B1),
				.a2(P14C1),
				.a3(P15A1),
				.a4(P15B1),
				.a5(P15C1),
				.a6(P16A1),
				.a7(P16B1),
				.a8(P16C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c114A7)
);

ninexnine_unit ninexnine_unit_5754(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A2),
				.a1(P14B2),
				.a2(P14C2),
				.a3(P15A2),
				.a4(P15B2),
				.a5(P15C2),
				.a6(P16A2),
				.a7(P16B2),
				.a8(P16C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c124A7)
);

ninexnine_unit ninexnine_unit_5755(
				.clk(clk),
				.rstn(rstn),
				.a0(P14A3),
				.a1(P14B3),
				.a2(P14C3),
				.a3(P15A3),
				.a4(P15B3),
				.a5(P15C3),
				.a6(P16A3),
				.a7(P16B3),
				.a8(P16C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c134A7)
);

assign C14A7=c104A7+c114A7+c124A7+c134A7;
assign A14A7=(C14A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5756(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B0),
				.a1(P14C0),
				.a2(P14D0),
				.a3(P15B0),
				.a4(P15C0),
				.a5(P15D0),
				.a6(P16B0),
				.a7(P16C0),
				.a8(P16D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c104B7)
);

ninexnine_unit ninexnine_unit_5757(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B1),
				.a1(P14C1),
				.a2(P14D1),
				.a3(P15B1),
				.a4(P15C1),
				.a5(P15D1),
				.a6(P16B1),
				.a7(P16C1),
				.a8(P16D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c114B7)
);

ninexnine_unit ninexnine_unit_5758(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B2),
				.a1(P14C2),
				.a2(P14D2),
				.a3(P15B2),
				.a4(P15C2),
				.a5(P15D2),
				.a6(P16B2),
				.a7(P16C2),
				.a8(P16D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c124B7)
);

ninexnine_unit ninexnine_unit_5759(
				.clk(clk),
				.rstn(rstn),
				.a0(P14B3),
				.a1(P14C3),
				.a2(P14D3),
				.a3(P15B3),
				.a4(P15C3),
				.a5(P15D3),
				.a6(P16B3),
				.a7(P16C3),
				.a8(P16D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c134B7)
);

assign C14B7=c104B7+c114B7+c124B7+c134B7;
assign A14B7=(C14B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5760(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C0),
				.a1(P14D0),
				.a2(P14E0),
				.a3(P15C0),
				.a4(P15D0),
				.a5(P15E0),
				.a6(P16C0),
				.a7(P16D0),
				.a8(P16E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c104C7)
);

ninexnine_unit ninexnine_unit_5761(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C1),
				.a1(P14D1),
				.a2(P14E1),
				.a3(P15C1),
				.a4(P15D1),
				.a5(P15E1),
				.a6(P16C1),
				.a7(P16D1),
				.a8(P16E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c114C7)
);

ninexnine_unit ninexnine_unit_5762(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C2),
				.a1(P14D2),
				.a2(P14E2),
				.a3(P15C2),
				.a4(P15D2),
				.a5(P15E2),
				.a6(P16C2),
				.a7(P16D2),
				.a8(P16E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c124C7)
);

ninexnine_unit ninexnine_unit_5763(
				.clk(clk),
				.rstn(rstn),
				.a0(P14C3),
				.a1(P14D3),
				.a2(P14E3),
				.a3(P15C3),
				.a4(P15D3),
				.a5(P15E3),
				.a6(P16C3),
				.a7(P16D3),
				.a8(P16E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c134C7)
);

assign C14C7=c104C7+c114C7+c124C7+c134C7;
assign A14C7=(C14C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5764(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D0),
				.a1(P14E0),
				.a2(P14F0),
				.a3(P15D0),
				.a4(P15E0),
				.a5(P15F0),
				.a6(P16D0),
				.a7(P16E0),
				.a8(P16F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c104D7)
);

ninexnine_unit ninexnine_unit_5765(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D1),
				.a1(P14E1),
				.a2(P14F1),
				.a3(P15D1),
				.a4(P15E1),
				.a5(P15F1),
				.a6(P16D1),
				.a7(P16E1),
				.a8(P16F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c114D7)
);

ninexnine_unit ninexnine_unit_5766(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D2),
				.a1(P14E2),
				.a2(P14F2),
				.a3(P15D2),
				.a4(P15E2),
				.a5(P15F2),
				.a6(P16D2),
				.a7(P16E2),
				.a8(P16F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c124D7)
);

ninexnine_unit ninexnine_unit_5767(
				.clk(clk),
				.rstn(rstn),
				.a0(P14D3),
				.a1(P14E3),
				.a2(P14F3),
				.a3(P15D3),
				.a4(P15E3),
				.a5(P15F3),
				.a6(P16D3),
				.a7(P16E3),
				.a8(P16F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c134D7)
);

assign C14D7=c104D7+c114D7+c124D7+c134D7;
assign A14D7=(C14D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1500),
				.a1(P1510),
				.a2(P1520),
				.a3(P1600),
				.a4(P1610),
				.a5(P1620),
				.a6(P1700),
				.a7(P1710),
				.a8(P1720),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10507)
);

ninexnine_unit ninexnine_unit_5769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1501),
				.a1(P1511),
				.a2(P1521),
				.a3(P1601),
				.a4(P1611),
				.a5(P1621),
				.a6(P1701),
				.a7(P1711),
				.a8(P1721),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11507)
);

ninexnine_unit ninexnine_unit_5770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1502),
				.a1(P1512),
				.a2(P1522),
				.a3(P1602),
				.a4(P1612),
				.a5(P1622),
				.a6(P1702),
				.a7(P1712),
				.a8(P1722),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12507)
);

ninexnine_unit ninexnine_unit_5771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1503),
				.a1(P1513),
				.a2(P1523),
				.a3(P1603),
				.a4(P1613),
				.a5(P1623),
				.a6(P1703),
				.a7(P1713),
				.a8(P1723),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13507)
);

assign C1507=c10507+c11507+c12507+c13507;
assign A1507=(C1507>=0)?1:0;

ninexnine_unit ninexnine_unit_5772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1510),
				.a1(P1520),
				.a2(P1530),
				.a3(P1610),
				.a4(P1620),
				.a5(P1630),
				.a6(P1710),
				.a7(P1720),
				.a8(P1730),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10517)
);

ninexnine_unit ninexnine_unit_5773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1511),
				.a1(P1521),
				.a2(P1531),
				.a3(P1611),
				.a4(P1621),
				.a5(P1631),
				.a6(P1711),
				.a7(P1721),
				.a8(P1731),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11517)
);

ninexnine_unit ninexnine_unit_5774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1512),
				.a1(P1522),
				.a2(P1532),
				.a3(P1612),
				.a4(P1622),
				.a5(P1632),
				.a6(P1712),
				.a7(P1722),
				.a8(P1732),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12517)
);

ninexnine_unit ninexnine_unit_5775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1513),
				.a1(P1523),
				.a2(P1533),
				.a3(P1613),
				.a4(P1623),
				.a5(P1633),
				.a6(P1713),
				.a7(P1723),
				.a8(P1733),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13517)
);

assign C1517=c10517+c11517+c12517+c13517;
assign A1517=(C1517>=0)?1:0;

ninexnine_unit ninexnine_unit_5776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1520),
				.a1(P1530),
				.a2(P1540),
				.a3(P1620),
				.a4(P1630),
				.a5(P1640),
				.a6(P1720),
				.a7(P1730),
				.a8(P1740),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10527)
);

ninexnine_unit ninexnine_unit_5777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1521),
				.a1(P1531),
				.a2(P1541),
				.a3(P1621),
				.a4(P1631),
				.a5(P1641),
				.a6(P1721),
				.a7(P1731),
				.a8(P1741),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11527)
);

ninexnine_unit ninexnine_unit_5778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1522),
				.a1(P1532),
				.a2(P1542),
				.a3(P1622),
				.a4(P1632),
				.a5(P1642),
				.a6(P1722),
				.a7(P1732),
				.a8(P1742),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12527)
);

ninexnine_unit ninexnine_unit_5779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1523),
				.a1(P1533),
				.a2(P1543),
				.a3(P1623),
				.a4(P1633),
				.a5(P1643),
				.a6(P1723),
				.a7(P1733),
				.a8(P1743),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13527)
);

assign C1527=c10527+c11527+c12527+c13527;
assign A1527=(C1527>=0)?1:0;

ninexnine_unit ninexnine_unit_5780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1530),
				.a1(P1540),
				.a2(P1550),
				.a3(P1630),
				.a4(P1640),
				.a5(P1650),
				.a6(P1730),
				.a7(P1740),
				.a8(P1750),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10537)
);

ninexnine_unit ninexnine_unit_5781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1531),
				.a1(P1541),
				.a2(P1551),
				.a3(P1631),
				.a4(P1641),
				.a5(P1651),
				.a6(P1731),
				.a7(P1741),
				.a8(P1751),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11537)
);

ninexnine_unit ninexnine_unit_5782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1532),
				.a1(P1542),
				.a2(P1552),
				.a3(P1632),
				.a4(P1642),
				.a5(P1652),
				.a6(P1732),
				.a7(P1742),
				.a8(P1752),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12537)
);

ninexnine_unit ninexnine_unit_5783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1533),
				.a1(P1543),
				.a2(P1553),
				.a3(P1633),
				.a4(P1643),
				.a5(P1653),
				.a6(P1733),
				.a7(P1743),
				.a8(P1753),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13537)
);

assign C1537=c10537+c11537+c12537+c13537;
assign A1537=(C1537>=0)?1:0;

ninexnine_unit ninexnine_unit_5784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1540),
				.a1(P1550),
				.a2(P1560),
				.a3(P1640),
				.a4(P1650),
				.a5(P1660),
				.a6(P1740),
				.a7(P1750),
				.a8(P1760),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10547)
);

ninexnine_unit ninexnine_unit_5785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1541),
				.a1(P1551),
				.a2(P1561),
				.a3(P1641),
				.a4(P1651),
				.a5(P1661),
				.a6(P1741),
				.a7(P1751),
				.a8(P1761),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11547)
);

ninexnine_unit ninexnine_unit_5786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1542),
				.a1(P1552),
				.a2(P1562),
				.a3(P1642),
				.a4(P1652),
				.a5(P1662),
				.a6(P1742),
				.a7(P1752),
				.a8(P1762),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12547)
);

ninexnine_unit ninexnine_unit_5787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1543),
				.a1(P1553),
				.a2(P1563),
				.a3(P1643),
				.a4(P1653),
				.a5(P1663),
				.a6(P1743),
				.a7(P1753),
				.a8(P1763),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13547)
);

assign C1547=c10547+c11547+c12547+c13547;
assign A1547=(C1547>=0)?1:0;

ninexnine_unit ninexnine_unit_5788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1550),
				.a1(P1560),
				.a2(P1570),
				.a3(P1650),
				.a4(P1660),
				.a5(P1670),
				.a6(P1750),
				.a7(P1760),
				.a8(P1770),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10557)
);

ninexnine_unit ninexnine_unit_5789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1551),
				.a1(P1561),
				.a2(P1571),
				.a3(P1651),
				.a4(P1661),
				.a5(P1671),
				.a6(P1751),
				.a7(P1761),
				.a8(P1771),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11557)
);

ninexnine_unit ninexnine_unit_5790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1552),
				.a1(P1562),
				.a2(P1572),
				.a3(P1652),
				.a4(P1662),
				.a5(P1672),
				.a6(P1752),
				.a7(P1762),
				.a8(P1772),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12557)
);

ninexnine_unit ninexnine_unit_5791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1553),
				.a1(P1563),
				.a2(P1573),
				.a3(P1653),
				.a4(P1663),
				.a5(P1673),
				.a6(P1753),
				.a7(P1763),
				.a8(P1773),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13557)
);

assign C1557=c10557+c11557+c12557+c13557;
assign A1557=(C1557>=0)?1:0;

ninexnine_unit ninexnine_unit_5792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1560),
				.a1(P1570),
				.a2(P1580),
				.a3(P1660),
				.a4(P1670),
				.a5(P1680),
				.a6(P1760),
				.a7(P1770),
				.a8(P1780),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10567)
);

ninexnine_unit ninexnine_unit_5793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1561),
				.a1(P1571),
				.a2(P1581),
				.a3(P1661),
				.a4(P1671),
				.a5(P1681),
				.a6(P1761),
				.a7(P1771),
				.a8(P1781),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11567)
);

ninexnine_unit ninexnine_unit_5794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1562),
				.a1(P1572),
				.a2(P1582),
				.a3(P1662),
				.a4(P1672),
				.a5(P1682),
				.a6(P1762),
				.a7(P1772),
				.a8(P1782),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12567)
);

ninexnine_unit ninexnine_unit_5795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1563),
				.a1(P1573),
				.a2(P1583),
				.a3(P1663),
				.a4(P1673),
				.a5(P1683),
				.a6(P1763),
				.a7(P1773),
				.a8(P1783),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13567)
);

assign C1567=c10567+c11567+c12567+c13567;
assign A1567=(C1567>=0)?1:0;

ninexnine_unit ninexnine_unit_5796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1570),
				.a1(P1580),
				.a2(P1590),
				.a3(P1670),
				.a4(P1680),
				.a5(P1690),
				.a6(P1770),
				.a7(P1780),
				.a8(P1790),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10577)
);

ninexnine_unit ninexnine_unit_5797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1571),
				.a1(P1581),
				.a2(P1591),
				.a3(P1671),
				.a4(P1681),
				.a5(P1691),
				.a6(P1771),
				.a7(P1781),
				.a8(P1791),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11577)
);

ninexnine_unit ninexnine_unit_5798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1572),
				.a1(P1582),
				.a2(P1592),
				.a3(P1672),
				.a4(P1682),
				.a5(P1692),
				.a6(P1772),
				.a7(P1782),
				.a8(P1792),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12577)
);

ninexnine_unit ninexnine_unit_5799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1573),
				.a1(P1583),
				.a2(P1593),
				.a3(P1673),
				.a4(P1683),
				.a5(P1693),
				.a6(P1773),
				.a7(P1783),
				.a8(P1793),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13577)
);

assign C1577=c10577+c11577+c12577+c13577;
assign A1577=(C1577>=0)?1:0;

ninexnine_unit ninexnine_unit_5800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1580),
				.a1(P1590),
				.a2(P15A0),
				.a3(P1680),
				.a4(P1690),
				.a5(P16A0),
				.a6(P1780),
				.a7(P1790),
				.a8(P17A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10587)
);

ninexnine_unit ninexnine_unit_5801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1581),
				.a1(P1591),
				.a2(P15A1),
				.a3(P1681),
				.a4(P1691),
				.a5(P16A1),
				.a6(P1781),
				.a7(P1791),
				.a8(P17A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11587)
);

ninexnine_unit ninexnine_unit_5802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1582),
				.a1(P1592),
				.a2(P15A2),
				.a3(P1682),
				.a4(P1692),
				.a5(P16A2),
				.a6(P1782),
				.a7(P1792),
				.a8(P17A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12587)
);

ninexnine_unit ninexnine_unit_5803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1583),
				.a1(P1593),
				.a2(P15A3),
				.a3(P1683),
				.a4(P1693),
				.a5(P16A3),
				.a6(P1783),
				.a7(P1793),
				.a8(P17A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13587)
);

assign C1587=c10587+c11587+c12587+c13587;
assign A1587=(C1587>=0)?1:0;

ninexnine_unit ninexnine_unit_5804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1590),
				.a1(P15A0),
				.a2(P15B0),
				.a3(P1690),
				.a4(P16A0),
				.a5(P16B0),
				.a6(P1790),
				.a7(P17A0),
				.a8(P17B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10597)
);

ninexnine_unit ninexnine_unit_5805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1591),
				.a1(P15A1),
				.a2(P15B1),
				.a3(P1691),
				.a4(P16A1),
				.a5(P16B1),
				.a6(P1791),
				.a7(P17A1),
				.a8(P17B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11597)
);

ninexnine_unit ninexnine_unit_5806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1592),
				.a1(P15A2),
				.a2(P15B2),
				.a3(P1692),
				.a4(P16A2),
				.a5(P16B2),
				.a6(P1792),
				.a7(P17A2),
				.a8(P17B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12597)
);

ninexnine_unit ninexnine_unit_5807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1593),
				.a1(P15A3),
				.a2(P15B3),
				.a3(P1693),
				.a4(P16A3),
				.a5(P16B3),
				.a6(P1793),
				.a7(P17A3),
				.a8(P17B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13597)
);

assign C1597=c10597+c11597+c12597+c13597;
assign A1597=(C1597>=0)?1:0;

ninexnine_unit ninexnine_unit_5808(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A0),
				.a1(P15B0),
				.a2(P15C0),
				.a3(P16A0),
				.a4(P16B0),
				.a5(P16C0),
				.a6(P17A0),
				.a7(P17B0),
				.a8(P17C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c105A7)
);

ninexnine_unit ninexnine_unit_5809(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A1),
				.a1(P15B1),
				.a2(P15C1),
				.a3(P16A1),
				.a4(P16B1),
				.a5(P16C1),
				.a6(P17A1),
				.a7(P17B1),
				.a8(P17C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c115A7)
);

ninexnine_unit ninexnine_unit_5810(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A2),
				.a1(P15B2),
				.a2(P15C2),
				.a3(P16A2),
				.a4(P16B2),
				.a5(P16C2),
				.a6(P17A2),
				.a7(P17B2),
				.a8(P17C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c125A7)
);

ninexnine_unit ninexnine_unit_5811(
				.clk(clk),
				.rstn(rstn),
				.a0(P15A3),
				.a1(P15B3),
				.a2(P15C3),
				.a3(P16A3),
				.a4(P16B3),
				.a5(P16C3),
				.a6(P17A3),
				.a7(P17B3),
				.a8(P17C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c135A7)
);

assign C15A7=c105A7+c115A7+c125A7+c135A7;
assign A15A7=(C15A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5812(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B0),
				.a1(P15C0),
				.a2(P15D0),
				.a3(P16B0),
				.a4(P16C0),
				.a5(P16D0),
				.a6(P17B0),
				.a7(P17C0),
				.a8(P17D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c105B7)
);

ninexnine_unit ninexnine_unit_5813(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B1),
				.a1(P15C1),
				.a2(P15D1),
				.a3(P16B1),
				.a4(P16C1),
				.a5(P16D1),
				.a6(P17B1),
				.a7(P17C1),
				.a8(P17D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c115B7)
);

ninexnine_unit ninexnine_unit_5814(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B2),
				.a1(P15C2),
				.a2(P15D2),
				.a3(P16B2),
				.a4(P16C2),
				.a5(P16D2),
				.a6(P17B2),
				.a7(P17C2),
				.a8(P17D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c125B7)
);

ninexnine_unit ninexnine_unit_5815(
				.clk(clk),
				.rstn(rstn),
				.a0(P15B3),
				.a1(P15C3),
				.a2(P15D3),
				.a3(P16B3),
				.a4(P16C3),
				.a5(P16D3),
				.a6(P17B3),
				.a7(P17C3),
				.a8(P17D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c135B7)
);

assign C15B7=c105B7+c115B7+c125B7+c135B7;
assign A15B7=(C15B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5816(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C0),
				.a1(P15D0),
				.a2(P15E0),
				.a3(P16C0),
				.a4(P16D0),
				.a5(P16E0),
				.a6(P17C0),
				.a7(P17D0),
				.a8(P17E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c105C7)
);

ninexnine_unit ninexnine_unit_5817(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C1),
				.a1(P15D1),
				.a2(P15E1),
				.a3(P16C1),
				.a4(P16D1),
				.a5(P16E1),
				.a6(P17C1),
				.a7(P17D1),
				.a8(P17E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c115C7)
);

ninexnine_unit ninexnine_unit_5818(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C2),
				.a1(P15D2),
				.a2(P15E2),
				.a3(P16C2),
				.a4(P16D2),
				.a5(P16E2),
				.a6(P17C2),
				.a7(P17D2),
				.a8(P17E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c125C7)
);

ninexnine_unit ninexnine_unit_5819(
				.clk(clk),
				.rstn(rstn),
				.a0(P15C3),
				.a1(P15D3),
				.a2(P15E3),
				.a3(P16C3),
				.a4(P16D3),
				.a5(P16E3),
				.a6(P17C3),
				.a7(P17D3),
				.a8(P17E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c135C7)
);

assign C15C7=c105C7+c115C7+c125C7+c135C7;
assign A15C7=(C15C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5820(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D0),
				.a1(P15E0),
				.a2(P15F0),
				.a3(P16D0),
				.a4(P16E0),
				.a5(P16F0),
				.a6(P17D0),
				.a7(P17E0),
				.a8(P17F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c105D7)
);

ninexnine_unit ninexnine_unit_5821(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D1),
				.a1(P15E1),
				.a2(P15F1),
				.a3(P16D1),
				.a4(P16E1),
				.a5(P16F1),
				.a6(P17D1),
				.a7(P17E1),
				.a8(P17F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c115D7)
);

ninexnine_unit ninexnine_unit_5822(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D2),
				.a1(P15E2),
				.a2(P15F2),
				.a3(P16D2),
				.a4(P16E2),
				.a5(P16F2),
				.a6(P17D2),
				.a7(P17E2),
				.a8(P17F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c125D7)
);

ninexnine_unit ninexnine_unit_5823(
				.clk(clk),
				.rstn(rstn),
				.a0(P15D3),
				.a1(P15E3),
				.a2(P15F3),
				.a3(P16D3),
				.a4(P16E3),
				.a5(P16F3),
				.a6(P17D3),
				.a7(P17E3),
				.a8(P17F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c135D7)
);

assign C15D7=c105D7+c115D7+c125D7+c135D7;
assign A15D7=(C15D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1600),
				.a1(P1610),
				.a2(P1620),
				.a3(P1700),
				.a4(P1710),
				.a5(P1720),
				.a6(P1800),
				.a7(P1810),
				.a8(P1820),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10607)
);

ninexnine_unit ninexnine_unit_5825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1601),
				.a1(P1611),
				.a2(P1621),
				.a3(P1701),
				.a4(P1711),
				.a5(P1721),
				.a6(P1801),
				.a7(P1811),
				.a8(P1821),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11607)
);

ninexnine_unit ninexnine_unit_5826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1602),
				.a1(P1612),
				.a2(P1622),
				.a3(P1702),
				.a4(P1712),
				.a5(P1722),
				.a6(P1802),
				.a7(P1812),
				.a8(P1822),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12607)
);

ninexnine_unit ninexnine_unit_5827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1603),
				.a1(P1613),
				.a2(P1623),
				.a3(P1703),
				.a4(P1713),
				.a5(P1723),
				.a6(P1803),
				.a7(P1813),
				.a8(P1823),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13607)
);

assign C1607=c10607+c11607+c12607+c13607;
assign A1607=(C1607>=0)?1:0;

ninexnine_unit ninexnine_unit_5828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1610),
				.a1(P1620),
				.a2(P1630),
				.a3(P1710),
				.a4(P1720),
				.a5(P1730),
				.a6(P1810),
				.a7(P1820),
				.a8(P1830),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10617)
);

ninexnine_unit ninexnine_unit_5829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1611),
				.a1(P1621),
				.a2(P1631),
				.a3(P1711),
				.a4(P1721),
				.a5(P1731),
				.a6(P1811),
				.a7(P1821),
				.a8(P1831),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11617)
);

ninexnine_unit ninexnine_unit_5830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1612),
				.a1(P1622),
				.a2(P1632),
				.a3(P1712),
				.a4(P1722),
				.a5(P1732),
				.a6(P1812),
				.a7(P1822),
				.a8(P1832),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12617)
);

ninexnine_unit ninexnine_unit_5831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1613),
				.a1(P1623),
				.a2(P1633),
				.a3(P1713),
				.a4(P1723),
				.a5(P1733),
				.a6(P1813),
				.a7(P1823),
				.a8(P1833),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13617)
);

assign C1617=c10617+c11617+c12617+c13617;
assign A1617=(C1617>=0)?1:0;

ninexnine_unit ninexnine_unit_5832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1620),
				.a1(P1630),
				.a2(P1640),
				.a3(P1720),
				.a4(P1730),
				.a5(P1740),
				.a6(P1820),
				.a7(P1830),
				.a8(P1840),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10627)
);

ninexnine_unit ninexnine_unit_5833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1621),
				.a1(P1631),
				.a2(P1641),
				.a3(P1721),
				.a4(P1731),
				.a5(P1741),
				.a6(P1821),
				.a7(P1831),
				.a8(P1841),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11627)
);

ninexnine_unit ninexnine_unit_5834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1622),
				.a1(P1632),
				.a2(P1642),
				.a3(P1722),
				.a4(P1732),
				.a5(P1742),
				.a6(P1822),
				.a7(P1832),
				.a8(P1842),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12627)
);

ninexnine_unit ninexnine_unit_5835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1623),
				.a1(P1633),
				.a2(P1643),
				.a3(P1723),
				.a4(P1733),
				.a5(P1743),
				.a6(P1823),
				.a7(P1833),
				.a8(P1843),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13627)
);

assign C1627=c10627+c11627+c12627+c13627;
assign A1627=(C1627>=0)?1:0;

ninexnine_unit ninexnine_unit_5836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1630),
				.a1(P1640),
				.a2(P1650),
				.a3(P1730),
				.a4(P1740),
				.a5(P1750),
				.a6(P1830),
				.a7(P1840),
				.a8(P1850),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10637)
);

ninexnine_unit ninexnine_unit_5837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1631),
				.a1(P1641),
				.a2(P1651),
				.a3(P1731),
				.a4(P1741),
				.a5(P1751),
				.a6(P1831),
				.a7(P1841),
				.a8(P1851),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11637)
);

ninexnine_unit ninexnine_unit_5838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1632),
				.a1(P1642),
				.a2(P1652),
				.a3(P1732),
				.a4(P1742),
				.a5(P1752),
				.a6(P1832),
				.a7(P1842),
				.a8(P1852),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12637)
);

ninexnine_unit ninexnine_unit_5839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1633),
				.a1(P1643),
				.a2(P1653),
				.a3(P1733),
				.a4(P1743),
				.a5(P1753),
				.a6(P1833),
				.a7(P1843),
				.a8(P1853),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13637)
);

assign C1637=c10637+c11637+c12637+c13637;
assign A1637=(C1637>=0)?1:0;

ninexnine_unit ninexnine_unit_5840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1640),
				.a1(P1650),
				.a2(P1660),
				.a3(P1740),
				.a4(P1750),
				.a5(P1760),
				.a6(P1840),
				.a7(P1850),
				.a8(P1860),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10647)
);

ninexnine_unit ninexnine_unit_5841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1641),
				.a1(P1651),
				.a2(P1661),
				.a3(P1741),
				.a4(P1751),
				.a5(P1761),
				.a6(P1841),
				.a7(P1851),
				.a8(P1861),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11647)
);

ninexnine_unit ninexnine_unit_5842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1642),
				.a1(P1652),
				.a2(P1662),
				.a3(P1742),
				.a4(P1752),
				.a5(P1762),
				.a6(P1842),
				.a7(P1852),
				.a8(P1862),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12647)
);

ninexnine_unit ninexnine_unit_5843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1643),
				.a1(P1653),
				.a2(P1663),
				.a3(P1743),
				.a4(P1753),
				.a5(P1763),
				.a6(P1843),
				.a7(P1853),
				.a8(P1863),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13647)
);

assign C1647=c10647+c11647+c12647+c13647;
assign A1647=(C1647>=0)?1:0;

ninexnine_unit ninexnine_unit_5844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1650),
				.a1(P1660),
				.a2(P1670),
				.a3(P1750),
				.a4(P1760),
				.a5(P1770),
				.a6(P1850),
				.a7(P1860),
				.a8(P1870),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10657)
);

ninexnine_unit ninexnine_unit_5845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1651),
				.a1(P1661),
				.a2(P1671),
				.a3(P1751),
				.a4(P1761),
				.a5(P1771),
				.a6(P1851),
				.a7(P1861),
				.a8(P1871),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11657)
);

ninexnine_unit ninexnine_unit_5846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1652),
				.a1(P1662),
				.a2(P1672),
				.a3(P1752),
				.a4(P1762),
				.a5(P1772),
				.a6(P1852),
				.a7(P1862),
				.a8(P1872),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12657)
);

ninexnine_unit ninexnine_unit_5847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1653),
				.a1(P1663),
				.a2(P1673),
				.a3(P1753),
				.a4(P1763),
				.a5(P1773),
				.a6(P1853),
				.a7(P1863),
				.a8(P1873),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13657)
);

assign C1657=c10657+c11657+c12657+c13657;
assign A1657=(C1657>=0)?1:0;

ninexnine_unit ninexnine_unit_5848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1660),
				.a1(P1670),
				.a2(P1680),
				.a3(P1760),
				.a4(P1770),
				.a5(P1780),
				.a6(P1860),
				.a7(P1870),
				.a8(P1880),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10667)
);

ninexnine_unit ninexnine_unit_5849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1661),
				.a1(P1671),
				.a2(P1681),
				.a3(P1761),
				.a4(P1771),
				.a5(P1781),
				.a6(P1861),
				.a7(P1871),
				.a8(P1881),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11667)
);

ninexnine_unit ninexnine_unit_5850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1662),
				.a1(P1672),
				.a2(P1682),
				.a3(P1762),
				.a4(P1772),
				.a5(P1782),
				.a6(P1862),
				.a7(P1872),
				.a8(P1882),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12667)
);

ninexnine_unit ninexnine_unit_5851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1663),
				.a1(P1673),
				.a2(P1683),
				.a3(P1763),
				.a4(P1773),
				.a5(P1783),
				.a6(P1863),
				.a7(P1873),
				.a8(P1883),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13667)
);

assign C1667=c10667+c11667+c12667+c13667;
assign A1667=(C1667>=0)?1:0;

ninexnine_unit ninexnine_unit_5852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1670),
				.a1(P1680),
				.a2(P1690),
				.a3(P1770),
				.a4(P1780),
				.a5(P1790),
				.a6(P1870),
				.a7(P1880),
				.a8(P1890),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10677)
);

ninexnine_unit ninexnine_unit_5853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1671),
				.a1(P1681),
				.a2(P1691),
				.a3(P1771),
				.a4(P1781),
				.a5(P1791),
				.a6(P1871),
				.a7(P1881),
				.a8(P1891),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11677)
);

ninexnine_unit ninexnine_unit_5854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1672),
				.a1(P1682),
				.a2(P1692),
				.a3(P1772),
				.a4(P1782),
				.a5(P1792),
				.a6(P1872),
				.a7(P1882),
				.a8(P1892),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12677)
);

ninexnine_unit ninexnine_unit_5855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1673),
				.a1(P1683),
				.a2(P1693),
				.a3(P1773),
				.a4(P1783),
				.a5(P1793),
				.a6(P1873),
				.a7(P1883),
				.a8(P1893),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13677)
);

assign C1677=c10677+c11677+c12677+c13677;
assign A1677=(C1677>=0)?1:0;

ninexnine_unit ninexnine_unit_5856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1680),
				.a1(P1690),
				.a2(P16A0),
				.a3(P1780),
				.a4(P1790),
				.a5(P17A0),
				.a6(P1880),
				.a7(P1890),
				.a8(P18A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10687)
);

ninexnine_unit ninexnine_unit_5857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1681),
				.a1(P1691),
				.a2(P16A1),
				.a3(P1781),
				.a4(P1791),
				.a5(P17A1),
				.a6(P1881),
				.a7(P1891),
				.a8(P18A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11687)
);

ninexnine_unit ninexnine_unit_5858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1682),
				.a1(P1692),
				.a2(P16A2),
				.a3(P1782),
				.a4(P1792),
				.a5(P17A2),
				.a6(P1882),
				.a7(P1892),
				.a8(P18A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12687)
);

ninexnine_unit ninexnine_unit_5859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1683),
				.a1(P1693),
				.a2(P16A3),
				.a3(P1783),
				.a4(P1793),
				.a5(P17A3),
				.a6(P1883),
				.a7(P1893),
				.a8(P18A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13687)
);

assign C1687=c10687+c11687+c12687+c13687;
assign A1687=(C1687>=0)?1:0;

ninexnine_unit ninexnine_unit_5860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1690),
				.a1(P16A0),
				.a2(P16B0),
				.a3(P1790),
				.a4(P17A0),
				.a5(P17B0),
				.a6(P1890),
				.a7(P18A0),
				.a8(P18B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10697)
);

ninexnine_unit ninexnine_unit_5861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1691),
				.a1(P16A1),
				.a2(P16B1),
				.a3(P1791),
				.a4(P17A1),
				.a5(P17B1),
				.a6(P1891),
				.a7(P18A1),
				.a8(P18B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11697)
);

ninexnine_unit ninexnine_unit_5862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1692),
				.a1(P16A2),
				.a2(P16B2),
				.a3(P1792),
				.a4(P17A2),
				.a5(P17B2),
				.a6(P1892),
				.a7(P18A2),
				.a8(P18B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12697)
);

ninexnine_unit ninexnine_unit_5863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1693),
				.a1(P16A3),
				.a2(P16B3),
				.a3(P1793),
				.a4(P17A3),
				.a5(P17B3),
				.a6(P1893),
				.a7(P18A3),
				.a8(P18B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13697)
);

assign C1697=c10697+c11697+c12697+c13697;
assign A1697=(C1697>=0)?1:0;

ninexnine_unit ninexnine_unit_5864(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A0),
				.a1(P16B0),
				.a2(P16C0),
				.a3(P17A0),
				.a4(P17B0),
				.a5(P17C0),
				.a6(P18A0),
				.a7(P18B0),
				.a8(P18C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c106A7)
);

ninexnine_unit ninexnine_unit_5865(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A1),
				.a1(P16B1),
				.a2(P16C1),
				.a3(P17A1),
				.a4(P17B1),
				.a5(P17C1),
				.a6(P18A1),
				.a7(P18B1),
				.a8(P18C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c116A7)
);

ninexnine_unit ninexnine_unit_5866(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A2),
				.a1(P16B2),
				.a2(P16C2),
				.a3(P17A2),
				.a4(P17B2),
				.a5(P17C2),
				.a6(P18A2),
				.a7(P18B2),
				.a8(P18C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c126A7)
);

ninexnine_unit ninexnine_unit_5867(
				.clk(clk),
				.rstn(rstn),
				.a0(P16A3),
				.a1(P16B3),
				.a2(P16C3),
				.a3(P17A3),
				.a4(P17B3),
				.a5(P17C3),
				.a6(P18A3),
				.a7(P18B3),
				.a8(P18C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c136A7)
);

assign C16A7=c106A7+c116A7+c126A7+c136A7;
assign A16A7=(C16A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5868(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B0),
				.a1(P16C0),
				.a2(P16D0),
				.a3(P17B0),
				.a4(P17C0),
				.a5(P17D0),
				.a6(P18B0),
				.a7(P18C0),
				.a8(P18D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c106B7)
);

ninexnine_unit ninexnine_unit_5869(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B1),
				.a1(P16C1),
				.a2(P16D1),
				.a3(P17B1),
				.a4(P17C1),
				.a5(P17D1),
				.a6(P18B1),
				.a7(P18C1),
				.a8(P18D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c116B7)
);

ninexnine_unit ninexnine_unit_5870(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B2),
				.a1(P16C2),
				.a2(P16D2),
				.a3(P17B2),
				.a4(P17C2),
				.a5(P17D2),
				.a6(P18B2),
				.a7(P18C2),
				.a8(P18D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c126B7)
);

ninexnine_unit ninexnine_unit_5871(
				.clk(clk),
				.rstn(rstn),
				.a0(P16B3),
				.a1(P16C3),
				.a2(P16D3),
				.a3(P17B3),
				.a4(P17C3),
				.a5(P17D3),
				.a6(P18B3),
				.a7(P18C3),
				.a8(P18D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c136B7)
);

assign C16B7=c106B7+c116B7+c126B7+c136B7;
assign A16B7=(C16B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5872(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C0),
				.a1(P16D0),
				.a2(P16E0),
				.a3(P17C0),
				.a4(P17D0),
				.a5(P17E0),
				.a6(P18C0),
				.a7(P18D0),
				.a8(P18E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c106C7)
);

ninexnine_unit ninexnine_unit_5873(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C1),
				.a1(P16D1),
				.a2(P16E1),
				.a3(P17C1),
				.a4(P17D1),
				.a5(P17E1),
				.a6(P18C1),
				.a7(P18D1),
				.a8(P18E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c116C7)
);

ninexnine_unit ninexnine_unit_5874(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C2),
				.a1(P16D2),
				.a2(P16E2),
				.a3(P17C2),
				.a4(P17D2),
				.a5(P17E2),
				.a6(P18C2),
				.a7(P18D2),
				.a8(P18E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c126C7)
);

ninexnine_unit ninexnine_unit_5875(
				.clk(clk),
				.rstn(rstn),
				.a0(P16C3),
				.a1(P16D3),
				.a2(P16E3),
				.a3(P17C3),
				.a4(P17D3),
				.a5(P17E3),
				.a6(P18C3),
				.a7(P18D3),
				.a8(P18E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c136C7)
);

assign C16C7=c106C7+c116C7+c126C7+c136C7;
assign A16C7=(C16C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5876(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D0),
				.a1(P16E0),
				.a2(P16F0),
				.a3(P17D0),
				.a4(P17E0),
				.a5(P17F0),
				.a6(P18D0),
				.a7(P18E0),
				.a8(P18F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c106D7)
);

ninexnine_unit ninexnine_unit_5877(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D1),
				.a1(P16E1),
				.a2(P16F1),
				.a3(P17D1),
				.a4(P17E1),
				.a5(P17F1),
				.a6(P18D1),
				.a7(P18E1),
				.a8(P18F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c116D7)
);

ninexnine_unit ninexnine_unit_5878(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D2),
				.a1(P16E2),
				.a2(P16F2),
				.a3(P17D2),
				.a4(P17E2),
				.a5(P17F2),
				.a6(P18D2),
				.a7(P18E2),
				.a8(P18F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c126D7)
);

ninexnine_unit ninexnine_unit_5879(
				.clk(clk),
				.rstn(rstn),
				.a0(P16D3),
				.a1(P16E3),
				.a2(P16F3),
				.a3(P17D3),
				.a4(P17E3),
				.a5(P17F3),
				.a6(P18D3),
				.a7(P18E3),
				.a8(P18F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c136D7)
);

assign C16D7=c106D7+c116D7+c126D7+c136D7;
assign A16D7=(C16D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1700),
				.a1(P1710),
				.a2(P1720),
				.a3(P1800),
				.a4(P1810),
				.a5(P1820),
				.a6(P1900),
				.a7(P1910),
				.a8(P1920),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10707)
);

ninexnine_unit ninexnine_unit_5881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1701),
				.a1(P1711),
				.a2(P1721),
				.a3(P1801),
				.a4(P1811),
				.a5(P1821),
				.a6(P1901),
				.a7(P1911),
				.a8(P1921),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11707)
);

ninexnine_unit ninexnine_unit_5882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1702),
				.a1(P1712),
				.a2(P1722),
				.a3(P1802),
				.a4(P1812),
				.a5(P1822),
				.a6(P1902),
				.a7(P1912),
				.a8(P1922),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12707)
);

ninexnine_unit ninexnine_unit_5883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1703),
				.a1(P1713),
				.a2(P1723),
				.a3(P1803),
				.a4(P1813),
				.a5(P1823),
				.a6(P1903),
				.a7(P1913),
				.a8(P1923),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13707)
);

assign C1707=c10707+c11707+c12707+c13707;
assign A1707=(C1707>=0)?1:0;

ninexnine_unit ninexnine_unit_5884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1710),
				.a1(P1720),
				.a2(P1730),
				.a3(P1810),
				.a4(P1820),
				.a5(P1830),
				.a6(P1910),
				.a7(P1920),
				.a8(P1930),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10717)
);

ninexnine_unit ninexnine_unit_5885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1711),
				.a1(P1721),
				.a2(P1731),
				.a3(P1811),
				.a4(P1821),
				.a5(P1831),
				.a6(P1911),
				.a7(P1921),
				.a8(P1931),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11717)
);

ninexnine_unit ninexnine_unit_5886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1712),
				.a1(P1722),
				.a2(P1732),
				.a3(P1812),
				.a4(P1822),
				.a5(P1832),
				.a6(P1912),
				.a7(P1922),
				.a8(P1932),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12717)
);

ninexnine_unit ninexnine_unit_5887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1713),
				.a1(P1723),
				.a2(P1733),
				.a3(P1813),
				.a4(P1823),
				.a5(P1833),
				.a6(P1913),
				.a7(P1923),
				.a8(P1933),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13717)
);

assign C1717=c10717+c11717+c12717+c13717;
assign A1717=(C1717>=0)?1:0;

ninexnine_unit ninexnine_unit_5888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1720),
				.a1(P1730),
				.a2(P1740),
				.a3(P1820),
				.a4(P1830),
				.a5(P1840),
				.a6(P1920),
				.a7(P1930),
				.a8(P1940),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10727)
);

ninexnine_unit ninexnine_unit_5889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1721),
				.a1(P1731),
				.a2(P1741),
				.a3(P1821),
				.a4(P1831),
				.a5(P1841),
				.a6(P1921),
				.a7(P1931),
				.a8(P1941),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11727)
);

ninexnine_unit ninexnine_unit_5890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1722),
				.a1(P1732),
				.a2(P1742),
				.a3(P1822),
				.a4(P1832),
				.a5(P1842),
				.a6(P1922),
				.a7(P1932),
				.a8(P1942),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12727)
);

ninexnine_unit ninexnine_unit_5891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1723),
				.a1(P1733),
				.a2(P1743),
				.a3(P1823),
				.a4(P1833),
				.a5(P1843),
				.a6(P1923),
				.a7(P1933),
				.a8(P1943),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13727)
);

assign C1727=c10727+c11727+c12727+c13727;
assign A1727=(C1727>=0)?1:0;

ninexnine_unit ninexnine_unit_5892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1730),
				.a1(P1740),
				.a2(P1750),
				.a3(P1830),
				.a4(P1840),
				.a5(P1850),
				.a6(P1930),
				.a7(P1940),
				.a8(P1950),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10737)
);

ninexnine_unit ninexnine_unit_5893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1731),
				.a1(P1741),
				.a2(P1751),
				.a3(P1831),
				.a4(P1841),
				.a5(P1851),
				.a6(P1931),
				.a7(P1941),
				.a8(P1951),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11737)
);

ninexnine_unit ninexnine_unit_5894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1732),
				.a1(P1742),
				.a2(P1752),
				.a3(P1832),
				.a4(P1842),
				.a5(P1852),
				.a6(P1932),
				.a7(P1942),
				.a8(P1952),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12737)
);

ninexnine_unit ninexnine_unit_5895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1733),
				.a1(P1743),
				.a2(P1753),
				.a3(P1833),
				.a4(P1843),
				.a5(P1853),
				.a6(P1933),
				.a7(P1943),
				.a8(P1953),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13737)
);

assign C1737=c10737+c11737+c12737+c13737;
assign A1737=(C1737>=0)?1:0;

ninexnine_unit ninexnine_unit_5896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1740),
				.a1(P1750),
				.a2(P1760),
				.a3(P1840),
				.a4(P1850),
				.a5(P1860),
				.a6(P1940),
				.a7(P1950),
				.a8(P1960),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10747)
);

ninexnine_unit ninexnine_unit_5897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1741),
				.a1(P1751),
				.a2(P1761),
				.a3(P1841),
				.a4(P1851),
				.a5(P1861),
				.a6(P1941),
				.a7(P1951),
				.a8(P1961),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11747)
);

ninexnine_unit ninexnine_unit_5898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1742),
				.a1(P1752),
				.a2(P1762),
				.a3(P1842),
				.a4(P1852),
				.a5(P1862),
				.a6(P1942),
				.a7(P1952),
				.a8(P1962),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12747)
);

ninexnine_unit ninexnine_unit_5899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1743),
				.a1(P1753),
				.a2(P1763),
				.a3(P1843),
				.a4(P1853),
				.a5(P1863),
				.a6(P1943),
				.a7(P1953),
				.a8(P1963),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13747)
);

assign C1747=c10747+c11747+c12747+c13747;
assign A1747=(C1747>=0)?1:0;

ninexnine_unit ninexnine_unit_5900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1750),
				.a1(P1760),
				.a2(P1770),
				.a3(P1850),
				.a4(P1860),
				.a5(P1870),
				.a6(P1950),
				.a7(P1960),
				.a8(P1970),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10757)
);

ninexnine_unit ninexnine_unit_5901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1751),
				.a1(P1761),
				.a2(P1771),
				.a3(P1851),
				.a4(P1861),
				.a5(P1871),
				.a6(P1951),
				.a7(P1961),
				.a8(P1971),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11757)
);

ninexnine_unit ninexnine_unit_5902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1752),
				.a1(P1762),
				.a2(P1772),
				.a3(P1852),
				.a4(P1862),
				.a5(P1872),
				.a6(P1952),
				.a7(P1962),
				.a8(P1972),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12757)
);

ninexnine_unit ninexnine_unit_5903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1753),
				.a1(P1763),
				.a2(P1773),
				.a3(P1853),
				.a4(P1863),
				.a5(P1873),
				.a6(P1953),
				.a7(P1963),
				.a8(P1973),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13757)
);

assign C1757=c10757+c11757+c12757+c13757;
assign A1757=(C1757>=0)?1:0;

ninexnine_unit ninexnine_unit_5904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1760),
				.a1(P1770),
				.a2(P1780),
				.a3(P1860),
				.a4(P1870),
				.a5(P1880),
				.a6(P1960),
				.a7(P1970),
				.a8(P1980),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10767)
);

ninexnine_unit ninexnine_unit_5905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1761),
				.a1(P1771),
				.a2(P1781),
				.a3(P1861),
				.a4(P1871),
				.a5(P1881),
				.a6(P1961),
				.a7(P1971),
				.a8(P1981),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11767)
);

ninexnine_unit ninexnine_unit_5906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1762),
				.a1(P1772),
				.a2(P1782),
				.a3(P1862),
				.a4(P1872),
				.a5(P1882),
				.a6(P1962),
				.a7(P1972),
				.a8(P1982),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12767)
);

ninexnine_unit ninexnine_unit_5907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1763),
				.a1(P1773),
				.a2(P1783),
				.a3(P1863),
				.a4(P1873),
				.a5(P1883),
				.a6(P1963),
				.a7(P1973),
				.a8(P1983),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13767)
);

assign C1767=c10767+c11767+c12767+c13767;
assign A1767=(C1767>=0)?1:0;

ninexnine_unit ninexnine_unit_5908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1770),
				.a1(P1780),
				.a2(P1790),
				.a3(P1870),
				.a4(P1880),
				.a5(P1890),
				.a6(P1970),
				.a7(P1980),
				.a8(P1990),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10777)
);

ninexnine_unit ninexnine_unit_5909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1771),
				.a1(P1781),
				.a2(P1791),
				.a3(P1871),
				.a4(P1881),
				.a5(P1891),
				.a6(P1971),
				.a7(P1981),
				.a8(P1991),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11777)
);

ninexnine_unit ninexnine_unit_5910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1772),
				.a1(P1782),
				.a2(P1792),
				.a3(P1872),
				.a4(P1882),
				.a5(P1892),
				.a6(P1972),
				.a7(P1982),
				.a8(P1992),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12777)
);

ninexnine_unit ninexnine_unit_5911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1773),
				.a1(P1783),
				.a2(P1793),
				.a3(P1873),
				.a4(P1883),
				.a5(P1893),
				.a6(P1973),
				.a7(P1983),
				.a8(P1993),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13777)
);

assign C1777=c10777+c11777+c12777+c13777;
assign A1777=(C1777>=0)?1:0;

ninexnine_unit ninexnine_unit_5912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1780),
				.a1(P1790),
				.a2(P17A0),
				.a3(P1880),
				.a4(P1890),
				.a5(P18A0),
				.a6(P1980),
				.a7(P1990),
				.a8(P19A0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10787)
);

ninexnine_unit ninexnine_unit_5913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1781),
				.a1(P1791),
				.a2(P17A1),
				.a3(P1881),
				.a4(P1891),
				.a5(P18A1),
				.a6(P1981),
				.a7(P1991),
				.a8(P19A1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11787)
);

ninexnine_unit ninexnine_unit_5914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1782),
				.a1(P1792),
				.a2(P17A2),
				.a3(P1882),
				.a4(P1892),
				.a5(P18A2),
				.a6(P1982),
				.a7(P1992),
				.a8(P19A2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12787)
);

ninexnine_unit ninexnine_unit_5915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1783),
				.a1(P1793),
				.a2(P17A3),
				.a3(P1883),
				.a4(P1893),
				.a5(P18A3),
				.a6(P1983),
				.a7(P1993),
				.a8(P19A3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13787)
);

assign C1787=c10787+c11787+c12787+c13787;
assign A1787=(C1787>=0)?1:0;

ninexnine_unit ninexnine_unit_5916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1790),
				.a1(P17A0),
				.a2(P17B0),
				.a3(P1890),
				.a4(P18A0),
				.a5(P18B0),
				.a6(P1990),
				.a7(P19A0),
				.a8(P19B0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10797)
);

ninexnine_unit ninexnine_unit_5917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1791),
				.a1(P17A1),
				.a2(P17B1),
				.a3(P1891),
				.a4(P18A1),
				.a5(P18B1),
				.a6(P1991),
				.a7(P19A1),
				.a8(P19B1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11797)
);

ninexnine_unit ninexnine_unit_5918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1792),
				.a1(P17A2),
				.a2(P17B2),
				.a3(P1892),
				.a4(P18A2),
				.a5(P18B2),
				.a6(P1992),
				.a7(P19A2),
				.a8(P19B2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12797)
);

ninexnine_unit ninexnine_unit_5919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1793),
				.a1(P17A3),
				.a2(P17B3),
				.a3(P1893),
				.a4(P18A3),
				.a5(P18B3),
				.a6(P1993),
				.a7(P19A3),
				.a8(P19B3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13797)
);

assign C1797=c10797+c11797+c12797+c13797;
assign A1797=(C1797>=0)?1:0;

ninexnine_unit ninexnine_unit_5920(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A0),
				.a1(P17B0),
				.a2(P17C0),
				.a3(P18A0),
				.a4(P18B0),
				.a5(P18C0),
				.a6(P19A0),
				.a7(P19B0),
				.a8(P19C0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c107A7)
);

ninexnine_unit ninexnine_unit_5921(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A1),
				.a1(P17B1),
				.a2(P17C1),
				.a3(P18A1),
				.a4(P18B1),
				.a5(P18C1),
				.a6(P19A1),
				.a7(P19B1),
				.a8(P19C1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c117A7)
);

ninexnine_unit ninexnine_unit_5922(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A2),
				.a1(P17B2),
				.a2(P17C2),
				.a3(P18A2),
				.a4(P18B2),
				.a5(P18C2),
				.a6(P19A2),
				.a7(P19B2),
				.a8(P19C2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c127A7)
);

ninexnine_unit ninexnine_unit_5923(
				.clk(clk),
				.rstn(rstn),
				.a0(P17A3),
				.a1(P17B3),
				.a2(P17C3),
				.a3(P18A3),
				.a4(P18B3),
				.a5(P18C3),
				.a6(P19A3),
				.a7(P19B3),
				.a8(P19C3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c137A7)
);

assign C17A7=c107A7+c117A7+c127A7+c137A7;
assign A17A7=(C17A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5924(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B0),
				.a1(P17C0),
				.a2(P17D0),
				.a3(P18B0),
				.a4(P18C0),
				.a5(P18D0),
				.a6(P19B0),
				.a7(P19C0),
				.a8(P19D0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c107B7)
);

ninexnine_unit ninexnine_unit_5925(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B1),
				.a1(P17C1),
				.a2(P17D1),
				.a3(P18B1),
				.a4(P18C1),
				.a5(P18D1),
				.a6(P19B1),
				.a7(P19C1),
				.a8(P19D1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c117B7)
);

ninexnine_unit ninexnine_unit_5926(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B2),
				.a1(P17C2),
				.a2(P17D2),
				.a3(P18B2),
				.a4(P18C2),
				.a5(P18D2),
				.a6(P19B2),
				.a7(P19C2),
				.a8(P19D2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c127B7)
);

ninexnine_unit ninexnine_unit_5927(
				.clk(clk),
				.rstn(rstn),
				.a0(P17B3),
				.a1(P17C3),
				.a2(P17D3),
				.a3(P18B3),
				.a4(P18C3),
				.a5(P18D3),
				.a6(P19B3),
				.a7(P19C3),
				.a8(P19D3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c137B7)
);

assign C17B7=c107B7+c117B7+c127B7+c137B7;
assign A17B7=(C17B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5928(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C0),
				.a1(P17D0),
				.a2(P17E0),
				.a3(P18C0),
				.a4(P18D0),
				.a5(P18E0),
				.a6(P19C0),
				.a7(P19D0),
				.a8(P19E0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c107C7)
);

ninexnine_unit ninexnine_unit_5929(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C1),
				.a1(P17D1),
				.a2(P17E1),
				.a3(P18C1),
				.a4(P18D1),
				.a5(P18E1),
				.a6(P19C1),
				.a7(P19D1),
				.a8(P19E1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c117C7)
);

ninexnine_unit ninexnine_unit_5930(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C2),
				.a1(P17D2),
				.a2(P17E2),
				.a3(P18C2),
				.a4(P18D2),
				.a5(P18E2),
				.a6(P19C2),
				.a7(P19D2),
				.a8(P19E2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c127C7)
);

ninexnine_unit ninexnine_unit_5931(
				.clk(clk),
				.rstn(rstn),
				.a0(P17C3),
				.a1(P17D3),
				.a2(P17E3),
				.a3(P18C3),
				.a4(P18D3),
				.a5(P18E3),
				.a6(P19C3),
				.a7(P19D3),
				.a8(P19E3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c137C7)
);

assign C17C7=c107C7+c117C7+c127C7+c137C7;
assign A17C7=(C17C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5932(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D0),
				.a1(P17E0),
				.a2(P17F0),
				.a3(P18D0),
				.a4(P18E0),
				.a5(P18F0),
				.a6(P19D0),
				.a7(P19E0),
				.a8(P19F0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c107D7)
);

ninexnine_unit ninexnine_unit_5933(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D1),
				.a1(P17E1),
				.a2(P17F1),
				.a3(P18D1),
				.a4(P18E1),
				.a5(P18F1),
				.a6(P19D1),
				.a7(P19E1),
				.a8(P19F1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c117D7)
);

ninexnine_unit ninexnine_unit_5934(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D2),
				.a1(P17E2),
				.a2(P17F2),
				.a3(P18D2),
				.a4(P18E2),
				.a5(P18F2),
				.a6(P19D2),
				.a7(P19E2),
				.a8(P19F2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c127D7)
);

ninexnine_unit ninexnine_unit_5935(
				.clk(clk),
				.rstn(rstn),
				.a0(P17D3),
				.a1(P17E3),
				.a2(P17F3),
				.a3(P18D3),
				.a4(P18E3),
				.a5(P18F3),
				.a6(P19D3),
				.a7(P19E3),
				.a8(P19F3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c137D7)
);

assign C17D7=c107D7+c117D7+c127D7+c137D7;
assign A17D7=(C17D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1800),
				.a1(P1810),
				.a2(P1820),
				.a3(P1900),
				.a4(P1910),
				.a5(P1920),
				.a6(P1A00),
				.a7(P1A10),
				.a8(P1A20),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10807)
);

ninexnine_unit ninexnine_unit_5937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1801),
				.a1(P1811),
				.a2(P1821),
				.a3(P1901),
				.a4(P1911),
				.a5(P1921),
				.a6(P1A01),
				.a7(P1A11),
				.a8(P1A21),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11807)
);

ninexnine_unit ninexnine_unit_5938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1802),
				.a1(P1812),
				.a2(P1822),
				.a3(P1902),
				.a4(P1912),
				.a5(P1922),
				.a6(P1A02),
				.a7(P1A12),
				.a8(P1A22),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12807)
);

ninexnine_unit ninexnine_unit_5939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1803),
				.a1(P1813),
				.a2(P1823),
				.a3(P1903),
				.a4(P1913),
				.a5(P1923),
				.a6(P1A03),
				.a7(P1A13),
				.a8(P1A23),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13807)
);

assign C1807=c10807+c11807+c12807+c13807;
assign A1807=(C1807>=0)?1:0;

ninexnine_unit ninexnine_unit_5940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1810),
				.a1(P1820),
				.a2(P1830),
				.a3(P1910),
				.a4(P1920),
				.a5(P1930),
				.a6(P1A10),
				.a7(P1A20),
				.a8(P1A30),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10817)
);

ninexnine_unit ninexnine_unit_5941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1811),
				.a1(P1821),
				.a2(P1831),
				.a3(P1911),
				.a4(P1921),
				.a5(P1931),
				.a6(P1A11),
				.a7(P1A21),
				.a8(P1A31),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11817)
);

ninexnine_unit ninexnine_unit_5942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1812),
				.a1(P1822),
				.a2(P1832),
				.a3(P1912),
				.a4(P1922),
				.a5(P1932),
				.a6(P1A12),
				.a7(P1A22),
				.a8(P1A32),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12817)
);

ninexnine_unit ninexnine_unit_5943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1813),
				.a1(P1823),
				.a2(P1833),
				.a3(P1913),
				.a4(P1923),
				.a5(P1933),
				.a6(P1A13),
				.a7(P1A23),
				.a8(P1A33),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13817)
);

assign C1817=c10817+c11817+c12817+c13817;
assign A1817=(C1817>=0)?1:0;

ninexnine_unit ninexnine_unit_5944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1820),
				.a1(P1830),
				.a2(P1840),
				.a3(P1920),
				.a4(P1930),
				.a5(P1940),
				.a6(P1A20),
				.a7(P1A30),
				.a8(P1A40),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10827)
);

ninexnine_unit ninexnine_unit_5945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1821),
				.a1(P1831),
				.a2(P1841),
				.a3(P1921),
				.a4(P1931),
				.a5(P1941),
				.a6(P1A21),
				.a7(P1A31),
				.a8(P1A41),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11827)
);

ninexnine_unit ninexnine_unit_5946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1822),
				.a1(P1832),
				.a2(P1842),
				.a3(P1922),
				.a4(P1932),
				.a5(P1942),
				.a6(P1A22),
				.a7(P1A32),
				.a8(P1A42),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12827)
);

ninexnine_unit ninexnine_unit_5947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1823),
				.a1(P1833),
				.a2(P1843),
				.a3(P1923),
				.a4(P1933),
				.a5(P1943),
				.a6(P1A23),
				.a7(P1A33),
				.a8(P1A43),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13827)
);

assign C1827=c10827+c11827+c12827+c13827;
assign A1827=(C1827>=0)?1:0;

ninexnine_unit ninexnine_unit_5948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1830),
				.a1(P1840),
				.a2(P1850),
				.a3(P1930),
				.a4(P1940),
				.a5(P1950),
				.a6(P1A30),
				.a7(P1A40),
				.a8(P1A50),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10837)
);

ninexnine_unit ninexnine_unit_5949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1831),
				.a1(P1841),
				.a2(P1851),
				.a3(P1931),
				.a4(P1941),
				.a5(P1951),
				.a6(P1A31),
				.a7(P1A41),
				.a8(P1A51),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11837)
);

ninexnine_unit ninexnine_unit_5950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1832),
				.a1(P1842),
				.a2(P1852),
				.a3(P1932),
				.a4(P1942),
				.a5(P1952),
				.a6(P1A32),
				.a7(P1A42),
				.a8(P1A52),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12837)
);

ninexnine_unit ninexnine_unit_5951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1833),
				.a1(P1843),
				.a2(P1853),
				.a3(P1933),
				.a4(P1943),
				.a5(P1953),
				.a6(P1A33),
				.a7(P1A43),
				.a8(P1A53),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13837)
);

assign C1837=c10837+c11837+c12837+c13837;
assign A1837=(C1837>=0)?1:0;

ninexnine_unit ninexnine_unit_5952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1840),
				.a1(P1850),
				.a2(P1860),
				.a3(P1940),
				.a4(P1950),
				.a5(P1960),
				.a6(P1A40),
				.a7(P1A50),
				.a8(P1A60),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10847)
);

ninexnine_unit ninexnine_unit_5953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1841),
				.a1(P1851),
				.a2(P1861),
				.a3(P1941),
				.a4(P1951),
				.a5(P1961),
				.a6(P1A41),
				.a7(P1A51),
				.a8(P1A61),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11847)
);

ninexnine_unit ninexnine_unit_5954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1842),
				.a1(P1852),
				.a2(P1862),
				.a3(P1942),
				.a4(P1952),
				.a5(P1962),
				.a6(P1A42),
				.a7(P1A52),
				.a8(P1A62),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12847)
);

ninexnine_unit ninexnine_unit_5955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1843),
				.a1(P1853),
				.a2(P1863),
				.a3(P1943),
				.a4(P1953),
				.a5(P1963),
				.a6(P1A43),
				.a7(P1A53),
				.a8(P1A63),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13847)
);

assign C1847=c10847+c11847+c12847+c13847;
assign A1847=(C1847>=0)?1:0;

ninexnine_unit ninexnine_unit_5956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1850),
				.a1(P1860),
				.a2(P1870),
				.a3(P1950),
				.a4(P1960),
				.a5(P1970),
				.a6(P1A50),
				.a7(P1A60),
				.a8(P1A70),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10857)
);

ninexnine_unit ninexnine_unit_5957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1851),
				.a1(P1861),
				.a2(P1871),
				.a3(P1951),
				.a4(P1961),
				.a5(P1971),
				.a6(P1A51),
				.a7(P1A61),
				.a8(P1A71),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11857)
);

ninexnine_unit ninexnine_unit_5958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1852),
				.a1(P1862),
				.a2(P1872),
				.a3(P1952),
				.a4(P1962),
				.a5(P1972),
				.a6(P1A52),
				.a7(P1A62),
				.a8(P1A72),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12857)
);

ninexnine_unit ninexnine_unit_5959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1853),
				.a1(P1863),
				.a2(P1873),
				.a3(P1953),
				.a4(P1963),
				.a5(P1973),
				.a6(P1A53),
				.a7(P1A63),
				.a8(P1A73),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13857)
);

assign C1857=c10857+c11857+c12857+c13857;
assign A1857=(C1857>=0)?1:0;

ninexnine_unit ninexnine_unit_5960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1860),
				.a1(P1870),
				.a2(P1880),
				.a3(P1960),
				.a4(P1970),
				.a5(P1980),
				.a6(P1A60),
				.a7(P1A70),
				.a8(P1A80),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10867)
);

ninexnine_unit ninexnine_unit_5961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1861),
				.a1(P1871),
				.a2(P1881),
				.a3(P1961),
				.a4(P1971),
				.a5(P1981),
				.a6(P1A61),
				.a7(P1A71),
				.a8(P1A81),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11867)
);

ninexnine_unit ninexnine_unit_5962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1862),
				.a1(P1872),
				.a2(P1882),
				.a3(P1962),
				.a4(P1972),
				.a5(P1982),
				.a6(P1A62),
				.a7(P1A72),
				.a8(P1A82),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12867)
);

ninexnine_unit ninexnine_unit_5963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1863),
				.a1(P1873),
				.a2(P1883),
				.a3(P1963),
				.a4(P1973),
				.a5(P1983),
				.a6(P1A63),
				.a7(P1A73),
				.a8(P1A83),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13867)
);

assign C1867=c10867+c11867+c12867+c13867;
assign A1867=(C1867>=0)?1:0;

ninexnine_unit ninexnine_unit_5964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1870),
				.a1(P1880),
				.a2(P1890),
				.a3(P1970),
				.a4(P1980),
				.a5(P1990),
				.a6(P1A70),
				.a7(P1A80),
				.a8(P1A90),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10877)
);

ninexnine_unit ninexnine_unit_5965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1871),
				.a1(P1881),
				.a2(P1891),
				.a3(P1971),
				.a4(P1981),
				.a5(P1991),
				.a6(P1A71),
				.a7(P1A81),
				.a8(P1A91),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11877)
);

ninexnine_unit ninexnine_unit_5966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1872),
				.a1(P1882),
				.a2(P1892),
				.a3(P1972),
				.a4(P1982),
				.a5(P1992),
				.a6(P1A72),
				.a7(P1A82),
				.a8(P1A92),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12877)
);

ninexnine_unit ninexnine_unit_5967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1873),
				.a1(P1883),
				.a2(P1893),
				.a3(P1973),
				.a4(P1983),
				.a5(P1993),
				.a6(P1A73),
				.a7(P1A83),
				.a8(P1A93),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13877)
);

assign C1877=c10877+c11877+c12877+c13877;
assign A1877=(C1877>=0)?1:0;

ninexnine_unit ninexnine_unit_5968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1880),
				.a1(P1890),
				.a2(P18A0),
				.a3(P1980),
				.a4(P1990),
				.a5(P19A0),
				.a6(P1A80),
				.a7(P1A90),
				.a8(P1AA0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10887)
);

ninexnine_unit ninexnine_unit_5969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1881),
				.a1(P1891),
				.a2(P18A1),
				.a3(P1981),
				.a4(P1991),
				.a5(P19A1),
				.a6(P1A81),
				.a7(P1A91),
				.a8(P1AA1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11887)
);

ninexnine_unit ninexnine_unit_5970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1882),
				.a1(P1892),
				.a2(P18A2),
				.a3(P1982),
				.a4(P1992),
				.a5(P19A2),
				.a6(P1A82),
				.a7(P1A92),
				.a8(P1AA2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12887)
);

ninexnine_unit ninexnine_unit_5971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1883),
				.a1(P1893),
				.a2(P18A3),
				.a3(P1983),
				.a4(P1993),
				.a5(P19A3),
				.a6(P1A83),
				.a7(P1A93),
				.a8(P1AA3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13887)
);

assign C1887=c10887+c11887+c12887+c13887;
assign A1887=(C1887>=0)?1:0;

ninexnine_unit ninexnine_unit_5972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1890),
				.a1(P18A0),
				.a2(P18B0),
				.a3(P1990),
				.a4(P19A0),
				.a5(P19B0),
				.a6(P1A90),
				.a7(P1AA0),
				.a8(P1AB0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10897)
);

ninexnine_unit ninexnine_unit_5973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1891),
				.a1(P18A1),
				.a2(P18B1),
				.a3(P1991),
				.a4(P19A1),
				.a5(P19B1),
				.a6(P1A91),
				.a7(P1AA1),
				.a8(P1AB1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11897)
);

ninexnine_unit ninexnine_unit_5974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1892),
				.a1(P18A2),
				.a2(P18B2),
				.a3(P1992),
				.a4(P19A2),
				.a5(P19B2),
				.a6(P1A92),
				.a7(P1AA2),
				.a8(P1AB2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12897)
);

ninexnine_unit ninexnine_unit_5975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1893),
				.a1(P18A3),
				.a2(P18B3),
				.a3(P1993),
				.a4(P19A3),
				.a5(P19B3),
				.a6(P1A93),
				.a7(P1AA3),
				.a8(P1AB3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13897)
);

assign C1897=c10897+c11897+c12897+c13897;
assign A1897=(C1897>=0)?1:0;

ninexnine_unit ninexnine_unit_5976(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A0),
				.a1(P18B0),
				.a2(P18C0),
				.a3(P19A0),
				.a4(P19B0),
				.a5(P19C0),
				.a6(P1AA0),
				.a7(P1AB0),
				.a8(P1AC0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c108A7)
);

ninexnine_unit ninexnine_unit_5977(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A1),
				.a1(P18B1),
				.a2(P18C1),
				.a3(P19A1),
				.a4(P19B1),
				.a5(P19C1),
				.a6(P1AA1),
				.a7(P1AB1),
				.a8(P1AC1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c118A7)
);

ninexnine_unit ninexnine_unit_5978(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A2),
				.a1(P18B2),
				.a2(P18C2),
				.a3(P19A2),
				.a4(P19B2),
				.a5(P19C2),
				.a6(P1AA2),
				.a7(P1AB2),
				.a8(P1AC2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c128A7)
);

ninexnine_unit ninexnine_unit_5979(
				.clk(clk),
				.rstn(rstn),
				.a0(P18A3),
				.a1(P18B3),
				.a2(P18C3),
				.a3(P19A3),
				.a4(P19B3),
				.a5(P19C3),
				.a6(P1AA3),
				.a7(P1AB3),
				.a8(P1AC3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c138A7)
);

assign C18A7=c108A7+c118A7+c128A7+c138A7;
assign A18A7=(C18A7>=0)?1:0;

ninexnine_unit ninexnine_unit_5980(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B0),
				.a1(P18C0),
				.a2(P18D0),
				.a3(P19B0),
				.a4(P19C0),
				.a5(P19D0),
				.a6(P1AB0),
				.a7(P1AC0),
				.a8(P1AD0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c108B7)
);

ninexnine_unit ninexnine_unit_5981(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B1),
				.a1(P18C1),
				.a2(P18D1),
				.a3(P19B1),
				.a4(P19C1),
				.a5(P19D1),
				.a6(P1AB1),
				.a7(P1AC1),
				.a8(P1AD1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c118B7)
);

ninexnine_unit ninexnine_unit_5982(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B2),
				.a1(P18C2),
				.a2(P18D2),
				.a3(P19B2),
				.a4(P19C2),
				.a5(P19D2),
				.a6(P1AB2),
				.a7(P1AC2),
				.a8(P1AD2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c128B7)
);

ninexnine_unit ninexnine_unit_5983(
				.clk(clk),
				.rstn(rstn),
				.a0(P18B3),
				.a1(P18C3),
				.a2(P18D3),
				.a3(P19B3),
				.a4(P19C3),
				.a5(P19D3),
				.a6(P1AB3),
				.a7(P1AC3),
				.a8(P1AD3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c138B7)
);

assign C18B7=c108B7+c118B7+c128B7+c138B7;
assign A18B7=(C18B7>=0)?1:0;

ninexnine_unit ninexnine_unit_5984(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C0),
				.a1(P18D0),
				.a2(P18E0),
				.a3(P19C0),
				.a4(P19D0),
				.a5(P19E0),
				.a6(P1AC0),
				.a7(P1AD0),
				.a8(P1AE0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c108C7)
);

ninexnine_unit ninexnine_unit_5985(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C1),
				.a1(P18D1),
				.a2(P18E1),
				.a3(P19C1),
				.a4(P19D1),
				.a5(P19E1),
				.a6(P1AC1),
				.a7(P1AD1),
				.a8(P1AE1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c118C7)
);

ninexnine_unit ninexnine_unit_5986(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C2),
				.a1(P18D2),
				.a2(P18E2),
				.a3(P19C2),
				.a4(P19D2),
				.a5(P19E2),
				.a6(P1AC2),
				.a7(P1AD2),
				.a8(P1AE2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c128C7)
);

ninexnine_unit ninexnine_unit_5987(
				.clk(clk),
				.rstn(rstn),
				.a0(P18C3),
				.a1(P18D3),
				.a2(P18E3),
				.a3(P19C3),
				.a4(P19D3),
				.a5(P19E3),
				.a6(P1AC3),
				.a7(P1AD3),
				.a8(P1AE3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c138C7)
);

assign C18C7=c108C7+c118C7+c128C7+c138C7;
assign A18C7=(C18C7>=0)?1:0;

ninexnine_unit ninexnine_unit_5988(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D0),
				.a1(P18E0),
				.a2(P18F0),
				.a3(P19D0),
				.a4(P19E0),
				.a5(P19F0),
				.a6(P1AD0),
				.a7(P1AE0),
				.a8(P1AF0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c108D7)
);

ninexnine_unit ninexnine_unit_5989(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D1),
				.a1(P18E1),
				.a2(P18F1),
				.a3(P19D1),
				.a4(P19E1),
				.a5(P19F1),
				.a6(P1AD1),
				.a7(P1AE1),
				.a8(P1AF1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c118D7)
);

ninexnine_unit ninexnine_unit_5990(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D2),
				.a1(P18E2),
				.a2(P18F2),
				.a3(P19D2),
				.a4(P19E2),
				.a5(P19F2),
				.a6(P1AD2),
				.a7(P1AE2),
				.a8(P1AF2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c128D7)
);

ninexnine_unit ninexnine_unit_5991(
				.clk(clk),
				.rstn(rstn),
				.a0(P18D3),
				.a1(P18E3),
				.a2(P18F3),
				.a3(P19D3),
				.a4(P19E3),
				.a5(P19F3),
				.a6(P1AD3),
				.a7(P1AE3),
				.a8(P1AF3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c138D7)
);

assign C18D7=c108D7+c118D7+c128D7+c138D7;
assign A18D7=(C18D7>=0)?1:0;

ninexnine_unit ninexnine_unit_5992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1900),
				.a1(P1910),
				.a2(P1920),
				.a3(P1A00),
				.a4(P1A10),
				.a5(P1A20),
				.a6(P1B00),
				.a7(P1B10),
				.a8(P1B20),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10907)
);

ninexnine_unit ninexnine_unit_5993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1901),
				.a1(P1911),
				.a2(P1921),
				.a3(P1A01),
				.a4(P1A11),
				.a5(P1A21),
				.a6(P1B01),
				.a7(P1B11),
				.a8(P1B21),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11907)
);

ninexnine_unit ninexnine_unit_5994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1902),
				.a1(P1912),
				.a2(P1922),
				.a3(P1A02),
				.a4(P1A12),
				.a5(P1A22),
				.a6(P1B02),
				.a7(P1B12),
				.a8(P1B22),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12907)
);

ninexnine_unit ninexnine_unit_5995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1903),
				.a1(P1913),
				.a2(P1923),
				.a3(P1A03),
				.a4(P1A13),
				.a5(P1A23),
				.a6(P1B03),
				.a7(P1B13),
				.a8(P1B23),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13907)
);

assign C1907=c10907+c11907+c12907+c13907;
assign A1907=(C1907>=0)?1:0;

ninexnine_unit ninexnine_unit_5996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1910),
				.a1(P1920),
				.a2(P1930),
				.a3(P1A10),
				.a4(P1A20),
				.a5(P1A30),
				.a6(P1B10),
				.a7(P1B20),
				.a8(P1B30),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10917)
);

ninexnine_unit ninexnine_unit_5997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1911),
				.a1(P1921),
				.a2(P1931),
				.a3(P1A11),
				.a4(P1A21),
				.a5(P1A31),
				.a6(P1B11),
				.a7(P1B21),
				.a8(P1B31),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11917)
);

ninexnine_unit ninexnine_unit_5998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1912),
				.a1(P1922),
				.a2(P1932),
				.a3(P1A12),
				.a4(P1A22),
				.a5(P1A32),
				.a6(P1B12),
				.a7(P1B22),
				.a8(P1B32),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12917)
);

ninexnine_unit ninexnine_unit_5999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1913),
				.a1(P1923),
				.a2(P1933),
				.a3(P1A13),
				.a4(P1A23),
				.a5(P1A33),
				.a6(P1B13),
				.a7(P1B23),
				.a8(P1B33),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13917)
);

assign C1917=c10917+c11917+c12917+c13917;
assign A1917=(C1917>=0)?1:0;

ninexnine_unit ninexnine_unit_6000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1920),
				.a1(P1930),
				.a2(P1940),
				.a3(P1A20),
				.a4(P1A30),
				.a5(P1A40),
				.a6(P1B20),
				.a7(P1B30),
				.a8(P1B40),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10927)
);

ninexnine_unit ninexnine_unit_6001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1921),
				.a1(P1931),
				.a2(P1941),
				.a3(P1A21),
				.a4(P1A31),
				.a5(P1A41),
				.a6(P1B21),
				.a7(P1B31),
				.a8(P1B41),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11927)
);

ninexnine_unit ninexnine_unit_6002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1922),
				.a1(P1932),
				.a2(P1942),
				.a3(P1A22),
				.a4(P1A32),
				.a5(P1A42),
				.a6(P1B22),
				.a7(P1B32),
				.a8(P1B42),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12927)
);

ninexnine_unit ninexnine_unit_6003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1923),
				.a1(P1933),
				.a2(P1943),
				.a3(P1A23),
				.a4(P1A33),
				.a5(P1A43),
				.a6(P1B23),
				.a7(P1B33),
				.a8(P1B43),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13927)
);

assign C1927=c10927+c11927+c12927+c13927;
assign A1927=(C1927>=0)?1:0;

ninexnine_unit ninexnine_unit_6004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1930),
				.a1(P1940),
				.a2(P1950),
				.a3(P1A30),
				.a4(P1A40),
				.a5(P1A50),
				.a6(P1B30),
				.a7(P1B40),
				.a8(P1B50),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10937)
);

ninexnine_unit ninexnine_unit_6005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1931),
				.a1(P1941),
				.a2(P1951),
				.a3(P1A31),
				.a4(P1A41),
				.a5(P1A51),
				.a6(P1B31),
				.a7(P1B41),
				.a8(P1B51),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11937)
);

ninexnine_unit ninexnine_unit_6006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1932),
				.a1(P1942),
				.a2(P1952),
				.a3(P1A32),
				.a4(P1A42),
				.a5(P1A52),
				.a6(P1B32),
				.a7(P1B42),
				.a8(P1B52),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12937)
);

ninexnine_unit ninexnine_unit_6007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1933),
				.a1(P1943),
				.a2(P1953),
				.a3(P1A33),
				.a4(P1A43),
				.a5(P1A53),
				.a6(P1B33),
				.a7(P1B43),
				.a8(P1B53),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13937)
);

assign C1937=c10937+c11937+c12937+c13937;
assign A1937=(C1937>=0)?1:0;

ninexnine_unit ninexnine_unit_6008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1940),
				.a1(P1950),
				.a2(P1960),
				.a3(P1A40),
				.a4(P1A50),
				.a5(P1A60),
				.a6(P1B40),
				.a7(P1B50),
				.a8(P1B60),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10947)
);

ninexnine_unit ninexnine_unit_6009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1941),
				.a1(P1951),
				.a2(P1961),
				.a3(P1A41),
				.a4(P1A51),
				.a5(P1A61),
				.a6(P1B41),
				.a7(P1B51),
				.a8(P1B61),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11947)
);

ninexnine_unit ninexnine_unit_6010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1942),
				.a1(P1952),
				.a2(P1962),
				.a3(P1A42),
				.a4(P1A52),
				.a5(P1A62),
				.a6(P1B42),
				.a7(P1B52),
				.a8(P1B62),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12947)
);

ninexnine_unit ninexnine_unit_6011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1943),
				.a1(P1953),
				.a2(P1963),
				.a3(P1A43),
				.a4(P1A53),
				.a5(P1A63),
				.a6(P1B43),
				.a7(P1B53),
				.a8(P1B63),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13947)
);

assign C1947=c10947+c11947+c12947+c13947;
assign A1947=(C1947>=0)?1:0;

ninexnine_unit ninexnine_unit_6012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1950),
				.a1(P1960),
				.a2(P1970),
				.a3(P1A50),
				.a4(P1A60),
				.a5(P1A70),
				.a6(P1B50),
				.a7(P1B60),
				.a8(P1B70),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10957)
);

ninexnine_unit ninexnine_unit_6013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1951),
				.a1(P1961),
				.a2(P1971),
				.a3(P1A51),
				.a4(P1A61),
				.a5(P1A71),
				.a6(P1B51),
				.a7(P1B61),
				.a8(P1B71),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11957)
);

ninexnine_unit ninexnine_unit_6014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1952),
				.a1(P1962),
				.a2(P1972),
				.a3(P1A52),
				.a4(P1A62),
				.a5(P1A72),
				.a6(P1B52),
				.a7(P1B62),
				.a8(P1B72),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12957)
);

ninexnine_unit ninexnine_unit_6015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1953),
				.a1(P1963),
				.a2(P1973),
				.a3(P1A53),
				.a4(P1A63),
				.a5(P1A73),
				.a6(P1B53),
				.a7(P1B63),
				.a8(P1B73),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13957)
);

assign C1957=c10957+c11957+c12957+c13957;
assign A1957=(C1957>=0)?1:0;

ninexnine_unit ninexnine_unit_6016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1960),
				.a1(P1970),
				.a2(P1980),
				.a3(P1A60),
				.a4(P1A70),
				.a5(P1A80),
				.a6(P1B60),
				.a7(P1B70),
				.a8(P1B80),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10967)
);

ninexnine_unit ninexnine_unit_6017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1961),
				.a1(P1971),
				.a2(P1981),
				.a3(P1A61),
				.a4(P1A71),
				.a5(P1A81),
				.a6(P1B61),
				.a7(P1B71),
				.a8(P1B81),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11967)
);

ninexnine_unit ninexnine_unit_6018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1962),
				.a1(P1972),
				.a2(P1982),
				.a3(P1A62),
				.a4(P1A72),
				.a5(P1A82),
				.a6(P1B62),
				.a7(P1B72),
				.a8(P1B82),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12967)
);

ninexnine_unit ninexnine_unit_6019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1963),
				.a1(P1973),
				.a2(P1983),
				.a3(P1A63),
				.a4(P1A73),
				.a5(P1A83),
				.a6(P1B63),
				.a7(P1B73),
				.a8(P1B83),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13967)
);

assign C1967=c10967+c11967+c12967+c13967;
assign A1967=(C1967>=0)?1:0;

ninexnine_unit ninexnine_unit_6020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1970),
				.a1(P1980),
				.a2(P1990),
				.a3(P1A70),
				.a4(P1A80),
				.a5(P1A90),
				.a6(P1B70),
				.a7(P1B80),
				.a8(P1B90),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10977)
);

ninexnine_unit ninexnine_unit_6021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1971),
				.a1(P1981),
				.a2(P1991),
				.a3(P1A71),
				.a4(P1A81),
				.a5(P1A91),
				.a6(P1B71),
				.a7(P1B81),
				.a8(P1B91),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11977)
);

ninexnine_unit ninexnine_unit_6022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1972),
				.a1(P1982),
				.a2(P1992),
				.a3(P1A72),
				.a4(P1A82),
				.a5(P1A92),
				.a6(P1B72),
				.a7(P1B82),
				.a8(P1B92),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12977)
);

ninexnine_unit ninexnine_unit_6023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1973),
				.a1(P1983),
				.a2(P1993),
				.a3(P1A73),
				.a4(P1A83),
				.a5(P1A93),
				.a6(P1B73),
				.a7(P1B83),
				.a8(P1B93),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13977)
);

assign C1977=c10977+c11977+c12977+c13977;
assign A1977=(C1977>=0)?1:0;

ninexnine_unit ninexnine_unit_6024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1980),
				.a1(P1990),
				.a2(P19A0),
				.a3(P1A80),
				.a4(P1A90),
				.a5(P1AA0),
				.a6(P1B80),
				.a7(P1B90),
				.a8(P1BA0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10987)
);

ninexnine_unit ninexnine_unit_6025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1981),
				.a1(P1991),
				.a2(P19A1),
				.a3(P1A81),
				.a4(P1A91),
				.a5(P1AA1),
				.a6(P1B81),
				.a7(P1B91),
				.a8(P1BA1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11987)
);

ninexnine_unit ninexnine_unit_6026(
				.clk(clk),
				.rstn(rstn),
				.a0(P1982),
				.a1(P1992),
				.a2(P19A2),
				.a3(P1A82),
				.a4(P1A92),
				.a5(P1AA2),
				.a6(P1B82),
				.a7(P1B92),
				.a8(P1BA2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12987)
);

ninexnine_unit ninexnine_unit_6027(
				.clk(clk),
				.rstn(rstn),
				.a0(P1983),
				.a1(P1993),
				.a2(P19A3),
				.a3(P1A83),
				.a4(P1A93),
				.a5(P1AA3),
				.a6(P1B83),
				.a7(P1B93),
				.a8(P1BA3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13987)
);

assign C1987=c10987+c11987+c12987+c13987;
assign A1987=(C1987>=0)?1:0;

ninexnine_unit ninexnine_unit_6028(
				.clk(clk),
				.rstn(rstn),
				.a0(P1990),
				.a1(P19A0),
				.a2(P19B0),
				.a3(P1A90),
				.a4(P1AA0),
				.a5(P1AB0),
				.a6(P1B90),
				.a7(P1BA0),
				.a8(P1BB0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10997)
);

ninexnine_unit ninexnine_unit_6029(
				.clk(clk),
				.rstn(rstn),
				.a0(P1991),
				.a1(P19A1),
				.a2(P19B1),
				.a3(P1A91),
				.a4(P1AA1),
				.a5(P1AB1),
				.a6(P1B91),
				.a7(P1BA1),
				.a8(P1BB1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11997)
);

ninexnine_unit ninexnine_unit_6030(
				.clk(clk),
				.rstn(rstn),
				.a0(P1992),
				.a1(P19A2),
				.a2(P19B2),
				.a3(P1A92),
				.a4(P1AA2),
				.a5(P1AB2),
				.a6(P1B92),
				.a7(P1BA2),
				.a8(P1BB2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12997)
);

ninexnine_unit ninexnine_unit_6031(
				.clk(clk),
				.rstn(rstn),
				.a0(P1993),
				.a1(P19A3),
				.a2(P19B3),
				.a3(P1A93),
				.a4(P1AA3),
				.a5(P1AB3),
				.a6(P1B93),
				.a7(P1BA3),
				.a8(P1BB3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13997)
);

assign C1997=c10997+c11997+c12997+c13997;
assign A1997=(C1997>=0)?1:0;

ninexnine_unit ninexnine_unit_6032(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A0),
				.a1(P19B0),
				.a2(P19C0),
				.a3(P1AA0),
				.a4(P1AB0),
				.a5(P1AC0),
				.a6(P1BA0),
				.a7(P1BB0),
				.a8(P1BC0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c109A7)
);

ninexnine_unit ninexnine_unit_6033(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A1),
				.a1(P19B1),
				.a2(P19C1),
				.a3(P1AA1),
				.a4(P1AB1),
				.a5(P1AC1),
				.a6(P1BA1),
				.a7(P1BB1),
				.a8(P1BC1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c119A7)
);

ninexnine_unit ninexnine_unit_6034(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A2),
				.a1(P19B2),
				.a2(P19C2),
				.a3(P1AA2),
				.a4(P1AB2),
				.a5(P1AC2),
				.a6(P1BA2),
				.a7(P1BB2),
				.a8(P1BC2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c129A7)
);

ninexnine_unit ninexnine_unit_6035(
				.clk(clk),
				.rstn(rstn),
				.a0(P19A3),
				.a1(P19B3),
				.a2(P19C3),
				.a3(P1AA3),
				.a4(P1AB3),
				.a5(P1AC3),
				.a6(P1BA3),
				.a7(P1BB3),
				.a8(P1BC3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c139A7)
);

assign C19A7=c109A7+c119A7+c129A7+c139A7;
assign A19A7=(C19A7>=0)?1:0;

ninexnine_unit ninexnine_unit_6036(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B0),
				.a1(P19C0),
				.a2(P19D0),
				.a3(P1AB0),
				.a4(P1AC0),
				.a5(P1AD0),
				.a6(P1BB0),
				.a7(P1BC0),
				.a8(P1BD0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c109B7)
);

ninexnine_unit ninexnine_unit_6037(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B1),
				.a1(P19C1),
				.a2(P19D1),
				.a3(P1AB1),
				.a4(P1AC1),
				.a5(P1AD1),
				.a6(P1BB1),
				.a7(P1BC1),
				.a8(P1BD1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c119B7)
);

ninexnine_unit ninexnine_unit_6038(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B2),
				.a1(P19C2),
				.a2(P19D2),
				.a3(P1AB2),
				.a4(P1AC2),
				.a5(P1AD2),
				.a6(P1BB2),
				.a7(P1BC2),
				.a8(P1BD2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c129B7)
);

ninexnine_unit ninexnine_unit_6039(
				.clk(clk),
				.rstn(rstn),
				.a0(P19B3),
				.a1(P19C3),
				.a2(P19D3),
				.a3(P1AB3),
				.a4(P1AC3),
				.a5(P1AD3),
				.a6(P1BB3),
				.a7(P1BC3),
				.a8(P1BD3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c139B7)
);

assign C19B7=c109B7+c119B7+c129B7+c139B7;
assign A19B7=(C19B7>=0)?1:0;

ninexnine_unit ninexnine_unit_6040(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C0),
				.a1(P19D0),
				.a2(P19E0),
				.a3(P1AC0),
				.a4(P1AD0),
				.a5(P1AE0),
				.a6(P1BC0),
				.a7(P1BD0),
				.a8(P1BE0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c109C7)
);

ninexnine_unit ninexnine_unit_6041(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C1),
				.a1(P19D1),
				.a2(P19E1),
				.a3(P1AC1),
				.a4(P1AD1),
				.a5(P1AE1),
				.a6(P1BC1),
				.a7(P1BD1),
				.a8(P1BE1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c119C7)
);

ninexnine_unit ninexnine_unit_6042(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C2),
				.a1(P19D2),
				.a2(P19E2),
				.a3(P1AC2),
				.a4(P1AD2),
				.a5(P1AE2),
				.a6(P1BC2),
				.a7(P1BD2),
				.a8(P1BE2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c129C7)
);

ninexnine_unit ninexnine_unit_6043(
				.clk(clk),
				.rstn(rstn),
				.a0(P19C3),
				.a1(P19D3),
				.a2(P19E3),
				.a3(P1AC3),
				.a4(P1AD3),
				.a5(P1AE3),
				.a6(P1BC3),
				.a7(P1BD3),
				.a8(P1BE3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c139C7)
);

assign C19C7=c109C7+c119C7+c129C7+c139C7;
assign A19C7=(C19C7>=0)?1:0;

ninexnine_unit ninexnine_unit_6044(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D0),
				.a1(P19E0),
				.a2(P19F0),
				.a3(P1AD0),
				.a4(P1AE0),
				.a5(P1AF0),
				.a6(P1BD0),
				.a7(P1BE0),
				.a8(P1BF0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c109D7)
);

ninexnine_unit ninexnine_unit_6045(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D1),
				.a1(P19E1),
				.a2(P19F1),
				.a3(P1AD1),
				.a4(P1AE1),
				.a5(P1AF1),
				.a6(P1BD1),
				.a7(P1BE1),
				.a8(P1BF1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c119D7)
);

ninexnine_unit ninexnine_unit_6046(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D2),
				.a1(P19E2),
				.a2(P19F2),
				.a3(P1AD2),
				.a4(P1AE2),
				.a5(P1AF2),
				.a6(P1BD2),
				.a7(P1BE2),
				.a8(P1BF2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c129D7)
);

ninexnine_unit ninexnine_unit_6047(
				.clk(clk),
				.rstn(rstn),
				.a0(P19D3),
				.a1(P19E3),
				.a2(P19F3),
				.a3(P1AD3),
				.a4(P1AE3),
				.a5(P1AF3),
				.a6(P1BD3),
				.a7(P1BE3),
				.a8(P1BF3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c139D7)
);

assign C19D7=c109D7+c119D7+c129D7+c139D7;
assign A19D7=(C19D7>=0)?1:0;

ninexnine_unit ninexnine_unit_6048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A00),
				.a1(P1A10),
				.a2(P1A20),
				.a3(P1B00),
				.a4(P1B10),
				.a5(P1B20),
				.a6(P1C00),
				.a7(P1C10),
				.a8(P1C20),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A07)
);

ninexnine_unit ninexnine_unit_6049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A01),
				.a1(P1A11),
				.a2(P1A21),
				.a3(P1B01),
				.a4(P1B11),
				.a5(P1B21),
				.a6(P1C01),
				.a7(P1C11),
				.a8(P1C21),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A07)
);

ninexnine_unit ninexnine_unit_6050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A02),
				.a1(P1A12),
				.a2(P1A22),
				.a3(P1B02),
				.a4(P1B12),
				.a5(P1B22),
				.a6(P1C02),
				.a7(P1C12),
				.a8(P1C22),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A07)
);

ninexnine_unit ninexnine_unit_6051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A03),
				.a1(P1A13),
				.a2(P1A23),
				.a3(P1B03),
				.a4(P1B13),
				.a5(P1B23),
				.a6(P1C03),
				.a7(P1C13),
				.a8(P1C23),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A07)
);

assign C1A07=c10A07+c11A07+c12A07+c13A07;
assign A1A07=(C1A07>=0)?1:0;

ninexnine_unit ninexnine_unit_6052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A10),
				.a1(P1A20),
				.a2(P1A30),
				.a3(P1B10),
				.a4(P1B20),
				.a5(P1B30),
				.a6(P1C10),
				.a7(P1C20),
				.a8(P1C30),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A17)
);

ninexnine_unit ninexnine_unit_6053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A11),
				.a1(P1A21),
				.a2(P1A31),
				.a3(P1B11),
				.a4(P1B21),
				.a5(P1B31),
				.a6(P1C11),
				.a7(P1C21),
				.a8(P1C31),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A17)
);

ninexnine_unit ninexnine_unit_6054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A12),
				.a1(P1A22),
				.a2(P1A32),
				.a3(P1B12),
				.a4(P1B22),
				.a5(P1B32),
				.a6(P1C12),
				.a7(P1C22),
				.a8(P1C32),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A17)
);

ninexnine_unit ninexnine_unit_6055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A13),
				.a1(P1A23),
				.a2(P1A33),
				.a3(P1B13),
				.a4(P1B23),
				.a5(P1B33),
				.a6(P1C13),
				.a7(P1C23),
				.a8(P1C33),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A17)
);

assign C1A17=c10A17+c11A17+c12A17+c13A17;
assign A1A17=(C1A17>=0)?1:0;

ninexnine_unit ninexnine_unit_6056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A20),
				.a1(P1A30),
				.a2(P1A40),
				.a3(P1B20),
				.a4(P1B30),
				.a5(P1B40),
				.a6(P1C20),
				.a7(P1C30),
				.a8(P1C40),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A27)
);

ninexnine_unit ninexnine_unit_6057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A21),
				.a1(P1A31),
				.a2(P1A41),
				.a3(P1B21),
				.a4(P1B31),
				.a5(P1B41),
				.a6(P1C21),
				.a7(P1C31),
				.a8(P1C41),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A27)
);

ninexnine_unit ninexnine_unit_6058(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A22),
				.a1(P1A32),
				.a2(P1A42),
				.a3(P1B22),
				.a4(P1B32),
				.a5(P1B42),
				.a6(P1C22),
				.a7(P1C32),
				.a8(P1C42),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A27)
);

ninexnine_unit ninexnine_unit_6059(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A23),
				.a1(P1A33),
				.a2(P1A43),
				.a3(P1B23),
				.a4(P1B33),
				.a5(P1B43),
				.a6(P1C23),
				.a7(P1C33),
				.a8(P1C43),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A27)
);

assign C1A27=c10A27+c11A27+c12A27+c13A27;
assign A1A27=(C1A27>=0)?1:0;

ninexnine_unit ninexnine_unit_6060(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A30),
				.a1(P1A40),
				.a2(P1A50),
				.a3(P1B30),
				.a4(P1B40),
				.a5(P1B50),
				.a6(P1C30),
				.a7(P1C40),
				.a8(P1C50),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A37)
);

ninexnine_unit ninexnine_unit_6061(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A31),
				.a1(P1A41),
				.a2(P1A51),
				.a3(P1B31),
				.a4(P1B41),
				.a5(P1B51),
				.a6(P1C31),
				.a7(P1C41),
				.a8(P1C51),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A37)
);

ninexnine_unit ninexnine_unit_6062(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A32),
				.a1(P1A42),
				.a2(P1A52),
				.a3(P1B32),
				.a4(P1B42),
				.a5(P1B52),
				.a6(P1C32),
				.a7(P1C42),
				.a8(P1C52),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A37)
);

ninexnine_unit ninexnine_unit_6063(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A33),
				.a1(P1A43),
				.a2(P1A53),
				.a3(P1B33),
				.a4(P1B43),
				.a5(P1B53),
				.a6(P1C33),
				.a7(P1C43),
				.a8(P1C53),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A37)
);

assign C1A37=c10A37+c11A37+c12A37+c13A37;
assign A1A37=(C1A37>=0)?1:0;

ninexnine_unit ninexnine_unit_6064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A40),
				.a1(P1A50),
				.a2(P1A60),
				.a3(P1B40),
				.a4(P1B50),
				.a5(P1B60),
				.a6(P1C40),
				.a7(P1C50),
				.a8(P1C60),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A47)
);

ninexnine_unit ninexnine_unit_6065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A41),
				.a1(P1A51),
				.a2(P1A61),
				.a3(P1B41),
				.a4(P1B51),
				.a5(P1B61),
				.a6(P1C41),
				.a7(P1C51),
				.a8(P1C61),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A47)
);

ninexnine_unit ninexnine_unit_6066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A42),
				.a1(P1A52),
				.a2(P1A62),
				.a3(P1B42),
				.a4(P1B52),
				.a5(P1B62),
				.a6(P1C42),
				.a7(P1C52),
				.a8(P1C62),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A47)
);

ninexnine_unit ninexnine_unit_6067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A43),
				.a1(P1A53),
				.a2(P1A63),
				.a3(P1B43),
				.a4(P1B53),
				.a5(P1B63),
				.a6(P1C43),
				.a7(P1C53),
				.a8(P1C63),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A47)
);

assign C1A47=c10A47+c11A47+c12A47+c13A47;
assign A1A47=(C1A47>=0)?1:0;

ninexnine_unit ninexnine_unit_6068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A50),
				.a1(P1A60),
				.a2(P1A70),
				.a3(P1B50),
				.a4(P1B60),
				.a5(P1B70),
				.a6(P1C50),
				.a7(P1C60),
				.a8(P1C70),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A57)
);

ninexnine_unit ninexnine_unit_6069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A51),
				.a1(P1A61),
				.a2(P1A71),
				.a3(P1B51),
				.a4(P1B61),
				.a5(P1B71),
				.a6(P1C51),
				.a7(P1C61),
				.a8(P1C71),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A57)
);

ninexnine_unit ninexnine_unit_6070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A52),
				.a1(P1A62),
				.a2(P1A72),
				.a3(P1B52),
				.a4(P1B62),
				.a5(P1B72),
				.a6(P1C52),
				.a7(P1C62),
				.a8(P1C72),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A57)
);

ninexnine_unit ninexnine_unit_6071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A53),
				.a1(P1A63),
				.a2(P1A73),
				.a3(P1B53),
				.a4(P1B63),
				.a5(P1B73),
				.a6(P1C53),
				.a7(P1C63),
				.a8(P1C73),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A57)
);

assign C1A57=c10A57+c11A57+c12A57+c13A57;
assign A1A57=(C1A57>=0)?1:0;

ninexnine_unit ninexnine_unit_6072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A60),
				.a1(P1A70),
				.a2(P1A80),
				.a3(P1B60),
				.a4(P1B70),
				.a5(P1B80),
				.a6(P1C60),
				.a7(P1C70),
				.a8(P1C80),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A67)
);

ninexnine_unit ninexnine_unit_6073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A61),
				.a1(P1A71),
				.a2(P1A81),
				.a3(P1B61),
				.a4(P1B71),
				.a5(P1B81),
				.a6(P1C61),
				.a7(P1C71),
				.a8(P1C81),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A67)
);

ninexnine_unit ninexnine_unit_6074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A62),
				.a1(P1A72),
				.a2(P1A82),
				.a3(P1B62),
				.a4(P1B72),
				.a5(P1B82),
				.a6(P1C62),
				.a7(P1C72),
				.a8(P1C82),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A67)
);

ninexnine_unit ninexnine_unit_6075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A63),
				.a1(P1A73),
				.a2(P1A83),
				.a3(P1B63),
				.a4(P1B73),
				.a5(P1B83),
				.a6(P1C63),
				.a7(P1C73),
				.a8(P1C83),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A67)
);

assign C1A67=c10A67+c11A67+c12A67+c13A67;
assign A1A67=(C1A67>=0)?1:0;

ninexnine_unit ninexnine_unit_6076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A70),
				.a1(P1A80),
				.a2(P1A90),
				.a3(P1B70),
				.a4(P1B80),
				.a5(P1B90),
				.a6(P1C70),
				.a7(P1C80),
				.a8(P1C90),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A77)
);

ninexnine_unit ninexnine_unit_6077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A71),
				.a1(P1A81),
				.a2(P1A91),
				.a3(P1B71),
				.a4(P1B81),
				.a5(P1B91),
				.a6(P1C71),
				.a7(P1C81),
				.a8(P1C91),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A77)
);

ninexnine_unit ninexnine_unit_6078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A72),
				.a1(P1A82),
				.a2(P1A92),
				.a3(P1B72),
				.a4(P1B82),
				.a5(P1B92),
				.a6(P1C72),
				.a7(P1C82),
				.a8(P1C92),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A77)
);

ninexnine_unit ninexnine_unit_6079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A73),
				.a1(P1A83),
				.a2(P1A93),
				.a3(P1B73),
				.a4(P1B83),
				.a5(P1B93),
				.a6(P1C73),
				.a7(P1C83),
				.a8(P1C93),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A77)
);

assign C1A77=c10A77+c11A77+c12A77+c13A77;
assign A1A77=(C1A77>=0)?1:0;

ninexnine_unit ninexnine_unit_6080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A80),
				.a1(P1A90),
				.a2(P1AA0),
				.a3(P1B80),
				.a4(P1B90),
				.a5(P1BA0),
				.a6(P1C80),
				.a7(P1C90),
				.a8(P1CA0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A87)
);

ninexnine_unit ninexnine_unit_6081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A81),
				.a1(P1A91),
				.a2(P1AA1),
				.a3(P1B81),
				.a4(P1B91),
				.a5(P1BA1),
				.a6(P1C81),
				.a7(P1C91),
				.a8(P1CA1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A87)
);

ninexnine_unit ninexnine_unit_6082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A82),
				.a1(P1A92),
				.a2(P1AA2),
				.a3(P1B82),
				.a4(P1B92),
				.a5(P1BA2),
				.a6(P1C82),
				.a7(P1C92),
				.a8(P1CA2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A87)
);

ninexnine_unit ninexnine_unit_6083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A83),
				.a1(P1A93),
				.a2(P1AA3),
				.a3(P1B83),
				.a4(P1B93),
				.a5(P1BA3),
				.a6(P1C83),
				.a7(P1C93),
				.a8(P1CA3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A87)
);

assign C1A87=c10A87+c11A87+c12A87+c13A87;
assign A1A87=(C1A87>=0)?1:0;

ninexnine_unit ninexnine_unit_6084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A90),
				.a1(P1AA0),
				.a2(P1AB0),
				.a3(P1B90),
				.a4(P1BA0),
				.a5(P1BB0),
				.a6(P1C90),
				.a7(P1CA0),
				.a8(P1CB0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10A97)
);

ninexnine_unit ninexnine_unit_6085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A91),
				.a1(P1AA1),
				.a2(P1AB1),
				.a3(P1B91),
				.a4(P1BA1),
				.a5(P1BB1),
				.a6(P1C91),
				.a7(P1CA1),
				.a8(P1CB1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11A97)
);

ninexnine_unit ninexnine_unit_6086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A92),
				.a1(P1AA2),
				.a2(P1AB2),
				.a3(P1B92),
				.a4(P1BA2),
				.a5(P1BB2),
				.a6(P1C92),
				.a7(P1CA2),
				.a8(P1CB2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12A97)
);

ninexnine_unit ninexnine_unit_6087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1A93),
				.a1(P1AA3),
				.a2(P1AB3),
				.a3(P1B93),
				.a4(P1BA3),
				.a5(P1BB3),
				.a6(P1C93),
				.a7(P1CA3),
				.a8(P1CB3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13A97)
);

assign C1A97=c10A97+c11A97+c12A97+c13A97;
assign A1A97=(C1A97>=0)?1:0;

ninexnine_unit ninexnine_unit_6088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA0),
				.a1(P1AB0),
				.a2(P1AC0),
				.a3(P1BA0),
				.a4(P1BB0),
				.a5(P1BC0),
				.a6(P1CA0),
				.a7(P1CB0),
				.a8(P1CC0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10AA7)
);

ninexnine_unit ninexnine_unit_6089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA1),
				.a1(P1AB1),
				.a2(P1AC1),
				.a3(P1BA1),
				.a4(P1BB1),
				.a5(P1BC1),
				.a6(P1CA1),
				.a7(P1CB1),
				.a8(P1CC1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11AA7)
);

ninexnine_unit ninexnine_unit_6090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA2),
				.a1(P1AB2),
				.a2(P1AC2),
				.a3(P1BA2),
				.a4(P1BB2),
				.a5(P1BC2),
				.a6(P1CA2),
				.a7(P1CB2),
				.a8(P1CC2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12AA7)
);

ninexnine_unit ninexnine_unit_6091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AA3),
				.a1(P1AB3),
				.a2(P1AC3),
				.a3(P1BA3),
				.a4(P1BB3),
				.a5(P1BC3),
				.a6(P1CA3),
				.a7(P1CB3),
				.a8(P1CC3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13AA7)
);

assign C1AA7=c10AA7+c11AA7+c12AA7+c13AA7;
assign A1AA7=(C1AA7>=0)?1:0;

ninexnine_unit ninexnine_unit_6092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB0),
				.a1(P1AC0),
				.a2(P1AD0),
				.a3(P1BB0),
				.a4(P1BC0),
				.a5(P1BD0),
				.a6(P1CB0),
				.a7(P1CC0),
				.a8(P1CD0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10AB7)
);

ninexnine_unit ninexnine_unit_6093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB1),
				.a1(P1AC1),
				.a2(P1AD1),
				.a3(P1BB1),
				.a4(P1BC1),
				.a5(P1BD1),
				.a6(P1CB1),
				.a7(P1CC1),
				.a8(P1CD1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11AB7)
);

ninexnine_unit ninexnine_unit_6094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB2),
				.a1(P1AC2),
				.a2(P1AD2),
				.a3(P1BB2),
				.a4(P1BC2),
				.a5(P1BD2),
				.a6(P1CB2),
				.a7(P1CC2),
				.a8(P1CD2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12AB7)
);

ninexnine_unit ninexnine_unit_6095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AB3),
				.a1(P1AC3),
				.a2(P1AD3),
				.a3(P1BB3),
				.a4(P1BC3),
				.a5(P1BD3),
				.a6(P1CB3),
				.a7(P1CC3),
				.a8(P1CD3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13AB7)
);

assign C1AB7=c10AB7+c11AB7+c12AB7+c13AB7;
assign A1AB7=(C1AB7>=0)?1:0;

ninexnine_unit ninexnine_unit_6096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC0),
				.a1(P1AD0),
				.a2(P1AE0),
				.a3(P1BC0),
				.a4(P1BD0),
				.a5(P1BE0),
				.a6(P1CC0),
				.a7(P1CD0),
				.a8(P1CE0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10AC7)
);

ninexnine_unit ninexnine_unit_6097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC1),
				.a1(P1AD1),
				.a2(P1AE1),
				.a3(P1BC1),
				.a4(P1BD1),
				.a5(P1BE1),
				.a6(P1CC1),
				.a7(P1CD1),
				.a8(P1CE1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11AC7)
);

ninexnine_unit ninexnine_unit_6098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC2),
				.a1(P1AD2),
				.a2(P1AE2),
				.a3(P1BC2),
				.a4(P1BD2),
				.a5(P1BE2),
				.a6(P1CC2),
				.a7(P1CD2),
				.a8(P1CE2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12AC7)
);

ninexnine_unit ninexnine_unit_6099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AC3),
				.a1(P1AD3),
				.a2(P1AE3),
				.a3(P1BC3),
				.a4(P1BD3),
				.a5(P1BE3),
				.a6(P1CC3),
				.a7(P1CD3),
				.a8(P1CE3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13AC7)
);

assign C1AC7=c10AC7+c11AC7+c12AC7+c13AC7;
assign A1AC7=(C1AC7>=0)?1:0;

ninexnine_unit ninexnine_unit_6100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD0),
				.a1(P1AE0),
				.a2(P1AF0),
				.a3(P1BD0),
				.a4(P1BE0),
				.a5(P1BF0),
				.a6(P1CD0),
				.a7(P1CE0),
				.a8(P1CF0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10AD7)
);

ninexnine_unit ninexnine_unit_6101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD1),
				.a1(P1AE1),
				.a2(P1AF1),
				.a3(P1BD1),
				.a4(P1BE1),
				.a5(P1BF1),
				.a6(P1CD1),
				.a7(P1CE1),
				.a8(P1CF1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11AD7)
);

ninexnine_unit ninexnine_unit_6102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD2),
				.a1(P1AE2),
				.a2(P1AF2),
				.a3(P1BD2),
				.a4(P1BE2),
				.a5(P1BF2),
				.a6(P1CD2),
				.a7(P1CE2),
				.a8(P1CF2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12AD7)
);

ninexnine_unit ninexnine_unit_6103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1AD3),
				.a1(P1AE3),
				.a2(P1AF3),
				.a3(P1BD3),
				.a4(P1BE3),
				.a5(P1BF3),
				.a6(P1CD3),
				.a7(P1CE3),
				.a8(P1CF3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13AD7)
);

assign C1AD7=c10AD7+c11AD7+c12AD7+c13AD7;
assign A1AD7=(C1AD7>=0)?1:0;

ninexnine_unit ninexnine_unit_6104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B00),
				.a1(P1B10),
				.a2(P1B20),
				.a3(P1C00),
				.a4(P1C10),
				.a5(P1C20),
				.a6(P1D00),
				.a7(P1D10),
				.a8(P1D20),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B07)
);

ninexnine_unit ninexnine_unit_6105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B01),
				.a1(P1B11),
				.a2(P1B21),
				.a3(P1C01),
				.a4(P1C11),
				.a5(P1C21),
				.a6(P1D01),
				.a7(P1D11),
				.a8(P1D21),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B07)
);

ninexnine_unit ninexnine_unit_6106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B02),
				.a1(P1B12),
				.a2(P1B22),
				.a3(P1C02),
				.a4(P1C12),
				.a5(P1C22),
				.a6(P1D02),
				.a7(P1D12),
				.a8(P1D22),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B07)
);

ninexnine_unit ninexnine_unit_6107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B03),
				.a1(P1B13),
				.a2(P1B23),
				.a3(P1C03),
				.a4(P1C13),
				.a5(P1C23),
				.a6(P1D03),
				.a7(P1D13),
				.a8(P1D23),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B07)
);

assign C1B07=c10B07+c11B07+c12B07+c13B07;
assign A1B07=(C1B07>=0)?1:0;

ninexnine_unit ninexnine_unit_6108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B10),
				.a1(P1B20),
				.a2(P1B30),
				.a3(P1C10),
				.a4(P1C20),
				.a5(P1C30),
				.a6(P1D10),
				.a7(P1D20),
				.a8(P1D30),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B17)
);

ninexnine_unit ninexnine_unit_6109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B11),
				.a1(P1B21),
				.a2(P1B31),
				.a3(P1C11),
				.a4(P1C21),
				.a5(P1C31),
				.a6(P1D11),
				.a7(P1D21),
				.a8(P1D31),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B17)
);

ninexnine_unit ninexnine_unit_6110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B12),
				.a1(P1B22),
				.a2(P1B32),
				.a3(P1C12),
				.a4(P1C22),
				.a5(P1C32),
				.a6(P1D12),
				.a7(P1D22),
				.a8(P1D32),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B17)
);

ninexnine_unit ninexnine_unit_6111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B13),
				.a1(P1B23),
				.a2(P1B33),
				.a3(P1C13),
				.a4(P1C23),
				.a5(P1C33),
				.a6(P1D13),
				.a7(P1D23),
				.a8(P1D33),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B17)
);

assign C1B17=c10B17+c11B17+c12B17+c13B17;
assign A1B17=(C1B17>=0)?1:0;

ninexnine_unit ninexnine_unit_6112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B20),
				.a1(P1B30),
				.a2(P1B40),
				.a3(P1C20),
				.a4(P1C30),
				.a5(P1C40),
				.a6(P1D20),
				.a7(P1D30),
				.a8(P1D40),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B27)
);

ninexnine_unit ninexnine_unit_6113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B21),
				.a1(P1B31),
				.a2(P1B41),
				.a3(P1C21),
				.a4(P1C31),
				.a5(P1C41),
				.a6(P1D21),
				.a7(P1D31),
				.a8(P1D41),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B27)
);

ninexnine_unit ninexnine_unit_6114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B22),
				.a1(P1B32),
				.a2(P1B42),
				.a3(P1C22),
				.a4(P1C32),
				.a5(P1C42),
				.a6(P1D22),
				.a7(P1D32),
				.a8(P1D42),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B27)
);

ninexnine_unit ninexnine_unit_6115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B23),
				.a1(P1B33),
				.a2(P1B43),
				.a3(P1C23),
				.a4(P1C33),
				.a5(P1C43),
				.a6(P1D23),
				.a7(P1D33),
				.a8(P1D43),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B27)
);

assign C1B27=c10B27+c11B27+c12B27+c13B27;
assign A1B27=(C1B27>=0)?1:0;

ninexnine_unit ninexnine_unit_6116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B30),
				.a1(P1B40),
				.a2(P1B50),
				.a3(P1C30),
				.a4(P1C40),
				.a5(P1C50),
				.a6(P1D30),
				.a7(P1D40),
				.a8(P1D50),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B37)
);

ninexnine_unit ninexnine_unit_6117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B31),
				.a1(P1B41),
				.a2(P1B51),
				.a3(P1C31),
				.a4(P1C41),
				.a5(P1C51),
				.a6(P1D31),
				.a7(P1D41),
				.a8(P1D51),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B37)
);

ninexnine_unit ninexnine_unit_6118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B32),
				.a1(P1B42),
				.a2(P1B52),
				.a3(P1C32),
				.a4(P1C42),
				.a5(P1C52),
				.a6(P1D32),
				.a7(P1D42),
				.a8(P1D52),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B37)
);

ninexnine_unit ninexnine_unit_6119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B33),
				.a1(P1B43),
				.a2(P1B53),
				.a3(P1C33),
				.a4(P1C43),
				.a5(P1C53),
				.a6(P1D33),
				.a7(P1D43),
				.a8(P1D53),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B37)
);

assign C1B37=c10B37+c11B37+c12B37+c13B37;
assign A1B37=(C1B37>=0)?1:0;

ninexnine_unit ninexnine_unit_6120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B40),
				.a1(P1B50),
				.a2(P1B60),
				.a3(P1C40),
				.a4(P1C50),
				.a5(P1C60),
				.a6(P1D40),
				.a7(P1D50),
				.a8(P1D60),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B47)
);

ninexnine_unit ninexnine_unit_6121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B41),
				.a1(P1B51),
				.a2(P1B61),
				.a3(P1C41),
				.a4(P1C51),
				.a5(P1C61),
				.a6(P1D41),
				.a7(P1D51),
				.a8(P1D61),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B47)
);

ninexnine_unit ninexnine_unit_6122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B42),
				.a1(P1B52),
				.a2(P1B62),
				.a3(P1C42),
				.a4(P1C52),
				.a5(P1C62),
				.a6(P1D42),
				.a7(P1D52),
				.a8(P1D62),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B47)
);

ninexnine_unit ninexnine_unit_6123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B43),
				.a1(P1B53),
				.a2(P1B63),
				.a3(P1C43),
				.a4(P1C53),
				.a5(P1C63),
				.a6(P1D43),
				.a7(P1D53),
				.a8(P1D63),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B47)
);

assign C1B47=c10B47+c11B47+c12B47+c13B47;
assign A1B47=(C1B47>=0)?1:0;

ninexnine_unit ninexnine_unit_6124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B50),
				.a1(P1B60),
				.a2(P1B70),
				.a3(P1C50),
				.a4(P1C60),
				.a5(P1C70),
				.a6(P1D50),
				.a7(P1D60),
				.a8(P1D70),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B57)
);

ninexnine_unit ninexnine_unit_6125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B51),
				.a1(P1B61),
				.a2(P1B71),
				.a3(P1C51),
				.a4(P1C61),
				.a5(P1C71),
				.a6(P1D51),
				.a7(P1D61),
				.a8(P1D71),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B57)
);

ninexnine_unit ninexnine_unit_6126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B52),
				.a1(P1B62),
				.a2(P1B72),
				.a3(P1C52),
				.a4(P1C62),
				.a5(P1C72),
				.a6(P1D52),
				.a7(P1D62),
				.a8(P1D72),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B57)
);

ninexnine_unit ninexnine_unit_6127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B53),
				.a1(P1B63),
				.a2(P1B73),
				.a3(P1C53),
				.a4(P1C63),
				.a5(P1C73),
				.a6(P1D53),
				.a7(P1D63),
				.a8(P1D73),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B57)
);

assign C1B57=c10B57+c11B57+c12B57+c13B57;
assign A1B57=(C1B57>=0)?1:0;

ninexnine_unit ninexnine_unit_6128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B60),
				.a1(P1B70),
				.a2(P1B80),
				.a3(P1C60),
				.a4(P1C70),
				.a5(P1C80),
				.a6(P1D60),
				.a7(P1D70),
				.a8(P1D80),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B67)
);

ninexnine_unit ninexnine_unit_6129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B61),
				.a1(P1B71),
				.a2(P1B81),
				.a3(P1C61),
				.a4(P1C71),
				.a5(P1C81),
				.a6(P1D61),
				.a7(P1D71),
				.a8(P1D81),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B67)
);

ninexnine_unit ninexnine_unit_6130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B62),
				.a1(P1B72),
				.a2(P1B82),
				.a3(P1C62),
				.a4(P1C72),
				.a5(P1C82),
				.a6(P1D62),
				.a7(P1D72),
				.a8(P1D82),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B67)
);

ninexnine_unit ninexnine_unit_6131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B63),
				.a1(P1B73),
				.a2(P1B83),
				.a3(P1C63),
				.a4(P1C73),
				.a5(P1C83),
				.a6(P1D63),
				.a7(P1D73),
				.a8(P1D83),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B67)
);

assign C1B67=c10B67+c11B67+c12B67+c13B67;
assign A1B67=(C1B67>=0)?1:0;

ninexnine_unit ninexnine_unit_6132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B70),
				.a1(P1B80),
				.a2(P1B90),
				.a3(P1C70),
				.a4(P1C80),
				.a5(P1C90),
				.a6(P1D70),
				.a7(P1D80),
				.a8(P1D90),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B77)
);

ninexnine_unit ninexnine_unit_6133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B71),
				.a1(P1B81),
				.a2(P1B91),
				.a3(P1C71),
				.a4(P1C81),
				.a5(P1C91),
				.a6(P1D71),
				.a7(P1D81),
				.a8(P1D91),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B77)
);

ninexnine_unit ninexnine_unit_6134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B72),
				.a1(P1B82),
				.a2(P1B92),
				.a3(P1C72),
				.a4(P1C82),
				.a5(P1C92),
				.a6(P1D72),
				.a7(P1D82),
				.a8(P1D92),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B77)
);

ninexnine_unit ninexnine_unit_6135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B73),
				.a1(P1B83),
				.a2(P1B93),
				.a3(P1C73),
				.a4(P1C83),
				.a5(P1C93),
				.a6(P1D73),
				.a7(P1D83),
				.a8(P1D93),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B77)
);

assign C1B77=c10B77+c11B77+c12B77+c13B77;
assign A1B77=(C1B77>=0)?1:0;

ninexnine_unit ninexnine_unit_6136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B80),
				.a1(P1B90),
				.a2(P1BA0),
				.a3(P1C80),
				.a4(P1C90),
				.a5(P1CA0),
				.a6(P1D80),
				.a7(P1D90),
				.a8(P1DA0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B87)
);

ninexnine_unit ninexnine_unit_6137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B81),
				.a1(P1B91),
				.a2(P1BA1),
				.a3(P1C81),
				.a4(P1C91),
				.a5(P1CA1),
				.a6(P1D81),
				.a7(P1D91),
				.a8(P1DA1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B87)
);

ninexnine_unit ninexnine_unit_6138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B82),
				.a1(P1B92),
				.a2(P1BA2),
				.a3(P1C82),
				.a4(P1C92),
				.a5(P1CA2),
				.a6(P1D82),
				.a7(P1D92),
				.a8(P1DA2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B87)
);

ninexnine_unit ninexnine_unit_6139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B83),
				.a1(P1B93),
				.a2(P1BA3),
				.a3(P1C83),
				.a4(P1C93),
				.a5(P1CA3),
				.a6(P1D83),
				.a7(P1D93),
				.a8(P1DA3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B87)
);

assign C1B87=c10B87+c11B87+c12B87+c13B87;
assign A1B87=(C1B87>=0)?1:0;

ninexnine_unit ninexnine_unit_6140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B90),
				.a1(P1BA0),
				.a2(P1BB0),
				.a3(P1C90),
				.a4(P1CA0),
				.a5(P1CB0),
				.a6(P1D90),
				.a7(P1DA0),
				.a8(P1DB0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10B97)
);

ninexnine_unit ninexnine_unit_6141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B91),
				.a1(P1BA1),
				.a2(P1BB1),
				.a3(P1C91),
				.a4(P1CA1),
				.a5(P1CB1),
				.a6(P1D91),
				.a7(P1DA1),
				.a8(P1DB1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11B97)
);

ninexnine_unit ninexnine_unit_6142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B92),
				.a1(P1BA2),
				.a2(P1BB2),
				.a3(P1C92),
				.a4(P1CA2),
				.a5(P1CB2),
				.a6(P1D92),
				.a7(P1DA2),
				.a8(P1DB2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12B97)
);

ninexnine_unit ninexnine_unit_6143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1B93),
				.a1(P1BA3),
				.a2(P1BB3),
				.a3(P1C93),
				.a4(P1CA3),
				.a5(P1CB3),
				.a6(P1D93),
				.a7(P1DA3),
				.a8(P1DB3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13B97)
);

assign C1B97=c10B97+c11B97+c12B97+c13B97;
assign A1B97=(C1B97>=0)?1:0;

ninexnine_unit ninexnine_unit_6144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA0),
				.a1(P1BB0),
				.a2(P1BC0),
				.a3(P1CA0),
				.a4(P1CB0),
				.a5(P1CC0),
				.a6(P1DA0),
				.a7(P1DB0),
				.a8(P1DC0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10BA7)
);

ninexnine_unit ninexnine_unit_6145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA1),
				.a1(P1BB1),
				.a2(P1BC1),
				.a3(P1CA1),
				.a4(P1CB1),
				.a5(P1CC1),
				.a6(P1DA1),
				.a7(P1DB1),
				.a8(P1DC1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11BA7)
);

ninexnine_unit ninexnine_unit_6146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA2),
				.a1(P1BB2),
				.a2(P1BC2),
				.a3(P1CA2),
				.a4(P1CB2),
				.a5(P1CC2),
				.a6(P1DA2),
				.a7(P1DB2),
				.a8(P1DC2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12BA7)
);

ninexnine_unit ninexnine_unit_6147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BA3),
				.a1(P1BB3),
				.a2(P1BC3),
				.a3(P1CA3),
				.a4(P1CB3),
				.a5(P1CC3),
				.a6(P1DA3),
				.a7(P1DB3),
				.a8(P1DC3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13BA7)
);

assign C1BA7=c10BA7+c11BA7+c12BA7+c13BA7;
assign A1BA7=(C1BA7>=0)?1:0;

ninexnine_unit ninexnine_unit_6148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB0),
				.a1(P1BC0),
				.a2(P1BD0),
				.a3(P1CB0),
				.a4(P1CC0),
				.a5(P1CD0),
				.a6(P1DB0),
				.a7(P1DC0),
				.a8(P1DD0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10BB7)
);

ninexnine_unit ninexnine_unit_6149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB1),
				.a1(P1BC1),
				.a2(P1BD1),
				.a3(P1CB1),
				.a4(P1CC1),
				.a5(P1CD1),
				.a6(P1DB1),
				.a7(P1DC1),
				.a8(P1DD1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11BB7)
);

ninexnine_unit ninexnine_unit_6150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB2),
				.a1(P1BC2),
				.a2(P1BD2),
				.a3(P1CB2),
				.a4(P1CC2),
				.a5(P1CD2),
				.a6(P1DB2),
				.a7(P1DC2),
				.a8(P1DD2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12BB7)
);

ninexnine_unit ninexnine_unit_6151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BB3),
				.a1(P1BC3),
				.a2(P1BD3),
				.a3(P1CB3),
				.a4(P1CC3),
				.a5(P1CD3),
				.a6(P1DB3),
				.a7(P1DC3),
				.a8(P1DD3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13BB7)
);

assign C1BB7=c10BB7+c11BB7+c12BB7+c13BB7;
assign A1BB7=(C1BB7>=0)?1:0;

ninexnine_unit ninexnine_unit_6152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC0),
				.a1(P1BD0),
				.a2(P1BE0),
				.a3(P1CC0),
				.a4(P1CD0),
				.a5(P1CE0),
				.a6(P1DC0),
				.a7(P1DD0),
				.a8(P1DE0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10BC7)
);

ninexnine_unit ninexnine_unit_6153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC1),
				.a1(P1BD1),
				.a2(P1BE1),
				.a3(P1CC1),
				.a4(P1CD1),
				.a5(P1CE1),
				.a6(P1DC1),
				.a7(P1DD1),
				.a8(P1DE1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11BC7)
);

ninexnine_unit ninexnine_unit_6154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC2),
				.a1(P1BD2),
				.a2(P1BE2),
				.a3(P1CC2),
				.a4(P1CD2),
				.a5(P1CE2),
				.a6(P1DC2),
				.a7(P1DD2),
				.a8(P1DE2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12BC7)
);

ninexnine_unit ninexnine_unit_6155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BC3),
				.a1(P1BD3),
				.a2(P1BE3),
				.a3(P1CC3),
				.a4(P1CD3),
				.a5(P1CE3),
				.a6(P1DC3),
				.a7(P1DD3),
				.a8(P1DE3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13BC7)
);

assign C1BC7=c10BC7+c11BC7+c12BC7+c13BC7;
assign A1BC7=(C1BC7>=0)?1:0;

ninexnine_unit ninexnine_unit_6156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD0),
				.a1(P1BE0),
				.a2(P1BF0),
				.a3(P1CD0),
				.a4(P1CE0),
				.a5(P1CF0),
				.a6(P1DD0),
				.a7(P1DE0),
				.a8(P1DF0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10BD7)
);

ninexnine_unit ninexnine_unit_6157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD1),
				.a1(P1BE1),
				.a2(P1BF1),
				.a3(P1CD1),
				.a4(P1CE1),
				.a5(P1CF1),
				.a6(P1DD1),
				.a7(P1DE1),
				.a8(P1DF1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11BD7)
);

ninexnine_unit ninexnine_unit_6158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD2),
				.a1(P1BE2),
				.a2(P1BF2),
				.a3(P1CD2),
				.a4(P1CE2),
				.a5(P1CF2),
				.a6(P1DD2),
				.a7(P1DE2),
				.a8(P1DF2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12BD7)
);

ninexnine_unit ninexnine_unit_6159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1BD3),
				.a1(P1BE3),
				.a2(P1BF3),
				.a3(P1CD3),
				.a4(P1CE3),
				.a5(P1CF3),
				.a6(P1DD3),
				.a7(P1DE3),
				.a8(P1DF3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13BD7)
);

assign C1BD7=c10BD7+c11BD7+c12BD7+c13BD7;
assign A1BD7=(C1BD7>=0)?1:0;

ninexnine_unit ninexnine_unit_6160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C00),
				.a1(P1C10),
				.a2(P1C20),
				.a3(P1D00),
				.a4(P1D10),
				.a5(P1D20),
				.a6(P1E00),
				.a7(P1E10),
				.a8(P1E20),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C07)
);

ninexnine_unit ninexnine_unit_6161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C01),
				.a1(P1C11),
				.a2(P1C21),
				.a3(P1D01),
				.a4(P1D11),
				.a5(P1D21),
				.a6(P1E01),
				.a7(P1E11),
				.a8(P1E21),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C07)
);

ninexnine_unit ninexnine_unit_6162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C02),
				.a1(P1C12),
				.a2(P1C22),
				.a3(P1D02),
				.a4(P1D12),
				.a5(P1D22),
				.a6(P1E02),
				.a7(P1E12),
				.a8(P1E22),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C07)
);

ninexnine_unit ninexnine_unit_6163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C03),
				.a1(P1C13),
				.a2(P1C23),
				.a3(P1D03),
				.a4(P1D13),
				.a5(P1D23),
				.a6(P1E03),
				.a7(P1E13),
				.a8(P1E23),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C07)
);

assign C1C07=c10C07+c11C07+c12C07+c13C07;
assign A1C07=(C1C07>=0)?1:0;

ninexnine_unit ninexnine_unit_6164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C10),
				.a1(P1C20),
				.a2(P1C30),
				.a3(P1D10),
				.a4(P1D20),
				.a5(P1D30),
				.a6(P1E10),
				.a7(P1E20),
				.a8(P1E30),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C17)
);

ninexnine_unit ninexnine_unit_6165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C11),
				.a1(P1C21),
				.a2(P1C31),
				.a3(P1D11),
				.a4(P1D21),
				.a5(P1D31),
				.a6(P1E11),
				.a7(P1E21),
				.a8(P1E31),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C17)
);

ninexnine_unit ninexnine_unit_6166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C12),
				.a1(P1C22),
				.a2(P1C32),
				.a3(P1D12),
				.a4(P1D22),
				.a5(P1D32),
				.a6(P1E12),
				.a7(P1E22),
				.a8(P1E32),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C17)
);

ninexnine_unit ninexnine_unit_6167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C13),
				.a1(P1C23),
				.a2(P1C33),
				.a3(P1D13),
				.a4(P1D23),
				.a5(P1D33),
				.a6(P1E13),
				.a7(P1E23),
				.a8(P1E33),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C17)
);

assign C1C17=c10C17+c11C17+c12C17+c13C17;
assign A1C17=(C1C17>=0)?1:0;

ninexnine_unit ninexnine_unit_6168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C20),
				.a1(P1C30),
				.a2(P1C40),
				.a3(P1D20),
				.a4(P1D30),
				.a5(P1D40),
				.a6(P1E20),
				.a7(P1E30),
				.a8(P1E40),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C27)
);

ninexnine_unit ninexnine_unit_6169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C21),
				.a1(P1C31),
				.a2(P1C41),
				.a3(P1D21),
				.a4(P1D31),
				.a5(P1D41),
				.a6(P1E21),
				.a7(P1E31),
				.a8(P1E41),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C27)
);

ninexnine_unit ninexnine_unit_6170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C22),
				.a1(P1C32),
				.a2(P1C42),
				.a3(P1D22),
				.a4(P1D32),
				.a5(P1D42),
				.a6(P1E22),
				.a7(P1E32),
				.a8(P1E42),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C27)
);

ninexnine_unit ninexnine_unit_6171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C23),
				.a1(P1C33),
				.a2(P1C43),
				.a3(P1D23),
				.a4(P1D33),
				.a5(P1D43),
				.a6(P1E23),
				.a7(P1E33),
				.a8(P1E43),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C27)
);

assign C1C27=c10C27+c11C27+c12C27+c13C27;
assign A1C27=(C1C27>=0)?1:0;

ninexnine_unit ninexnine_unit_6172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C30),
				.a1(P1C40),
				.a2(P1C50),
				.a3(P1D30),
				.a4(P1D40),
				.a5(P1D50),
				.a6(P1E30),
				.a7(P1E40),
				.a8(P1E50),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C37)
);

ninexnine_unit ninexnine_unit_6173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C31),
				.a1(P1C41),
				.a2(P1C51),
				.a3(P1D31),
				.a4(P1D41),
				.a5(P1D51),
				.a6(P1E31),
				.a7(P1E41),
				.a8(P1E51),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C37)
);

ninexnine_unit ninexnine_unit_6174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C32),
				.a1(P1C42),
				.a2(P1C52),
				.a3(P1D32),
				.a4(P1D42),
				.a5(P1D52),
				.a6(P1E32),
				.a7(P1E42),
				.a8(P1E52),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C37)
);

ninexnine_unit ninexnine_unit_6175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C33),
				.a1(P1C43),
				.a2(P1C53),
				.a3(P1D33),
				.a4(P1D43),
				.a5(P1D53),
				.a6(P1E33),
				.a7(P1E43),
				.a8(P1E53),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C37)
);

assign C1C37=c10C37+c11C37+c12C37+c13C37;
assign A1C37=(C1C37>=0)?1:0;

ninexnine_unit ninexnine_unit_6176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C40),
				.a1(P1C50),
				.a2(P1C60),
				.a3(P1D40),
				.a4(P1D50),
				.a5(P1D60),
				.a6(P1E40),
				.a7(P1E50),
				.a8(P1E60),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C47)
);

ninexnine_unit ninexnine_unit_6177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C41),
				.a1(P1C51),
				.a2(P1C61),
				.a3(P1D41),
				.a4(P1D51),
				.a5(P1D61),
				.a6(P1E41),
				.a7(P1E51),
				.a8(P1E61),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C47)
);

ninexnine_unit ninexnine_unit_6178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C42),
				.a1(P1C52),
				.a2(P1C62),
				.a3(P1D42),
				.a4(P1D52),
				.a5(P1D62),
				.a6(P1E42),
				.a7(P1E52),
				.a8(P1E62),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C47)
);

ninexnine_unit ninexnine_unit_6179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C43),
				.a1(P1C53),
				.a2(P1C63),
				.a3(P1D43),
				.a4(P1D53),
				.a5(P1D63),
				.a6(P1E43),
				.a7(P1E53),
				.a8(P1E63),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C47)
);

assign C1C47=c10C47+c11C47+c12C47+c13C47;
assign A1C47=(C1C47>=0)?1:0;

ninexnine_unit ninexnine_unit_6180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C50),
				.a1(P1C60),
				.a2(P1C70),
				.a3(P1D50),
				.a4(P1D60),
				.a5(P1D70),
				.a6(P1E50),
				.a7(P1E60),
				.a8(P1E70),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C57)
);

ninexnine_unit ninexnine_unit_6181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C51),
				.a1(P1C61),
				.a2(P1C71),
				.a3(P1D51),
				.a4(P1D61),
				.a5(P1D71),
				.a6(P1E51),
				.a7(P1E61),
				.a8(P1E71),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C57)
);

ninexnine_unit ninexnine_unit_6182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C52),
				.a1(P1C62),
				.a2(P1C72),
				.a3(P1D52),
				.a4(P1D62),
				.a5(P1D72),
				.a6(P1E52),
				.a7(P1E62),
				.a8(P1E72),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C57)
);

ninexnine_unit ninexnine_unit_6183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C53),
				.a1(P1C63),
				.a2(P1C73),
				.a3(P1D53),
				.a4(P1D63),
				.a5(P1D73),
				.a6(P1E53),
				.a7(P1E63),
				.a8(P1E73),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C57)
);

assign C1C57=c10C57+c11C57+c12C57+c13C57;
assign A1C57=(C1C57>=0)?1:0;

ninexnine_unit ninexnine_unit_6184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C60),
				.a1(P1C70),
				.a2(P1C80),
				.a3(P1D60),
				.a4(P1D70),
				.a5(P1D80),
				.a6(P1E60),
				.a7(P1E70),
				.a8(P1E80),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C67)
);

ninexnine_unit ninexnine_unit_6185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C61),
				.a1(P1C71),
				.a2(P1C81),
				.a3(P1D61),
				.a4(P1D71),
				.a5(P1D81),
				.a6(P1E61),
				.a7(P1E71),
				.a8(P1E81),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C67)
);

ninexnine_unit ninexnine_unit_6186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C62),
				.a1(P1C72),
				.a2(P1C82),
				.a3(P1D62),
				.a4(P1D72),
				.a5(P1D82),
				.a6(P1E62),
				.a7(P1E72),
				.a8(P1E82),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C67)
);

ninexnine_unit ninexnine_unit_6187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C63),
				.a1(P1C73),
				.a2(P1C83),
				.a3(P1D63),
				.a4(P1D73),
				.a5(P1D83),
				.a6(P1E63),
				.a7(P1E73),
				.a8(P1E83),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C67)
);

assign C1C67=c10C67+c11C67+c12C67+c13C67;
assign A1C67=(C1C67>=0)?1:0;

ninexnine_unit ninexnine_unit_6188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C70),
				.a1(P1C80),
				.a2(P1C90),
				.a3(P1D70),
				.a4(P1D80),
				.a5(P1D90),
				.a6(P1E70),
				.a7(P1E80),
				.a8(P1E90),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C77)
);

ninexnine_unit ninexnine_unit_6189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C71),
				.a1(P1C81),
				.a2(P1C91),
				.a3(P1D71),
				.a4(P1D81),
				.a5(P1D91),
				.a6(P1E71),
				.a7(P1E81),
				.a8(P1E91),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C77)
);

ninexnine_unit ninexnine_unit_6190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C72),
				.a1(P1C82),
				.a2(P1C92),
				.a3(P1D72),
				.a4(P1D82),
				.a5(P1D92),
				.a6(P1E72),
				.a7(P1E82),
				.a8(P1E92),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C77)
);

ninexnine_unit ninexnine_unit_6191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C73),
				.a1(P1C83),
				.a2(P1C93),
				.a3(P1D73),
				.a4(P1D83),
				.a5(P1D93),
				.a6(P1E73),
				.a7(P1E83),
				.a8(P1E93),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C77)
);

assign C1C77=c10C77+c11C77+c12C77+c13C77;
assign A1C77=(C1C77>=0)?1:0;

ninexnine_unit ninexnine_unit_6192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C80),
				.a1(P1C90),
				.a2(P1CA0),
				.a3(P1D80),
				.a4(P1D90),
				.a5(P1DA0),
				.a6(P1E80),
				.a7(P1E90),
				.a8(P1EA0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C87)
);

ninexnine_unit ninexnine_unit_6193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C81),
				.a1(P1C91),
				.a2(P1CA1),
				.a3(P1D81),
				.a4(P1D91),
				.a5(P1DA1),
				.a6(P1E81),
				.a7(P1E91),
				.a8(P1EA1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C87)
);

ninexnine_unit ninexnine_unit_6194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C82),
				.a1(P1C92),
				.a2(P1CA2),
				.a3(P1D82),
				.a4(P1D92),
				.a5(P1DA2),
				.a6(P1E82),
				.a7(P1E92),
				.a8(P1EA2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C87)
);

ninexnine_unit ninexnine_unit_6195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C83),
				.a1(P1C93),
				.a2(P1CA3),
				.a3(P1D83),
				.a4(P1D93),
				.a5(P1DA3),
				.a6(P1E83),
				.a7(P1E93),
				.a8(P1EA3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C87)
);

assign C1C87=c10C87+c11C87+c12C87+c13C87;
assign A1C87=(C1C87>=0)?1:0;

ninexnine_unit ninexnine_unit_6196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C90),
				.a1(P1CA0),
				.a2(P1CB0),
				.a3(P1D90),
				.a4(P1DA0),
				.a5(P1DB0),
				.a6(P1E90),
				.a7(P1EA0),
				.a8(P1EB0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10C97)
);

ninexnine_unit ninexnine_unit_6197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C91),
				.a1(P1CA1),
				.a2(P1CB1),
				.a3(P1D91),
				.a4(P1DA1),
				.a5(P1DB1),
				.a6(P1E91),
				.a7(P1EA1),
				.a8(P1EB1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11C97)
);

ninexnine_unit ninexnine_unit_6198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C92),
				.a1(P1CA2),
				.a2(P1CB2),
				.a3(P1D92),
				.a4(P1DA2),
				.a5(P1DB2),
				.a6(P1E92),
				.a7(P1EA2),
				.a8(P1EB2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12C97)
);

ninexnine_unit ninexnine_unit_6199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1C93),
				.a1(P1CA3),
				.a2(P1CB3),
				.a3(P1D93),
				.a4(P1DA3),
				.a5(P1DB3),
				.a6(P1E93),
				.a7(P1EA3),
				.a8(P1EB3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13C97)
);

assign C1C97=c10C97+c11C97+c12C97+c13C97;
assign A1C97=(C1C97>=0)?1:0;

ninexnine_unit ninexnine_unit_6200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA0),
				.a1(P1CB0),
				.a2(P1CC0),
				.a3(P1DA0),
				.a4(P1DB0),
				.a5(P1DC0),
				.a6(P1EA0),
				.a7(P1EB0),
				.a8(P1EC0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10CA7)
);

ninexnine_unit ninexnine_unit_6201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA1),
				.a1(P1CB1),
				.a2(P1CC1),
				.a3(P1DA1),
				.a4(P1DB1),
				.a5(P1DC1),
				.a6(P1EA1),
				.a7(P1EB1),
				.a8(P1EC1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11CA7)
);

ninexnine_unit ninexnine_unit_6202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA2),
				.a1(P1CB2),
				.a2(P1CC2),
				.a3(P1DA2),
				.a4(P1DB2),
				.a5(P1DC2),
				.a6(P1EA2),
				.a7(P1EB2),
				.a8(P1EC2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12CA7)
);

ninexnine_unit ninexnine_unit_6203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CA3),
				.a1(P1CB3),
				.a2(P1CC3),
				.a3(P1DA3),
				.a4(P1DB3),
				.a5(P1DC3),
				.a6(P1EA3),
				.a7(P1EB3),
				.a8(P1EC3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13CA7)
);

assign C1CA7=c10CA7+c11CA7+c12CA7+c13CA7;
assign A1CA7=(C1CA7>=0)?1:0;

ninexnine_unit ninexnine_unit_6204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB0),
				.a1(P1CC0),
				.a2(P1CD0),
				.a3(P1DB0),
				.a4(P1DC0),
				.a5(P1DD0),
				.a6(P1EB0),
				.a7(P1EC0),
				.a8(P1ED0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10CB7)
);

ninexnine_unit ninexnine_unit_6205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB1),
				.a1(P1CC1),
				.a2(P1CD1),
				.a3(P1DB1),
				.a4(P1DC1),
				.a5(P1DD1),
				.a6(P1EB1),
				.a7(P1EC1),
				.a8(P1ED1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11CB7)
);

ninexnine_unit ninexnine_unit_6206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB2),
				.a1(P1CC2),
				.a2(P1CD2),
				.a3(P1DB2),
				.a4(P1DC2),
				.a5(P1DD2),
				.a6(P1EB2),
				.a7(P1EC2),
				.a8(P1ED2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12CB7)
);

ninexnine_unit ninexnine_unit_6207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CB3),
				.a1(P1CC3),
				.a2(P1CD3),
				.a3(P1DB3),
				.a4(P1DC3),
				.a5(P1DD3),
				.a6(P1EB3),
				.a7(P1EC3),
				.a8(P1ED3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13CB7)
);

assign C1CB7=c10CB7+c11CB7+c12CB7+c13CB7;
assign A1CB7=(C1CB7>=0)?1:0;

ninexnine_unit ninexnine_unit_6208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC0),
				.a1(P1CD0),
				.a2(P1CE0),
				.a3(P1DC0),
				.a4(P1DD0),
				.a5(P1DE0),
				.a6(P1EC0),
				.a7(P1ED0),
				.a8(P1EE0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10CC7)
);

ninexnine_unit ninexnine_unit_6209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC1),
				.a1(P1CD1),
				.a2(P1CE1),
				.a3(P1DC1),
				.a4(P1DD1),
				.a5(P1DE1),
				.a6(P1EC1),
				.a7(P1ED1),
				.a8(P1EE1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11CC7)
);

ninexnine_unit ninexnine_unit_6210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC2),
				.a1(P1CD2),
				.a2(P1CE2),
				.a3(P1DC2),
				.a4(P1DD2),
				.a5(P1DE2),
				.a6(P1EC2),
				.a7(P1ED2),
				.a8(P1EE2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12CC7)
);

ninexnine_unit ninexnine_unit_6211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CC3),
				.a1(P1CD3),
				.a2(P1CE3),
				.a3(P1DC3),
				.a4(P1DD3),
				.a5(P1DE3),
				.a6(P1EC3),
				.a7(P1ED3),
				.a8(P1EE3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13CC7)
);

assign C1CC7=c10CC7+c11CC7+c12CC7+c13CC7;
assign A1CC7=(C1CC7>=0)?1:0;

ninexnine_unit ninexnine_unit_6212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD0),
				.a1(P1CE0),
				.a2(P1CF0),
				.a3(P1DD0),
				.a4(P1DE0),
				.a5(P1DF0),
				.a6(P1ED0),
				.a7(P1EE0),
				.a8(P1EF0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10CD7)
);

ninexnine_unit ninexnine_unit_6213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD1),
				.a1(P1CE1),
				.a2(P1CF1),
				.a3(P1DD1),
				.a4(P1DE1),
				.a5(P1DF1),
				.a6(P1ED1),
				.a7(P1EE1),
				.a8(P1EF1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11CD7)
);

ninexnine_unit ninexnine_unit_6214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD2),
				.a1(P1CE2),
				.a2(P1CF2),
				.a3(P1DD2),
				.a4(P1DE2),
				.a5(P1DF2),
				.a6(P1ED2),
				.a7(P1EE2),
				.a8(P1EF2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12CD7)
);

ninexnine_unit ninexnine_unit_6215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1CD3),
				.a1(P1CE3),
				.a2(P1CF3),
				.a3(P1DD3),
				.a4(P1DE3),
				.a5(P1DF3),
				.a6(P1ED3),
				.a7(P1EE3),
				.a8(P1EF3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13CD7)
);

assign C1CD7=c10CD7+c11CD7+c12CD7+c13CD7;
assign A1CD7=(C1CD7>=0)?1:0;

ninexnine_unit ninexnine_unit_6216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D00),
				.a1(P1D10),
				.a2(P1D20),
				.a3(P1E00),
				.a4(P1E10),
				.a5(P1E20),
				.a6(P1F00),
				.a7(P1F10),
				.a8(P1F20),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D07)
);

ninexnine_unit ninexnine_unit_6217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D01),
				.a1(P1D11),
				.a2(P1D21),
				.a3(P1E01),
				.a4(P1E11),
				.a5(P1E21),
				.a6(P1F01),
				.a7(P1F11),
				.a8(P1F21),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D07)
);

ninexnine_unit ninexnine_unit_6218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D02),
				.a1(P1D12),
				.a2(P1D22),
				.a3(P1E02),
				.a4(P1E12),
				.a5(P1E22),
				.a6(P1F02),
				.a7(P1F12),
				.a8(P1F22),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D07)
);

ninexnine_unit ninexnine_unit_6219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D03),
				.a1(P1D13),
				.a2(P1D23),
				.a3(P1E03),
				.a4(P1E13),
				.a5(P1E23),
				.a6(P1F03),
				.a7(P1F13),
				.a8(P1F23),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D07)
);

assign C1D07=c10D07+c11D07+c12D07+c13D07;
assign A1D07=(C1D07>=0)?1:0;

ninexnine_unit ninexnine_unit_6220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D10),
				.a1(P1D20),
				.a2(P1D30),
				.a3(P1E10),
				.a4(P1E20),
				.a5(P1E30),
				.a6(P1F10),
				.a7(P1F20),
				.a8(P1F30),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D17)
);

ninexnine_unit ninexnine_unit_6221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D11),
				.a1(P1D21),
				.a2(P1D31),
				.a3(P1E11),
				.a4(P1E21),
				.a5(P1E31),
				.a6(P1F11),
				.a7(P1F21),
				.a8(P1F31),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D17)
);

ninexnine_unit ninexnine_unit_6222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D12),
				.a1(P1D22),
				.a2(P1D32),
				.a3(P1E12),
				.a4(P1E22),
				.a5(P1E32),
				.a6(P1F12),
				.a7(P1F22),
				.a8(P1F32),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D17)
);

ninexnine_unit ninexnine_unit_6223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D13),
				.a1(P1D23),
				.a2(P1D33),
				.a3(P1E13),
				.a4(P1E23),
				.a5(P1E33),
				.a6(P1F13),
				.a7(P1F23),
				.a8(P1F33),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D17)
);

assign C1D17=c10D17+c11D17+c12D17+c13D17;
assign A1D17=(C1D17>=0)?1:0;

ninexnine_unit ninexnine_unit_6224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D20),
				.a1(P1D30),
				.a2(P1D40),
				.a3(P1E20),
				.a4(P1E30),
				.a5(P1E40),
				.a6(P1F20),
				.a7(P1F30),
				.a8(P1F40),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D27)
);

ninexnine_unit ninexnine_unit_6225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D21),
				.a1(P1D31),
				.a2(P1D41),
				.a3(P1E21),
				.a4(P1E31),
				.a5(P1E41),
				.a6(P1F21),
				.a7(P1F31),
				.a8(P1F41),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D27)
);

ninexnine_unit ninexnine_unit_6226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D22),
				.a1(P1D32),
				.a2(P1D42),
				.a3(P1E22),
				.a4(P1E32),
				.a5(P1E42),
				.a6(P1F22),
				.a7(P1F32),
				.a8(P1F42),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D27)
);

ninexnine_unit ninexnine_unit_6227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D23),
				.a1(P1D33),
				.a2(P1D43),
				.a3(P1E23),
				.a4(P1E33),
				.a5(P1E43),
				.a6(P1F23),
				.a7(P1F33),
				.a8(P1F43),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D27)
);

assign C1D27=c10D27+c11D27+c12D27+c13D27;
assign A1D27=(C1D27>=0)?1:0;

ninexnine_unit ninexnine_unit_6228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D30),
				.a1(P1D40),
				.a2(P1D50),
				.a3(P1E30),
				.a4(P1E40),
				.a5(P1E50),
				.a6(P1F30),
				.a7(P1F40),
				.a8(P1F50),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D37)
);

ninexnine_unit ninexnine_unit_6229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D31),
				.a1(P1D41),
				.a2(P1D51),
				.a3(P1E31),
				.a4(P1E41),
				.a5(P1E51),
				.a6(P1F31),
				.a7(P1F41),
				.a8(P1F51),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D37)
);

ninexnine_unit ninexnine_unit_6230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D32),
				.a1(P1D42),
				.a2(P1D52),
				.a3(P1E32),
				.a4(P1E42),
				.a5(P1E52),
				.a6(P1F32),
				.a7(P1F42),
				.a8(P1F52),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D37)
);

ninexnine_unit ninexnine_unit_6231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D33),
				.a1(P1D43),
				.a2(P1D53),
				.a3(P1E33),
				.a4(P1E43),
				.a5(P1E53),
				.a6(P1F33),
				.a7(P1F43),
				.a8(P1F53),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D37)
);

assign C1D37=c10D37+c11D37+c12D37+c13D37;
assign A1D37=(C1D37>=0)?1:0;

ninexnine_unit ninexnine_unit_6232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D40),
				.a1(P1D50),
				.a2(P1D60),
				.a3(P1E40),
				.a4(P1E50),
				.a5(P1E60),
				.a6(P1F40),
				.a7(P1F50),
				.a8(P1F60),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D47)
);

ninexnine_unit ninexnine_unit_6233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D41),
				.a1(P1D51),
				.a2(P1D61),
				.a3(P1E41),
				.a4(P1E51),
				.a5(P1E61),
				.a6(P1F41),
				.a7(P1F51),
				.a8(P1F61),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D47)
);

ninexnine_unit ninexnine_unit_6234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D42),
				.a1(P1D52),
				.a2(P1D62),
				.a3(P1E42),
				.a4(P1E52),
				.a5(P1E62),
				.a6(P1F42),
				.a7(P1F52),
				.a8(P1F62),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D47)
);

ninexnine_unit ninexnine_unit_6235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D43),
				.a1(P1D53),
				.a2(P1D63),
				.a3(P1E43),
				.a4(P1E53),
				.a5(P1E63),
				.a6(P1F43),
				.a7(P1F53),
				.a8(P1F63),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D47)
);

assign C1D47=c10D47+c11D47+c12D47+c13D47;
assign A1D47=(C1D47>=0)?1:0;

ninexnine_unit ninexnine_unit_6236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D50),
				.a1(P1D60),
				.a2(P1D70),
				.a3(P1E50),
				.a4(P1E60),
				.a5(P1E70),
				.a6(P1F50),
				.a7(P1F60),
				.a8(P1F70),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D57)
);

ninexnine_unit ninexnine_unit_6237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D51),
				.a1(P1D61),
				.a2(P1D71),
				.a3(P1E51),
				.a4(P1E61),
				.a5(P1E71),
				.a6(P1F51),
				.a7(P1F61),
				.a8(P1F71),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D57)
);

ninexnine_unit ninexnine_unit_6238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D52),
				.a1(P1D62),
				.a2(P1D72),
				.a3(P1E52),
				.a4(P1E62),
				.a5(P1E72),
				.a6(P1F52),
				.a7(P1F62),
				.a8(P1F72),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D57)
);

ninexnine_unit ninexnine_unit_6239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D53),
				.a1(P1D63),
				.a2(P1D73),
				.a3(P1E53),
				.a4(P1E63),
				.a5(P1E73),
				.a6(P1F53),
				.a7(P1F63),
				.a8(P1F73),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D57)
);

assign C1D57=c10D57+c11D57+c12D57+c13D57;
assign A1D57=(C1D57>=0)?1:0;

ninexnine_unit ninexnine_unit_6240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D60),
				.a1(P1D70),
				.a2(P1D80),
				.a3(P1E60),
				.a4(P1E70),
				.a5(P1E80),
				.a6(P1F60),
				.a7(P1F70),
				.a8(P1F80),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D67)
);

ninexnine_unit ninexnine_unit_6241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D61),
				.a1(P1D71),
				.a2(P1D81),
				.a3(P1E61),
				.a4(P1E71),
				.a5(P1E81),
				.a6(P1F61),
				.a7(P1F71),
				.a8(P1F81),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D67)
);

ninexnine_unit ninexnine_unit_6242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D62),
				.a1(P1D72),
				.a2(P1D82),
				.a3(P1E62),
				.a4(P1E72),
				.a5(P1E82),
				.a6(P1F62),
				.a7(P1F72),
				.a8(P1F82),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D67)
);

ninexnine_unit ninexnine_unit_6243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D63),
				.a1(P1D73),
				.a2(P1D83),
				.a3(P1E63),
				.a4(P1E73),
				.a5(P1E83),
				.a6(P1F63),
				.a7(P1F73),
				.a8(P1F83),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D67)
);

assign C1D67=c10D67+c11D67+c12D67+c13D67;
assign A1D67=(C1D67>=0)?1:0;

ninexnine_unit ninexnine_unit_6244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D70),
				.a1(P1D80),
				.a2(P1D90),
				.a3(P1E70),
				.a4(P1E80),
				.a5(P1E90),
				.a6(P1F70),
				.a7(P1F80),
				.a8(P1F90),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D77)
);

ninexnine_unit ninexnine_unit_6245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D71),
				.a1(P1D81),
				.a2(P1D91),
				.a3(P1E71),
				.a4(P1E81),
				.a5(P1E91),
				.a6(P1F71),
				.a7(P1F81),
				.a8(P1F91),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D77)
);

ninexnine_unit ninexnine_unit_6246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D72),
				.a1(P1D82),
				.a2(P1D92),
				.a3(P1E72),
				.a4(P1E82),
				.a5(P1E92),
				.a6(P1F72),
				.a7(P1F82),
				.a8(P1F92),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D77)
);

ninexnine_unit ninexnine_unit_6247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D73),
				.a1(P1D83),
				.a2(P1D93),
				.a3(P1E73),
				.a4(P1E83),
				.a5(P1E93),
				.a6(P1F73),
				.a7(P1F83),
				.a8(P1F93),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D77)
);

assign C1D77=c10D77+c11D77+c12D77+c13D77;
assign A1D77=(C1D77>=0)?1:0;

ninexnine_unit ninexnine_unit_6248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D80),
				.a1(P1D90),
				.a2(P1DA0),
				.a3(P1E80),
				.a4(P1E90),
				.a5(P1EA0),
				.a6(P1F80),
				.a7(P1F90),
				.a8(P1FA0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D87)
);

ninexnine_unit ninexnine_unit_6249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D81),
				.a1(P1D91),
				.a2(P1DA1),
				.a3(P1E81),
				.a4(P1E91),
				.a5(P1EA1),
				.a6(P1F81),
				.a7(P1F91),
				.a8(P1FA1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D87)
);

ninexnine_unit ninexnine_unit_6250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D82),
				.a1(P1D92),
				.a2(P1DA2),
				.a3(P1E82),
				.a4(P1E92),
				.a5(P1EA2),
				.a6(P1F82),
				.a7(P1F92),
				.a8(P1FA2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D87)
);

ninexnine_unit ninexnine_unit_6251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D83),
				.a1(P1D93),
				.a2(P1DA3),
				.a3(P1E83),
				.a4(P1E93),
				.a5(P1EA3),
				.a6(P1F83),
				.a7(P1F93),
				.a8(P1FA3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D87)
);

assign C1D87=c10D87+c11D87+c12D87+c13D87;
assign A1D87=(C1D87>=0)?1:0;

ninexnine_unit ninexnine_unit_6252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D90),
				.a1(P1DA0),
				.a2(P1DB0),
				.a3(P1E90),
				.a4(P1EA0),
				.a5(P1EB0),
				.a6(P1F90),
				.a7(P1FA0),
				.a8(P1FB0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10D97)
);

ninexnine_unit ninexnine_unit_6253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D91),
				.a1(P1DA1),
				.a2(P1DB1),
				.a3(P1E91),
				.a4(P1EA1),
				.a5(P1EB1),
				.a6(P1F91),
				.a7(P1FA1),
				.a8(P1FB1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11D97)
);

ninexnine_unit ninexnine_unit_6254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D92),
				.a1(P1DA2),
				.a2(P1DB2),
				.a3(P1E92),
				.a4(P1EA2),
				.a5(P1EB2),
				.a6(P1F92),
				.a7(P1FA2),
				.a8(P1FB2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12D97)
);

ninexnine_unit ninexnine_unit_6255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1D93),
				.a1(P1DA3),
				.a2(P1DB3),
				.a3(P1E93),
				.a4(P1EA3),
				.a5(P1EB3),
				.a6(P1F93),
				.a7(P1FA3),
				.a8(P1FB3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13D97)
);

assign C1D97=c10D97+c11D97+c12D97+c13D97;
assign A1D97=(C1D97>=0)?1:0;

ninexnine_unit ninexnine_unit_6256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA0),
				.a1(P1DB0),
				.a2(P1DC0),
				.a3(P1EA0),
				.a4(P1EB0),
				.a5(P1EC0),
				.a6(P1FA0),
				.a7(P1FB0),
				.a8(P1FC0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10DA7)
);

ninexnine_unit ninexnine_unit_6257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA1),
				.a1(P1DB1),
				.a2(P1DC1),
				.a3(P1EA1),
				.a4(P1EB1),
				.a5(P1EC1),
				.a6(P1FA1),
				.a7(P1FB1),
				.a8(P1FC1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11DA7)
);

ninexnine_unit ninexnine_unit_6258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA2),
				.a1(P1DB2),
				.a2(P1DC2),
				.a3(P1EA2),
				.a4(P1EB2),
				.a5(P1EC2),
				.a6(P1FA2),
				.a7(P1FB2),
				.a8(P1FC2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12DA7)
);

ninexnine_unit ninexnine_unit_6259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DA3),
				.a1(P1DB3),
				.a2(P1DC3),
				.a3(P1EA3),
				.a4(P1EB3),
				.a5(P1EC3),
				.a6(P1FA3),
				.a7(P1FB3),
				.a8(P1FC3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13DA7)
);

assign C1DA7=c10DA7+c11DA7+c12DA7+c13DA7;
assign A1DA7=(C1DA7>=0)?1:0;

ninexnine_unit ninexnine_unit_6260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB0),
				.a1(P1DC0),
				.a2(P1DD0),
				.a3(P1EB0),
				.a4(P1EC0),
				.a5(P1ED0),
				.a6(P1FB0),
				.a7(P1FC0),
				.a8(P1FD0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10DB7)
);

ninexnine_unit ninexnine_unit_6261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB1),
				.a1(P1DC1),
				.a2(P1DD1),
				.a3(P1EB1),
				.a4(P1EC1),
				.a5(P1ED1),
				.a6(P1FB1),
				.a7(P1FC1),
				.a8(P1FD1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11DB7)
);

ninexnine_unit ninexnine_unit_6262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB2),
				.a1(P1DC2),
				.a2(P1DD2),
				.a3(P1EB2),
				.a4(P1EC2),
				.a5(P1ED2),
				.a6(P1FB2),
				.a7(P1FC2),
				.a8(P1FD2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12DB7)
);

ninexnine_unit ninexnine_unit_6263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DB3),
				.a1(P1DC3),
				.a2(P1DD3),
				.a3(P1EB3),
				.a4(P1EC3),
				.a5(P1ED3),
				.a6(P1FB3),
				.a7(P1FC3),
				.a8(P1FD3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13DB7)
);

assign C1DB7=c10DB7+c11DB7+c12DB7+c13DB7;
assign A1DB7=(C1DB7>=0)?1:0;

ninexnine_unit ninexnine_unit_6264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC0),
				.a1(P1DD0),
				.a2(P1DE0),
				.a3(P1EC0),
				.a4(P1ED0),
				.a5(P1EE0),
				.a6(P1FC0),
				.a7(P1FD0),
				.a8(P1FE0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10DC7)
);

ninexnine_unit ninexnine_unit_6265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC1),
				.a1(P1DD1),
				.a2(P1DE1),
				.a3(P1EC1),
				.a4(P1ED1),
				.a5(P1EE1),
				.a6(P1FC1),
				.a7(P1FD1),
				.a8(P1FE1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11DC7)
);

ninexnine_unit ninexnine_unit_6266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC2),
				.a1(P1DD2),
				.a2(P1DE2),
				.a3(P1EC2),
				.a4(P1ED2),
				.a5(P1EE2),
				.a6(P1FC2),
				.a7(P1FD2),
				.a8(P1FE2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12DC7)
);

ninexnine_unit ninexnine_unit_6267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DC3),
				.a1(P1DD3),
				.a2(P1DE3),
				.a3(P1EC3),
				.a4(P1ED3),
				.a5(P1EE3),
				.a6(P1FC3),
				.a7(P1FD3),
				.a8(P1FE3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13DC7)
);

assign C1DC7=c10DC7+c11DC7+c12DC7+c13DC7;
assign A1DC7=(C1DC7>=0)?1:0;

ninexnine_unit ninexnine_unit_6268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD0),
				.a1(P1DE0),
				.a2(P1DF0),
				.a3(P1ED0),
				.a4(P1EE0),
				.a5(P1EF0),
				.a6(P1FD0),
				.a7(P1FE0),
				.a8(P1FF0),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10DD7)
);

ninexnine_unit ninexnine_unit_6269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD1),
				.a1(P1DE1),
				.a2(P1DF1),
				.a3(P1ED1),
				.a4(P1EE1),
				.a5(P1EF1),
				.a6(P1FD1),
				.a7(P1FE1),
				.a8(P1FF1),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11DD7)
);

ninexnine_unit ninexnine_unit_6270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD2),
				.a1(P1DE2),
				.a2(P1DF2),
				.a3(P1ED2),
				.a4(P1EE2),
				.a5(P1EF2),
				.a6(P1FD2),
				.a7(P1FE2),
				.a8(P1FF2),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12DD7)
);

ninexnine_unit ninexnine_unit_6271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1DD3),
				.a1(P1DE3),
				.a2(P1DF3),
				.a3(P1ED3),
				.a4(P1EE3),
				.a5(P1EF3),
				.a6(P1FD3),
				.a7(P1FE3),
				.a8(P1FF3),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13DD7)
);

assign C1DD7=c10DD7+c11DD7+c12DD7+c13DD7;
assign A1DD7=(C1DD7>=0)?1:0;

maxpool maxpool_0(
				.clk(clk),
				.rstn(rstn),
				.a0(A1000),
				.a1(A1010),
				.a2(A1100),
				.a3(A1110),
				.p(P2000)
);

maxpool maxpool_1(
				.clk(clk),
				.rstn(rstn),
				.a0(A1020),
				.a1(A1030),
				.a2(A1120),
				.a3(A1130),
				.p(P2010)
);

maxpool maxpool_2(
				.clk(clk),
				.rstn(rstn),
				.a0(A1040),
				.a1(A1050),
				.a2(A1140),
				.a3(A1150),
				.p(P2020)
);

maxpool maxpool_3(
				.clk(clk),
				.rstn(rstn),
				.a0(A1060),
				.a1(A1070),
				.a2(A1160),
				.a3(A1170),
				.p(P2030)
);

maxpool maxpool_4(
				.clk(clk),
				.rstn(rstn),
				.a0(A1080),
				.a1(A1090),
				.a2(A1180),
				.a3(A1190),
				.p(P2040)
);

maxpool maxpool_5(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A0),
				.a1(A10B0),
				.a2(A11A0),
				.a3(A11B0),
				.p(P2050)
);

maxpool maxpool_6(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C0),
				.a1(A10D0),
				.a2(A11C0),
				.a3(A11D0),
				.p(P2060)
);

maxpool maxpool_7(
				.clk(clk),
				.rstn(rstn),
				.a0(A1200),
				.a1(A1210),
				.a2(A1300),
				.a3(A1310),
				.p(P2100)
);

maxpool maxpool_8(
				.clk(clk),
				.rstn(rstn),
				.a0(A1220),
				.a1(A1230),
				.a2(A1320),
				.a3(A1330),
				.p(P2110)
);

maxpool maxpool_9(
				.clk(clk),
				.rstn(rstn),
				.a0(A1240),
				.a1(A1250),
				.a2(A1340),
				.a3(A1350),
				.p(P2120)
);

maxpool maxpool_10(
				.clk(clk),
				.rstn(rstn),
				.a0(A1260),
				.a1(A1270),
				.a2(A1360),
				.a3(A1370),
				.p(P2130)
);

maxpool maxpool_11(
				.clk(clk),
				.rstn(rstn),
				.a0(A1280),
				.a1(A1290),
				.a2(A1380),
				.a3(A1390),
				.p(P2140)
);

maxpool maxpool_12(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A0),
				.a1(A12B0),
				.a2(A13A0),
				.a3(A13B0),
				.p(P2150)
);

maxpool maxpool_13(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C0),
				.a1(A12D0),
				.a2(A13C0),
				.a3(A13D0),
				.p(P2160)
);

maxpool maxpool_14(
				.clk(clk),
				.rstn(rstn),
				.a0(A1400),
				.a1(A1410),
				.a2(A1500),
				.a3(A1510),
				.p(P2200)
);

maxpool maxpool_15(
				.clk(clk),
				.rstn(rstn),
				.a0(A1420),
				.a1(A1430),
				.a2(A1520),
				.a3(A1530),
				.p(P2210)
);

maxpool maxpool_16(
				.clk(clk),
				.rstn(rstn),
				.a0(A1440),
				.a1(A1450),
				.a2(A1540),
				.a3(A1550),
				.p(P2220)
);

maxpool maxpool_17(
				.clk(clk),
				.rstn(rstn),
				.a0(A1460),
				.a1(A1470),
				.a2(A1560),
				.a3(A1570),
				.p(P2230)
);

maxpool maxpool_18(
				.clk(clk),
				.rstn(rstn),
				.a0(A1480),
				.a1(A1490),
				.a2(A1580),
				.a3(A1590),
				.p(P2240)
);

maxpool maxpool_19(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A0),
				.a1(A14B0),
				.a2(A15A0),
				.a3(A15B0),
				.p(P2250)
);

maxpool maxpool_20(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C0),
				.a1(A14D0),
				.a2(A15C0),
				.a3(A15D0),
				.p(P2260)
);

maxpool maxpool_21(
				.clk(clk),
				.rstn(rstn),
				.a0(A1600),
				.a1(A1610),
				.a2(A1700),
				.a3(A1710),
				.p(P2300)
);

maxpool maxpool_22(
				.clk(clk),
				.rstn(rstn),
				.a0(A1620),
				.a1(A1630),
				.a2(A1720),
				.a3(A1730),
				.p(P2310)
);

maxpool maxpool_23(
				.clk(clk),
				.rstn(rstn),
				.a0(A1640),
				.a1(A1650),
				.a2(A1740),
				.a3(A1750),
				.p(P2320)
);

maxpool maxpool_24(
				.clk(clk),
				.rstn(rstn),
				.a0(A1660),
				.a1(A1670),
				.a2(A1760),
				.a3(A1770),
				.p(P2330)
);

maxpool maxpool_25(
				.clk(clk),
				.rstn(rstn),
				.a0(A1680),
				.a1(A1690),
				.a2(A1780),
				.a3(A1790),
				.p(P2340)
);

maxpool maxpool_26(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A0),
				.a1(A16B0),
				.a2(A17A0),
				.a3(A17B0),
				.p(P2350)
);

maxpool maxpool_27(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C0),
				.a1(A16D0),
				.a2(A17C0),
				.a3(A17D0),
				.p(P2360)
);

maxpool maxpool_28(
				.clk(clk),
				.rstn(rstn),
				.a0(A1800),
				.a1(A1810),
				.a2(A1900),
				.a3(A1910),
				.p(P2400)
);

maxpool maxpool_29(
				.clk(clk),
				.rstn(rstn),
				.a0(A1820),
				.a1(A1830),
				.a2(A1920),
				.a3(A1930),
				.p(P2410)
);

maxpool maxpool_30(
				.clk(clk),
				.rstn(rstn),
				.a0(A1840),
				.a1(A1850),
				.a2(A1940),
				.a3(A1950),
				.p(P2420)
);

maxpool maxpool_31(
				.clk(clk),
				.rstn(rstn),
				.a0(A1860),
				.a1(A1870),
				.a2(A1960),
				.a3(A1970),
				.p(P2430)
);

maxpool maxpool_32(
				.clk(clk),
				.rstn(rstn),
				.a0(A1880),
				.a1(A1890),
				.a2(A1980),
				.a3(A1990),
				.p(P2440)
);

maxpool maxpool_33(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A0),
				.a1(A18B0),
				.a2(A19A0),
				.a3(A19B0),
				.p(P2450)
);

maxpool maxpool_34(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C0),
				.a1(A18D0),
				.a2(A19C0),
				.a3(A19D0),
				.p(P2460)
);

maxpool maxpool_35(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A00),
				.a1(A1A10),
				.a2(A1B00),
				.a3(A1B10),
				.p(P2500)
);

maxpool maxpool_36(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A20),
				.a1(A1A30),
				.a2(A1B20),
				.a3(A1B30),
				.p(P2510)
);

maxpool maxpool_37(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A40),
				.a1(A1A50),
				.a2(A1B40),
				.a3(A1B50),
				.p(P2520)
);

maxpool maxpool_38(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A60),
				.a1(A1A70),
				.a2(A1B60),
				.a3(A1B70),
				.p(P2530)
);

maxpool maxpool_39(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A80),
				.a1(A1A90),
				.a2(A1B80),
				.a3(A1B90),
				.p(P2540)
);

maxpool maxpool_40(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA0),
				.a1(A1AB0),
				.a2(A1BA0),
				.a3(A1BB0),
				.p(P2550)
);

maxpool maxpool_41(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC0),
				.a1(A1AD0),
				.a2(A1BC0),
				.a3(A1BD0),
				.p(P2560)
);

maxpool maxpool_42(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C00),
				.a1(A1C10),
				.a2(A1D00),
				.a3(A1D10),
				.p(P2600)
);

maxpool maxpool_43(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C20),
				.a1(A1C30),
				.a2(A1D20),
				.a3(A1D30),
				.p(P2610)
);

maxpool maxpool_44(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C40),
				.a1(A1C50),
				.a2(A1D40),
				.a3(A1D50),
				.p(P2620)
);

maxpool maxpool_45(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C60),
				.a1(A1C70),
				.a2(A1D60),
				.a3(A1D70),
				.p(P2630)
);

maxpool maxpool_46(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C80),
				.a1(A1C90),
				.a2(A1D80),
				.a3(A1D90),
				.p(P2640)
);

maxpool maxpool_47(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA0),
				.a1(A1CB0),
				.a2(A1DA0),
				.a3(A1DB0),
				.p(P2650)
);

maxpool maxpool_48(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC0),
				.a1(A1CD0),
				.a2(A1DC0),
				.a3(A1DD0),
				.p(P2660)
);

maxpool maxpool_49(
				.clk(clk),
				.rstn(rstn),
				.a0(A1001),
				.a1(A1011),
				.a2(A1101),
				.a3(A1111),
				.p(P2001)
);

maxpool maxpool_50(
				.clk(clk),
				.rstn(rstn),
				.a0(A1021),
				.a1(A1031),
				.a2(A1121),
				.a3(A1131),
				.p(P2011)
);

maxpool maxpool_51(
				.clk(clk),
				.rstn(rstn),
				.a0(A1041),
				.a1(A1051),
				.a2(A1141),
				.a3(A1151),
				.p(P2021)
);

maxpool maxpool_52(
				.clk(clk),
				.rstn(rstn),
				.a0(A1061),
				.a1(A1071),
				.a2(A1161),
				.a3(A1171),
				.p(P2031)
);

maxpool maxpool_53(
				.clk(clk),
				.rstn(rstn),
				.a0(A1081),
				.a1(A1091),
				.a2(A1181),
				.a3(A1191),
				.p(P2041)
);

maxpool maxpool_54(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A1),
				.a1(A10B1),
				.a2(A11A1),
				.a3(A11B1),
				.p(P2051)
);

maxpool maxpool_55(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C1),
				.a1(A10D1),
				.a2(A11C1),
				.a3(A11D1),
				.p(P2061)
);

maxpool maxpool_56(
				.clk(clk),
				.rstn(rstn),
				.a0(A1201),
				.a1(A1211),
				.a2(A1301),
				.a3(A1311),
				.p(P2101)
);

maxpool maxpool_57(
				.clk(clk),
				.rstn(rstn),
				.a0(A1221),
				.a1(A1231),
				.a2(A1321),
				.a3(A1331),
				.p(P2111)
);

maxpool maxpool_58(
				.clk(clk),
				.rstn(rstn),
				.a0(A1241),
				.a1(A1251),
				.a2(A1341),
				.a3(A1351),
				.p(P2121)
);

maxpool maxpool_59(
				.clk(clk),
				.rstn(rstn),
				.a0(A1261),
				.a1(A1271),
				.a2(A1361),
				.a3(A1371),
				.p(P2131)
);

maxpool maxpool_60(
				.clk(clk),
				.rstn(rstn),
				.a0(A1281),
				.a1(A1291),
				.a2(A1381),
				.a3(A1391),
				.p(P2141)
);

maxpool maxpool_61(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A1),
				.a1(A12B1),
				.a2(A13A1),
				.a3(A13B1),
				.p(P2151)
);

maxpool maxpool_62(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C1),
				.a1(A12D1),
				.a2(A13C1),
				.a3(A13D1),
				.p(P2161)
);

maxpool maxpool_63(
				.clk(clk),
				.rstn(rstn),
				.a0(A1401),
				.a1(A1411),
				.a2(A1501),
				.a3(A1511),
				.p(P2201)
);

maxpool maxpool_64(
				.clk(clk),
				.rstn(rstn),
				.a0(A1421),
				.a1(A1431),
				.a2(A1521),
				.a3(A1531),
				.p(P2211)
);

maxpool maxpool_65(
				.clk(clk),
				.rstn(rstn),
				.a0(A1441),
				.a1(A1451),
				.a2(A1541),
				.a3(A1551),
				.p(P2221)
);

maxpool maxpool_66(
				.clk(clk),
				.rstn(rstn),
				.a0(A1461),
				.a1(A1471),
				.a2(A1561),
				.a3(A1571),
				.p(P2231)
);

maxpool maxpool_67(
				.clk(clk),
				.rstn(rstn),
				.a0(A1481),
				.a1(A1491),
				.a2(A1581),
				.a3(A1591),
				.p(P2241)
);

maxpool maxpool_68(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A1),
				.a1(A14B1),
				.a2(A15A1),
				.a3(A15B1),
				.p(P2251)
);

maxpool maxpool_69(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C1),
				.a1(A14D1),
				.a2(A15C1),
				.a3(A15D1),
				.p(P2261)
);

maxpool maxpool_70(
				.clk(clk),
				.rstn(rstn),
				.a0(A1601),
				.a1(A1611),
				.a2(A1701),
				.a3(A1711),
				.p(P2301)
);

maxpool maxpool_71(
				.clk(clk),
				.rstn(rstn),
				.a0(A1621),
				.a1(A1631),
				.a2(A1721),
				.a3(A1731),
				.p(P2311)
);

maxpool maxpool_72(
				.clk(clk),
				.rstn(rstn),
				.a0(A1641),
				.a1(A1651),
				.a2(A1741),
				.a3(A1751),
				.p(P2321)
);

maxpool maxpool_73(
				.clk(clk),
				.rstn(rstn),
				.a0(A1661),
				.a1(A1671),
				.a2(A1761),
				.a3(A1771),
				.p(P2331)
);

maxpool maxpool_74(
				.clk(clk),
				.rstn(rstn),
				.a0(A1681),
				.a1(A1691),
				.a2(A1781),
				.a3(A1791),
				.p(P2341)
);

maxpool maxpool_75(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A1),
				.a1(A16B1),
				.a2(A17A1),
				.a3(A17B1),
				.p(P2351)
);

maxpool maxpool_76(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C1),
				.a1(A16D1),
				.a2(A17C1),
				.a3(A17D1),
				.p(P2361)
);

maxpool maxpool_77(
				.clk(clk),
				.rstn(rstn),
				.a0(A1801),
				.a1(A1811),
				.a2(A1901),
				.a3(A1911),
				.p(P2401)
);

maxpool maxpool_78(
				.clk(clk),
				.rstn(rstn),
				.a0(A1821),
				.a1(A1831),
				.a2(A1921),
				.a3(A1931),
				.p(P2411)
);

maxpool maxpool_79(
				.clk(clk),
				.rstn(rstn),
				.a0(A1841),
				.a1(A1851),
				.a2(A1941),
				.a3(A1951),
				.p(P2421)
);

maxpool maxpool_80(
				.clk(clk),
				.rstn(rstn),
				.a0(A1861),
				.a1(A1871),
				.a2(A1961),
				.a3(A1971),
				.p(P2431)
);

maxpool maxpool_81(
				.clk(clk),
				.rstn(rstn),
				.a0(A1881),
				.a1(A1891),
				.a2(A1981),
				.a3(A1991),
				.p(P2441)
);

maxpool maxpool_82(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A1),
				.a1(A18B1),
				.a2(A19A1),
				.a3(A19B1),
				.p(P2451)
);

maxpool maxpool_83(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C1),
				.a1(A18D1),
				.a2(A19C1),
				.a3(A19D1),
				.p(P2461)
);

maxpool maxpool_84(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A01),
				.a1(A1A11),
				.a2(A1B01),
				.a3(A1B11),
				.p(P2501)
);

maxpool maxpool_85(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A21),
				.a1(A1A31),
				.a2(A1B21),
				.a3(A1B31),
				.p(P2511)
);

maxpool maxpool_86(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A41),
				.a1(A1A51),
				.a2(A1B41),
				.a3(A1B51),
				.p(P2521)
);

maxpool maxpool_87(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A61),
				.a1(A1A71),
				.a2(A1B61),
				.a3(A1B71),
				.p(P2531)
);

maxpool maxpool_88(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A81),
				.a1(A1A91),
				.a2(A1B81),
				.a3(A1B91),
				.p(P2541)
);

maxpool maxpool_89(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA1),
				.a1(A1AB1),
				.a2(A1BA1),
				.a3(A1BB1),
				.p(P2551)
);

maxpool maxpool_90(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC1),
				.a1(A1AD1),
				.a2(A1BC1),
				.a3(A1BD1),
				.p(P2561)
);

maxpool maxpool_91(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C01),
				.a1(A1C11),
				.a2(A1D01),
				.a3(A1D11),
				.p(P2601)
);

maxpool maxpool_92(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C21),
				.a1(A1C31),
				.a2(A1D21),
				.a3(A1D31),
				.p(P2611)
);

maxpool maxpool_93(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C41),
				.a1(A1C51),
				.a2(A1D41),
				.a3(A1D51),
				.p(P2621)
);

maxpool maxpool_94(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C61),
				.a1(A1C71),
				.a2(A1D61),
				.a3(A1D71),
				.p(P2631)
);

maxpool maxpool_95(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C81),
				.a1(A1C91),
				.a2(A1D81),
				.a3(A1D91),
				.p(P2641)
);

maxpool maxpool_96(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA1),
				.a1(A1CB1),
				.a2(A1DA1),
				.a3(A1DB1),
				.p(P2651)
);

maxpool maxpool_97(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC1),
				.a1(A1CD1),
				.a2(A1DC1),
				.a3(A1DD1),
				.p(P2661)
);

maxpool maxpool_98(
				.clk(clk),
				.rstn(rstn),
				.a0(A1002),
				.a1(A1012),
				.a2(A1102),
				.a3(A1112),
				.p(P2002)
);

maxpool maxpool_99(
				.clk(clk),
				.rstn(rstn),
				.a0(A1022),
				.a1(A1032),
				.a2(A1122),
				.a3(A1132),
				.p(P2012)
);

maxpool maxpool_100(
				.clk(clk),
				.rstn(rstn),
				.a0(A1042),
				.a1(A1052),
				.a2(A1142),
				.a3(A1152),
				.p(P2022)
);

maxpool maxpool_101(
				.clk(clk),
				.rstn(rstn),
				.a0(A1062),
				.a1(A1072),
				.a2(A1162),
				.a3(A1172),
				.p(P2032)
);

maxpool maxpool_102(
				.clk(clk),
				.rstn(rstn),
				.a0(A1082),
				.a1(A1092),
				.a2(A1182),
				.a3(A1192),
				.p(P2042)
);

maxpool maxpool_103(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A2),
				.a1(A10B2),
				.a2(A11A2),
				.a3(A11B2),
				.p(P2052)
);

maxpool maxpool_104(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C2),
				.a1(A10D2),
				.a2(A11C2),
				.a3(A11D2),
				.p(P2062)
);

maxpool maxpool_105(
				.clk(clk),
				.rstn(rstn),
				.a0(A1202),
				.a1(A1212),
				.a2(A1302),
				.a3(A1312),
				.p(P2102)
);

maxpool maxpool_106(
				.clk(clk),
				.rstn(rstn),
				.a0(A1222),
				.a1(A1232),
				.a2(A1322),
				.a3(A1332),
				.p(P2112)
);

maxpool maxpool_107(
				.clk(clk),
				.rstn(rstn),
				.a0(A1242),
				.a1(A1252),
				.a2(A1342),
				.a3(A1352),
				.p(P2122)
);

maxpool maxpool_108(
				.clk(clk),
				.rstn(rstn),
				.a0(A1262),
				.a1(A1272),
				.a2(A1362),
				.a3(A1372),
				.p(P2132)
);

maxpool maxpool_109(
				.clk(clk),
				.rstn(rstn),
				.a0(A1282),
				.a1(A1292),
				.a2(A1382),
				.a3(A1392),
				.p(P2142)
);

maxpool maxpool_110(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A2),
				.a1(A12B2),
				.a2(A13A2),
				.a3(A13B2),
				.p(P2152)
);

maxpool maxpool_111(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C2),
				.a1(A12D2),
				.a2(A13C2),
				.a3(A13D2),
				.p(P2162)
);

maxpool maxpool_112(
				.clk(clk),
				.rstn(rstn),
				.a0(A1402),
				.a1(A1412),
				.a2(A1502),
				.a3(A1512),
				.p(P2202)
);

maxpool maxpool_113(
				.clk(clk),
				.rstn(rstn),
				.a0(A1422),
				.a1(A1432),
				.a2(A1522),
				.a3(A1532),
				.p(P2212)
);

maxpool maxpool_114(
				.clk(clk),
				.rstn(rstn),
				.a0(A1442),
				.a1(A1452),
				.a2(A1542),
				.a3(A1552),
				.p(P2222)
);

maxpool maxpool_115(
				.clk(clk),
				.rstn(rstn),
				.a0(A1462),
				.a1(A1472),
				.a2(A1562),
				.a3(A1572),
				.p(P2232)
);

maxpool maxpool_116(
				.clk(clk),
				.rstn(rstn),
				.a0(A1482),
				.a1(A1492),
				.a2(A1582),
				.a3(A1592),
				.p(P2242)
);

maxpool maxpool_117(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A2),
				.a1(A14B2),
				.a2(A15A2),
				.a3(A15B2),
				.p(P2252)
);

maxpool maxpool_118(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C2),
				.a1(A14D2),
				.a2(A15C2),
				.a3(A15D2),
				.p(P2262)
);

maxpool maxpool_119(
				.clk(clk),
				.rstn(rstn),
				.a0(A1602),
				.a1(A1612),
				.a2(A1702),
				.a3(A1712),
				.p(P2302)
);

maxpool maxpool_120(
				.clk(clk),
				.rstn(rstn),
				.a0(A1622),
				.a1(A1632),
				.a2(A1722),
				.a3(A1732),
				.p(P2312)
);

maxpool maxpool_121(
				.clk(clk),
				.rstn(rstn),
				.a0(A1642),
				.a1(A1652),
				.a2(A1742),
				.a3(A1752),
				.p(P2322)
);

maxpool maxpool_122(
				.clk(clk),
				.rstn(rstn),
				.a0(A1662),
				.a1(A1672),
				.a2(A1762),
				.a3(A1772),
				.p(P2332)
);

maxpool maxpool_123(
				.clk(clk),
				.rstn(rstn),
				.a0(A1682),
				.a1(A1692),
				.a2(A1782),
				.a3(A1792),
				.p(P2342)
);

maxpool maxpool_124(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A2),
				.a1(A16B2),
				.a2(A17A2),
				.a3(A17B2),
				.p(P2352)
);

maxpool maxpool_125(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C2),
				.a1(A16D2),
				.a2(A17C2),
				.a3(A17D2),
				.p(P2362)
);

maxpool maxpool_126(
				.clk(clk),
				.rstn(rstn),
				.a0(A1802),
				.a1(A1812),
				.a2(A1902),
				.a3(A1912),
				.p(P2402)
);

maxpool maxpool_127(
				.clk(clk),
				.rstn(rstn),
				.a0(A1822),
				.a1(A1832),
				.a2(A1922),
				.a3(A1932),
				.p(P2412)
);

maxpool maxpool_128(
				.clk(clk),
				.rstn(rstn),
				.a0(A1842),
				.a1(A1852),
				.a2(A1942),
				.a3(A1952),
				.p(P2422)
);

maxpool maxpool_129(
				.clk(clk),
				.rstn(rstn),
				.a0(A1862),
				.a1(A1872),
				.a2(A1962),
				.a3(A1972),
				.p(P2432)
);

maxpool maxpool_130(
				.clk(clk),
				.rstn(rstn),
				.a0(A1882),
				.a1(A1892),
				.a2(A1982),
				.a3(A1992),
				.p(P2442)
);

maxpool maxpool_131(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A2),
				.a1(A18B2),
				.a2(A19A2),
				.a3(A19B2),
				.p(P2452)
);

maxpool maxpool_132(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C2),
				.a1(A18D2),
				.a2(A19C2),
				.a3(A19D2),
				.p(P2462)
);

maxpool maxpool_133(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A02),
				.a1(A1A12),
				.a2(A1B02),
				.a3(A1B12),
				.p(P2502)
);

maxpool maxpool_134(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A22),
				.a1(A1A32),
				.a2(A1B22),
				.a3(A1B32),
				.p(P2512)
);

maxpool maxpool_135(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A42),
				.a1(A1A52),
				.a2(A1B42),
				.a3(A1B52),
				.p(P2522)
);

maxpool maxpool_136(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A62),
				.a1(A1A72),
				.a2(A1B62),
				.a3(A1B72),
				.p(P2532)
);

maxpool maxpool_137(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A82),
				.a1(A1A92),
				.a2(A1B82),
				.a3(A1B92),
				.p(P2542)
);

maxpool maxpool_138(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA2),
				.a1(A1AB2),
				.a2(A1BA2),
				.a3(A1BB2),
				.p(P2552)
);

maxpool maxpool_139(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC2),
				.a1(A1AD2),
				.a2(A1BC2),
				.a3(A1BD2),
				.p(P2562)
);

maxpool maxpool_140(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C02),
				.a1(A1C12),
				.a2(A1D02),
				.a3(A1D12),
				.p(P2602)
);

maxpool maxpool_141(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C22),
				.a1(A1C32),
				.a2(A1D22),
				.a3(A1D32),
				.p(P2612)
);

maxpool maxpool_142(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C42),
				.a1(A1C52),
				.a2(A1D42),
				.a3(A1D52),
				.p(P2622)
);

maxpool maxpool_143(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C62),
				.a1(A1C72),
				.a2(A1D62),
				.a3(A1D72),
				.p(P2632)
);

maxpool maxpool_144(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C82),
				.a1(A1C92),
				.a2(A1D82),
				.a3(A1D92),
				.p(P2642)
);

maxpool maxpool_145(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA2),
				.a1(A1CB2),
				.a2(A1DA2),
				.a3(A1DB2),
				.p(P2652)
);

maxpool maxpool_146(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC2),
				.a1(A1CD2),
				.a2(A1DC2),
				.a3(A1DD2),
				.p(P2662)
);

maxpool maxpool_147(
				.clk(clk),
				.rstn(rstn),
				.a0(A1003),
				.a1(A1013),
				.a2(A1103),
				.a3(A1113),
				.p(P2003)
);

maxpool maxpool_148(
				.clk(clk),
				.rstn(rstn),
				.a0(A1023),
				.a1(A1033),
				.a2(A1123),
				.a3(A1133),
				.p(P2013)
);

maxpool maxpool_149(
				.clk(clk),
				.rstn(rstn),
				.a0(A1043),
				.a1(A1053),
				.a2(A1143),
				.a3(A1153),
				.p(P2023)
);

maxpool maxpool_150(
				.clk(clk),
				.rstn(rstn),
				.a0(A1063),
				.a1(A1073),
				.a2(A1163),
				.a3(A1173),
				.p(P2033)
);

maxpool maxpool_151(
				.clk(clk),
				.rstn(rstn),
				.a0(A1083),
				.a1(A1093),
				.a2(A1183),
				.a3(A1193),
				.p(P2043)
);

maxpool maxpool_152(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A3),
				.a1(A10B3),
				.a2(A11A3),
				.a3(A11B3),
				.p(P2053)
);

maxpool maxpool_153(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C3),
				.a1(A10D3),
				.a2(A11C3),
				.a3(A11D3),
				.p(P2063)
);

maxpool maxpool_154(
				.clk(clk),
				.rstn(rstn),
				.a0(A1203),
				.a1(A1213),
				.a2(A1303),
				.a3(A1313),
				.p(P2103)
);

maxpool maxpool_155(
				.clk(clk),
				.rstn(rstn),
				.a0(A1223),
				.a1(A1233),
				.a2(A1323),
				.a3(A1333),
				.p(P2113)
);

maxpool maxpool_156(
				.clk(clk),
				.rstn(rstn),
				.a0(A1243),
				.a1(A1253),
				.a2(A1343),
				.a3(A1353),
				.p(P2123)
);

maxpool maxpool_157(
				.clk(clk),
				.rstn(rstn),
				.a0(A1263),
				.a1(A1273),
				.a2(A1363),
				.a3(A1373),
				.p(P2133)
);

maxpool maxpool_158(
				.clk(clk),
				.rstn(rstn),
				.a0(A1283),
				.a1(A1293),
				.a2(A1383),
				.a3(A1393),
				.p(P2143)
);

maxpool maxpool_159(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A3),
				.a1(A12B3),
				.a2(A13A3),
				.a3(A13B3),
				.p(P2153)
);

maxpool maxpool_160(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C3),
				.a1(A12D3),
				.a2(A13C3),
				.a3(A13D3),
				.p(P2163)
);

maxpool maxpool_161(
				.clk(clk),
				.rstn(rstn),
				.a0(A1403),
				.a1(A1413),
				.a2(A1503),
				.a3(A1513),
				.p(P2203)
);

maxpool maxpool_162(
				.clk(clk),
				.rstn(rstn),
				.a0(A1423),
				.a1(A1433),
				.a2(A1523),
				.a3(A1533),
				.p(P2213)
);

maxpool maxpool_163(
				.clk(clk),
				.rstn(rstn),
				.a0(A1443),
				.a1(A1453),
				.a2(A1543),
				.a3(A1553),
				.p(P2223)
);

maxpool maxpool_164(
				.clk(clk),
				.rstn(rstn),
				.a0(A1463),
				.a1(A1473),
				.a2(A1563),
				.a3(A1573),
				.p(P2233)
);

maxpool maxpool_165(
				.clk(clk),
				.rstn(rstn),
				.a0(A1483),
				.a1(A1493),
				.a2(A1583),
				.a3(A1593),
				.p(P2243)
);

maxpool maxpool_166(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A3),
				.a1(A14B3),
				.a2(A15A3),
				.a3(A15B3),
				.p(P2253)
);

maxpool maxpool_167(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C3),
				.a1(A14D3),
				.a2(A15C3),
				.a3(A15D3),
				.p(P2263)
);

maxpool maxpool_168(
				.clk(clk),
				.rstn(rstn),
				.a0(A1603),
				.a1(A1613),
				.a2(A1703),
				.a3(A1713),
				.p(P2303)
);

maxpool maxpool_169(
				.clk(clk),
				.rstn(rstn),
				.a0(A1623),
				.a1(A1633),
				.a2(A1723),
				.a3(A1733),
				.p(P2313)
);

maxpool maxpool_170(
				.clk(clk),
				.rstn(rstn),
				.a0(A1643),
				.a1(A1653),
				.a2(A1743),
				.a3(A1753),
				.p(P2323)
);

maxpool maxpool_171(
				.clk(clk),
				.rstn(rstn),
				.a0(A1663),
				.a1(A1673),
				.a2(A1763),
				.a3(A1773),
				.p(P2333)
);

maxpool maxpool_172(
				.clk(clk),
				.rstn(rstn),
				.a0(A1683),
				.a1(A1693),
				.a2(A1783),
				.a3(A1793),
				.p(P2343)
);

maxpool maxpool_173(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A3),
				.a1(A16B3),
				.a2(A17A3),
				.a3(A17B3),
				.p(P2353)
);

maxpool maxpool_174(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C3),
				.a1(A16D3),
				.a2(A17C3),
				.a3(A17D3),
				.p(P2363)
);

maxpool maxpool_175(
				.clk(clk),
				.rstn(rstn),
				.a0(A1803),
				.a1(A1813),
				.a2(A1903),
				.a3(A1913),
				.p(P2403)
);

maxpool maxpool_176(
				.clk(clk),
				.rstn(rstn),
				.a0(A1823),
				.a1(A1833),
				.a2(A1923),
				.a3(A1933),
				.p(P2413)
);

maxpool maxpool_177(
				.clk(clk),
				.rstn(rstn),
				.a0(A1843),
				.a1(A1853),
				.a2(A1943),
				.a3(A1953),
				.p(P2423)
);

maxpool maxpool_178(
				.clk(clk),
				.rstn(rstn),
				.a0(A1863),
				.a1(A1873),
				.a2(A1963),
				.a3(A1973),
				.p(P2433)
);

maxpool maxpool_179(
				.clk(clk),
				.rstn(rstn),
				.a0(A1883),
				.a1(A1893),
				.a2(A1983),
				.a3(A1993),
				.p(P2443)
);

maxpool maxpool_180(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A3),
				.a1(A18B3),
				.a2(A19A3),
				.a3(A19B3),
				.p(P2453)
);

maxpool maxpool_181(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C3),
				.a1(A18D3),
				.a2(A19C3),
				.a3(A19D3),
				.p(P2463)
);

maxpool maxpool_182(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A03),
				.a1(A1A13),
				.a2(A1B03),
				.a3(A1B13),
				.p(P2503)
);

maxpool maxpool_183(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A23),
				.a1(A1A33),
				.a2(A1B23),
				.a3(A1B33),
				.p(P2513)
);

maxpool maxpool_184(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A43),
				.a1(A1A53),
				.a2(A1B43),
				.a3(A1B53),
				.p(P2523)
);

maxpool maxpool_185(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A63),
				.a1(A1A73),
				.a2(A1B63),
				.a3(A1B73),
				.p(P2533)
);

maxpool maxpool_186(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A83),
				.a1(A1A93),
				.a2(A1B83),
				.a3(A1B93),
				.p(P2543)
);

maxpool maxpool_187(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA3),
				.a1(A1AB3),
				.a2(A1BA3),
				.a3(A1BB3),
				.p(P2553)
);

maxpool maxpool_188(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC3),
				.a1(A1AD3),
				.a2(A1BC3),
				.a3(A1BD3),
				.p(P2563)
);

maxpool maxpool_189(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C03),
				.a1(A1C13),
				.a2(A1D03),
				.a3(A1D13),
				.p(P2603)
);

maxpool maxpool_190(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C23),
				.a1(A1C33),
				.a2(A1D23),
				.a3(A1D33),
				.p(P2613)
);

maxpool maxpool_191(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C43),
				.a1(A1C53),
				.a2(A1D43),
				.a3(A1D53),
				.p(P2623)
);

maxpool maxpool_192(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C63),
				.a1(A1C73),
				.a2(A1D63),
				.a3(A1D73),
				.p(P2633)
);

maxpool maxpool_193(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C83),
				.a1(A1C93),
				.a2(A1D83),
				.a3(A1D93),
				.p(P2643)
);

maxpool maxpool_194(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA3),
				.a1(A1CB3),
				.a2(A1DA3),
				.a3(A1DB3),
				.p(P2653)
);

maxpool maxpool_195(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC3),
				.a1(A1CD3),
				.a2(A1DC3),
				.a3(A1DD3),
				.p(P2663)
);

maxpool maxpool_196(
				.clk(clk),
				.rstn(rstn),
				.a0(A1004),
				.a1(A1014),
				.a2(A1104),
				.a3(A1114),
				.p(P2004)
);

maxpool maxpool_197(
				.clk(clk),
				.rstn(rstn),
				.a0(A1024),
				.a1(A1034),
				.a2(A1124),
				.a3(A1134),
				.p(P2014)
);

maxpool maxpool_198(
				.clk(clk),
				.rstn(rstn),
				.a0(A1044),
				.a1(A1054),
				.a2(A1144),
				.a3(A1154),
				.p(P2024)
);

maxpool maxpool_199(
				.clk(clk),
				.rstn(rstn),
				.a0(A1064),
				.a1(A1074),
				.a2(A1164),
				.a3(A1174),
				.p(P2034)
);

maxpool maxpool_200(
				.clk(clk),
				.rstn(rstn),
				.a0(A1084),
				.a1(A1094),
				.a2(A1184),
				.a3(A1194),
				.p(P2044)
);

maxpool maxpool_201(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A4),
				.a1(A10B4),
				.a2(A11A4),
				.a3(A11B4),
				.p(P2054)
);

maxpool maxpool_202(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C4),
				.a1(A10D4),
				.a2(A11C4),
				.a3(A11D4),
				.p(P2064)
);

maxpool maxpool_203(
				.clk(clk),
				.rstn(rstn),
				.a0(A1204),
				.a1(A1214),
				.a2(A1304),
				.a3(A1314),
				.p(P2104)
);

maxpool maxpool_204(
				.clk(clk),
				.rstn(rstn),
				.a0(A1224),
				.a1(A1234),
				.a2(A1324),
				.a3(A1334),
				.p(P2114)
);

maxpool maxpool_205(
				.clk(clk),
				.rstn(rstn),
				.a0(A1244),
				.a1(A1254),
				.a2(A1344),
				.a3(A1354),
				.p(P2124)
);

maxpool maxpool_206(
				.clk(clk),
				.rstn(rstn),
				.a0(A1264),
				.a1(A1274),
				.a2(A1364),
				.a3(A1374),
				.p(P2134)
);

maxpool maxpool_207(
				.clk(clk),
				.rstn(rstn),
				.a0(A1284),
				.a1(A1294),
				.a2(A1384),
				.a3(A1394),
				.p(P2144)
);

maxpool maxpool_208(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A4),
				.a1(A12B4),
				.a2(A13A4),
				.a3(A13B4),
				.p(P2154)
);

maxpool maxpool_209(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C4),
				.a1(A12D4),
				.a2(A13C4),
				.a3(A13D4),
				.p(P2164)
);

maxpool maxpool_210(
				.clk(clk),
				.rstn(rstn),
				.a0(A1404),
				.a1(A1414),
				.a2(A1504),
				.a3(A1514),
				.p(P2204)
);

maxpool maxpool_211(
				.clk(clk),
				.rstn(rstn),
				.a0(A1424),
				.a1(A1434),
				.a2(A1524),
				.a3(A1534),
				.p(P2214)
);

maxpool maxpool_212(
				.clk(clk),
				.rstn(rstn),
				.a0(A1444),
				.a1(A1454),
				.a2(A1544),
				.a3(A1554),
				.p(P2224)
);

maxpool maxpool_213(
				.clk(clk),
				.rstn(rstn),
				.a0(A1464),
				.a1(A1474),
				.a2(A1564),
				.a3(A1574),
				.p(P2234)
);

maxpool maxpool_214(
				.clk(clk),
				.rstn(rstn),
				.a0(A1484),
				.a1(A1494),
				.a2(A1584),
				.a3(A1594),
				.p(P2244)
);

maxpool maxpool_215(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A4),
				.a1(A14B4),
				.a2(A15A4),
				.a3(A15B4),
				.p(P2254)
);

maxpool maxpool_216(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C4),
				.a1(A14D4),
				.a2(A15C4),
				.a3(A15D4),
				.p(P2264)
);

maxpool maxpool_217(
				.clk(clk),
				.rstn(rstn),
				.a0(A1604),
				.a1(A1614),
				.a2(A1704),
				.a3(A1714),
				.p(P2304)
);

maxpool maxpool_218(
				.clk(clk),
				.rstn(rstn),
				.a0(A1624),
				.a1(A1634),
				.a2(A1724),
				.a3(A1734),
				.p(P2314)
);

maxpool maxpool_219(
				.clk(clk),
				.rstn(rstn),
				.a0(A1644),
				.a1(A1654),
				.a2(A1744),
				.a3(A1754),
				.p(P2324)
);

maxpool maxpool_220(
				.clk(clk),
				.rstn(rstn),
				.a0(A1664),
				.a1(A1674),
				.a2(A1764),
				.a3(A1774),
				.p(P2334)
);

maxpool maxpool_221(
				.clk(clk),
				.rstn(rstn),
				.a0(A1684),
				.a1(A1694),
				.a2(A1784),
				.a3(A1794),
				.p(P2344)
);

maxpool maxpool_222(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A4),
				.a1(A16B4),
				.a2(A17A4),
				.a3(A17B4),
				.p(P2354)
);

maxpool maxpool_223(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C4),
				.a1(A16D4),
				.a2(A17C4),
				.a3(A17D4),
				.p(P2364)
);

maxpool maxpool_224(
				.clk(clk),
				.rstn(rstn),
				.a0(A1804),
				.a1(A1814),
				.a2(A1904),
				.a3(A1914),
				.p(P2404)
);

maxpool maxpool_225(
				.clk(clk),
				.rstn(rstn),
				.a0(A1824),
				.a1(A1834),
				.a2(A1924),
				.a3(A1934),
				.p(P2414)
);

maxpool maxpool_226(
				.clk(clk),
				.rstn(rstn),
				.a0(A1844),
				.a1(A1854),
				.a2(A1944),
				.a3(A1954),
				.p(P2424)
);

maxpool maxpool_227(
				.clk(clk),
				.rstn(rstn),
				.a0(A1864),
				.a1(A1874),
				.a2(A1964),
				.a3(A1974),
				.p(P2434)
);

maxpool maxpool_228(
				.clk(clk),
				.rstn(rstn),
				.a0(A1884),
				.a1(A1894),
				.a2(A1984),
				.a3(A1994),
				.p(P2444)
);

maxpool maxpool_229(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A4),
				.a1(A18B4),
				.a2(A19A4),
				.a3(A19B4),
				.p(P2454)
);

maxpool maxpool_230(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C4),
				.a1(A18D4),
				.a2(A19C4),
				.a3(A19D4),
				.p(P2464)
);

maxpool maxpool_231(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A04),
				.a1(A1A14),
				.a2(A1B04),
				.a3(A1B14),
				.p(P2504)
);

maxpool maxpool_232(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A24),
				.a1(A1A34),
				.a2(A1B24),
				.a3(A1B34),
				.p(P2514)
);

maxpool maxpool_233(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A44),
				.a1(A1A54),
				.a2(A1B44),
				.a3(A1B54),
				.p(P2524)
);

maxpool maxpool_234(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A64),
				.a1(A1A74),
				.a2(A1B64),
				.a3(A1B74),
				.p(P2534)
);

maxpool maxpool_235(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A84),
				.a1(A1A94),
				.a2(A1B84),
				.a3(A1B94),
				.p(P2544)
);

maxpool maxpool_236(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA4),
				.a1(A1AB4),
				.a2(A1BA4),
				.a3(A1BB4),
				.p(P2554)
);

maxpool maxpool_237(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC4),
				.a1(A1AD4),
				.a2(A1BC4),
				.a3(A1BD4),
				.p(P2564)
);

maxpool maxpool_238(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C04),
				.a1(A1C14),
				.a2(A1D04),
				.a3(A1D14),
				.p(P2604)
);

maxpool maxpool_239(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C24),
				.a1(A1C34),
				.a2(A1D24),
				.a3(A1D34),
				.p(P2614)
);

maxpool maxpool_240(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C44),
				.a1(A1C54),
				.a2(A1D44),
				.a3(A1D54),
				.p(P2624)
);

maxpool maxpool_241(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C64),
				.a1(A1C74),
				.a2(A1D64),
				.a3(A1D74),
				.p(P2634)
);

maxpool maxpool_242(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C84),
				.a1(A1C94),
				.a2(A1D84),
				.a3(A1D94),
				.p(P2644)
);

maxpool maxpool_243(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA4),
				.a1(A1CB4),
				.a2(A1DA4),
				.a3(A1DB4),
				.p(P2654)
);

maxpool maxpool_244(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC4),
				.a1(A1CD4),
				.a2(A1DC4),
				.a3(A1DD4),
				.p(P2664)
);

maxpool maxpool_245(
				.clk(clk),
				.rstn(rstn),
				.a0(A1005),
				.a1(A1015),
				.a2(A1105),
				.a3(A1115),
				.p(P2005)
);

maxpool maxpool_246(
				.clk(clk),
				.rstn(rstn),
				.a0(A1025),
				.a1(A1035),
				.a2(A1125),
				.a3(A1135),
				.p(P2015)
);

maxpool maxpool_247(
				.clk(clk),
				.rstn(rstn),
				.a0(A1045),
				.a1(A1055),
				.a2(A1145),
				.a3(A1155),
				.p(P2025)
);

maxpool maxpool_248(
				.clk(clk),
				.rstn(rstn),
				.a0(A1065),
				.a1(A1075),
				.a2(A1165),
				.a3(A1175),
				.p(P2035)
);

maxpool maxpool_249(
				.clk(clk),
				.rstn(rstn),
				.a0(A1085),
				.a1(A1095),
				.a2(A1185),
				.a3(A1195),
				.p(P2045)
);

maxpool maxpool_250(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A5),
				.a1(A10B5),
				.a2(A11A5),
				.a3(A11B5),
				.p(P2055)
);

maxpool maxpool_251(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C5),
				.a1(A10D5),
				.a2(A11C5),
				.a3(A11D5),
				.p(P2065)
);

maxpool maxpool_252(
				.clk(clk),
				.rstn(rstn),
				.a0(A1205),
				.a1(A1215),
				.a2(A1305),
				.a3(A1315),
				.p(P2105)
);

maxpool maxpool_253(
				.clk(clk),
				.rstn(rstn),
				.a0(A1225),
				.a1(A1235),
				.a2(A1325),
				.a3(A1335),
				.p(P2115)
);

maxpool maxpool_254(
				.clk(clk),
				.rstn(rstn),
				.a0(A1245),
				.a1(A1255),
				.a2(A1345),
				.a3(A1355),
				.p(P2125)
);

maxpool maxpool_255(
				.clk(clk),
				.rstn(rstn),
				.a0(A1265),
				.a1(A1275),
				.a2(A1365),
				.a3(A1375),
				.p(P2135)
);

maxpool maxpool_256(
				.clk(clk),
				.rstn(rstn),
				.a0(A1285),
				.a1(A1295),
				.a2(A1385),
				.a3(A1395),
				.p(P2145)
);

maxpool maxpool_257(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A5),
				.a1(A12B5),
				.a2(A13A5),
				.a3(A13B5),
				.p(P2155)
);

maxpool maxpool_258(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C5),
				.a1(A12D5),
				.a2(A13C5),
				.a3(A13D5),
				.p(P2165)
);

maxpool maxpool_259(
				.clk(clk),
				.rstn(rstn),
				.a0(A1405),
				.a1(A1415),
				.a2(A1505),
				.a3(A1515),
				.p(P2205)
);

maxpool maxpool_260(
				.clk(clk),
				.rstn(rstn),
				.a0(A1425),
				.a1(A1435),
				.a2(A1525),
				.a3(A1535),
				.p(P2215)
);

maxpool maxpool_261(
				.clk(clk),
				.rstn(rstn),
				.a0(A1445),
				.a1(A1455),
				.a2(A1545),
				.a3(A1555),
				.p(P2225)
);

maxpool maxpool_262(
				.clk(clk),
				.rstn(rstn),
				.a0(A1465),
				.a1(A1475),
				.a2(A1565),
				.a3(A1575),
				.p(P2235)
);

maxpool maxpool_263(
				.clk(clk),
				.rstn(rstn),
				.a0(A1485),
				.a1(A1495),
				.a2(A1585),
				.a3(A1595),
				.p(P2245)
);

maxpool maxpool_264(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A5),
				.a1(A14B5),
				.a2(A15A5),
				.a3(A15B5),
				.p(P2255)
);

maxpool maxpool_265(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C5),
				.a1(A14D5),
				.a2(A15C5),
				.a3(A15D5),
				.p(P2265)
);

maxpool maxpool_266(
				.clk(clk),
				.rstn(rstn),
				.a0(A1605),
				.a1(A1615),
				.a2(A1705),
				.a3(A1715),
				.p(P2305)
);

maxpool maxpool_267(
				.clk(clk),
				.rstn(rstn),
				.a0(A1625),
				.a1(A1635),
				.a2(A1725),
				.a3(A1735),
				.p(P2315)
);

maxpool maxpool_268(
				.clk(clk),
				.rstn(rstn),
				.a0(A1645),
				.a1(A1655),
				.a2(A1745),
				.a3(A1755),
				.p(P2325)
);

maxpool maxpool_269(
				.clk(clk),
				.rstn(rstn),
				.a0(A1665),
				.a1(A1675),
				.a2(A1765),
				.a3(A1775),
				.p(P2335)
);

maxpool maxpool_270(
				.clk(clk),
				.rstn(rstn),
				.a0(A1685),
				.a1(A1695),
				.a2(A1785),
				.a3(A1795),
				.p(P2345)
);

maxpool maxpool_271(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A5),
				.a1(A16B5),
				.a2(A17A5),
				.a3(A17B5),
				.p(P2355)
);

maxpool maxpool_272(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C5),
				.a1(A16D5),
				.a2(A17C5),
				.a3(A17D5),
				.p(P2365)
);

maxpool maxpool_273(
				.clk(clk),
				.rstn(rstn),
				.a0(A1805),
				.a1(A1815),
				.a2(A1905),
				.a3(A1915),
				.p(P2405)
);

maxpool maxpool_274(
				.clk(clk),
				.rstn(rstn),
				.a0(A1825),
				.a1(A1835),
				.a2(A1925),
				.a3(A1935),
				.p(P2415)
);

maxpool maxpool_275(
				.clk(clk),
				.rstn(rstn),
				.a0(A1845),
				.a1(A1855),
				.a2(A1945),
				.a3(A1955),
				.p(P2425)
);

maxpool maxpool_276(
				.clk(clk),
				.rstn(rstn),
				.a0(A1865),
				.a1(A1875),
				.a2(A1965),
				.a3(A1975),
				.p(P2435)
);

maxpool maxpool_277(
				.clk(clk),
				.rstn(rstn),
				.a0(A1885),
				.a1(A1895),
				.a2(A1985),
				.a3(A1995),
				.p(P2445)
);

maxpool maxpool_278(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A5),
				.a1(A18B5),
				.a2(A19A5),
				.a3(A19B5),
				.p(P2455)
);

maxpool maxpool_279(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C5),
				.a1(A18D5),
				.a2(A19C5),
				.a3(A19D5),
				.p(P2465)
);

maxpool maxpool_280(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A05),
				.a1(A1A15),
				.a2(A1B05),
				.a3(A1B15),
				.p(P2505)
);

maxpool maxpool_281(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A25),
				.a1(A1A35),
				.a2(A1B25),
				.a3(A1B35),
				.p(P2515)
);

maxpool maxpool_282(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A45),
				.a1(A1A55),
				.a2(A1B45),
				.a3(A1B55),
				.p(P2525)
);

maxpool maxpool_283(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A65),
				.a1(A1A75),
				.a2(A1B65),
				.a3(A1B75),
				.p(P2535)
);

maxpool maxpool_284(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A85),
				.a1(A1A95),
				.a2(A1B85),
				.a3(A1B95),
				.p(P2545)
);

maxpool maxpool_285(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA5),
				.a1(A1AB5),
				.a2(A1BA5),
				.a3(A1BB5),
				.p(P2555)
);

maxpool maxpool_286(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC5),
				.a1(A1AD5),
				.a2(A1BC5),
				.a3(A1BD5),
				.p(P2565)
);

maxpool maxpool_287(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C05),
				.a1(A1C15),
				.a2(A1D05),
				.a3(A1D15),
				.p(P2605)
);

maxpool maxpool_288(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C25),
				.a1(A1C35),
				.a2(A1D25),
				.a3(A1D35),
				.p(P2615)
);

maxpool maxpool_289(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C45),
				.a1(A1C55),
				.a2(A1D45),
				.a3(A1D55),
				.p(P2625)
);

maxpool maxpool_290(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C65),
				.a1(A1C75),
				.a2(A1D65),
				.a3(A1D75),
				.p(P2635)
);

maxpool maxpool_291(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C85),
				.a1(A1C95),
				.a2(A1D85),
				.a3(A1D95),
				.p(P2645)
);

maxpool maxpool_292(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA5),
				.a1(A1CB5),
				.a2(A1DA5),
				.a3(A1DB5),
				.p(P2655)
);

maxpool maxpool_293(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC5),
				.a1(A1CD5),
				.a2(A1DC5),
				.a3(A1DD5),
				.p(P2665)
);

maxpool maxpool_294(
				.clk(clk),
				.rstn(rstn),
				.a0(A1006),
				.a1(A1016),
				.a2(A1106),
				.a3(A1116),
				.p(P2006)
);

maxpool maxpool_295(
				.clk(clk),
				.rstn(rstn),
				.a0(A1026),
				.a1(A1036),
				.a2(A1126),
				.a3(A1136),
				.p(P2016)
);

maxpool maxpool_296(
				.clk(clk),
				.rstn(rstn),
				.a0(A1046),
				.a1(A1056),
				.a2(A1146),
				.a3(A1156),
				.p(P2026)
);

maxpool maxpool_297(
				.clk(clk),
				.rstn(rstn),
				.a0(A1066),
				.a1(A1076),
				.a2(A1166),
				.a3(A1176),
				.p(P2036)
);

maxpool maxpool_298(
				.clk(clk),
				.rstn(rstn),
				.a0(A1086),
				.a1(A1096),
				.a2(A1186),
				.a3(A1196),
				.p(P2046)
);

maxpool maxpool_299(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A6),
				.a1(A10B6),
				.a2(A11A6),
				.a3(A11B6),
				.p(P2056)
);

maxpool maxpool_300(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C6),
				.a1(A10D6),
				.a2(A11C6),
				.a3(A11D6),
				.p(P2066)
);

maxpool maxpool_301(
				.clk(clk),
				.rstn(rstn),
				.a0(A1206),
				.a1(A1216),
				.a2(A1306),
				.a3(A1316),
				.p(P2106)
);

maxpool maxpool_302(
				.clk(clk),
				.rstn(rstn),
				.a0(A1226),
				.a1(A1236),
				.a2(A1326),
				.a3(A1336),
				.p(P2116)
);

maxpool maxpool_303(
				.clk(clk),
				.rstn(rstn),
				.a0(A1246),
				.a1(A1256),
				.a2(A1346),
				.a3(A1356),
				.p(P2126)
);

maxpool maxpool_304(
				.clk(clk),
				.rstn(rstn),
				.a0(A1266),
				.a1(A1276),
				.a2(A1366),
				.a3(A1376),
				.p(P2136)
);

maxpool maxpool_305(
				.clk(clk),
				.rstn(rstn),
				.a0(A1286),
				.a1(A1296),
				.a2(A1386),
				.a3(A1396),
				.p(P2146)
);

maxpool maxpool_306(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A6),
				.a1(A12B6),
				.a2(A13A6),
				.a3(A13B6),
				.p(P2156)
);

maxpool maxpool_307(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C6),
				.a1(A12D6),
				.a2(A13C6),
				.a3(A13D6),
				.p(P2166)
);

maxpool maxpool_308(
				.clk(clk),
				.rstn(rstn),
				.a0(A1406),
				.a1(A1416),
				.a2(A1506),
				.a3(A1516),
				.p(P2206)
);

maxpool maxpool_309(
				.clk(clk),
				.rstn(rstn),
				.a0(A1426),
				.a1(A1436),
				.a2(A1526),
				.a3(A1536),
				.p(P2216)
);

maxpool maxpool_310(
				.clk(clk),
				.rstn(rstn),
				.a0(A1446),
				.a1(A1456),
				.a2(A1546),
				.a3(A1556),
				.p(P2226)
);

maxpool maxpool_311(
				.clk(clk),
				.rstn(rstn),
				.a0(A1466),
				.a1(A1476),
				.a2(A1566),
				.a3(A1576),
				.p(P2236)
);

maxpool maxpool_312(
				.clk(clk),
				.rstn(rstn),
				.a0(A1486),
				.a1(A1496),
				.a2(A1586),
				.a3(A1596),
				.p(P2246)
);

maxpool maxpool_313(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A6),
				.a1(A14B6),
				.a2(A15A6),
				.a3(A15B6),
				.p(P2256)
);

maxpool maxpool_314(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C6),
				.a1(A14D6),
				.a2(A15C6),
				.a3(A15D6),
				.p(P2266)
);

maxpool maxpool_315(
				.clk(clk),
				.rstn(rstn),
				.a0(A1606),
				.a1(A1616),
				.a2(A1706),
				.a3(A1716),
				.p(P2306)
);

maxpool maxpool_316(
				.clk(clk),
				.rstn(rstn),
				.a0(A1626),
				.a1(A1636),
				.a2(A1726),
				.a3(A1736),
				.p(P2316)
);

maxpool maxpool_317(
				.clk(clk),
				.rstn(rstn),
				.a0(A1646),
				.a1(A1656),
				.a2(A1746),
				.a3(A1756),
				.p(P2326)
);

maxpool maxpool_318(
				.clk(clk),
				.rstn(rstn),
				.a0(A1666),
				.a1(A1676),
				.a2(A1766),
				.a3(A1776),
				.p(P2336)
);

maxpool maxpool_319(
				.clk(clk),
				.rstn(rstn),
				.a0(A1686),
				.a1(A1696),
				.a2(A1786),
				.a3(A1796),
				.p(P2346)
);

maxpool maxpool_320(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A6),
				.a1(A16B6),
				.a2(A17A6),
				.a3(A17B6),
				.p(P2356)
);

maxpool maxpool_321(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C6),
				.a1(A16D6),
				.a2(A17C6),
				.a3(A17D6),
				.p(P2366)
);

maxpool maxpool_322(
				.clk(clk),
				.rstn(rstn),
				.a0(A1806),
				.a1(A1816),
				.a2(A1906),
				.a3(A1916),
				.p(P2406)
);

maxpool maxpool_323(
				.clk(clk),
				.rstn(rstn),
				.a0(A1826),
				.a1(A1836),
				.a2(A1926),
				.a3(A1936),
				.p(P2416)
);

maxpool maxpool_324(
				.clk(clk),
				.rstn(rstn),
				.a0(A1846),
				.a1(A1856),
				.a2(A1946),
				.a3(A1956),
				.p(P2426)
);

maxpool maxpool_325(
				.clk(clk),
				.rstn(rstn),
				.a0(A1866),
				.a1(A1876),
				.a2(A1966),
				.a3(A1976),
				.p(P2436)
);

maxpool maxpool_326(
				.clk(clk),
				.rstn(rstn),
				.a0(A1886),
				.a1(A1896),
				.a2(A1986),
				.a3(A1996),
				.p(P2446)
);

maxpool maxpool_327(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A6),
				.a1(A18B6),
				.a2(A19A6),
				.a3(A19B6),
				.p(P2456)
);

maxpool maxpool_328(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C6),
				.a1(A18D6),
				.a2(A19C6),
				.a3(A19D6),
				.p(P2466)
);

maxpool maxpool_329(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A06),
				.a1(A1A16),
				.a2(A1B06),
				.a3(A1B16),
				.p(P2506)
);

maxpool maxpool_330(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A26),
				.a1(A1A36),
				.a2(A1B26),
				.a3(A1B36),
				.p(P2516)
);

maxpool maxpool_331(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A46),
				.a1(A1A56),
				.a2(A1B46),
				.a3(A1B56),
				.p(P2526)
);

maxpool maxpool_332(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A66),
				.a1(A1A76),
				.a2(A1B66),
				.a3(A1B76),
				.p(P2536)
);

maxpool maxpool_333(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A86),
				.a1(A1A96),
				.a2(A1B86),
				.a3(A1B96),
				.p(P2546)
);

maxpool maxpool_334(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA6),
				.a1(A1AB6),
				.a2(A1BA6),
				.a3(A1BB6),
				.p(P2556)
);

maxpool maxpool_335(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC6),
				.a1(A1AD6),
				.a2(A1BC6),
				.a3(A1BD6),
				.p(P2566)
);

maxpool maxpool_336(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C06),
				.a1(A1C16),
				.a2(A1D06),
				.a3(A1D16),
				.p(P2606)
);

maxpool maxpool_337(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C26),
				.a1(A1C36),
				.a2(A1D26),
				.a3(A1D36),
				.p(P2616)
);

maxpool maxpool_338(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C46),
				.a1(A1C56),
				.a2(A1D46),
				.a3(A1D56),
				.p(P2626)
);

maxpool maxpool_339(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C66),
				.a1(A1C76),
				.a2(A1D66),
				.a3(A1D76),
				.p(P2636)
);

maxpool maxpool_340(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C86),
				.a1(A1C96),
				.a2(A1D86),
				.a3(A1D96),
				.p(P2646)
);

maxpool maxpool_341(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA6),
				.a1(A1CB6),
				.a2(A1DA6),
				.a3(A1DB6),
				.p(P2656)
);

maxpool maxpool_342(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC6),
				.a1(A1CD6),
				.a2(A1DC6),
				.a3(A1DD6),
				.p(P2666)
);

maxpool maxpool_343(
				.clk(clk),
				.rstn(rstn),
				.a0(A1007),
				.a1(A1017),
				.a2(A1107),
				.a3(A1117),
				.p(P2007)
);

maxpool maxpool_344(
				.clk(clk),
				.rstn(rstn),
				.a0(A1027),
				.a1(A1037),
				.a2(A1127),
				.a3(A1137),
				.p(P2017)
);

maxpool maxpool_345(
				.clk(clk),
				.rstn(rstn),
				.a0(A1047),
				.a1(A1057),
				.a2(A1147),
				.a3(A1157),
				.p(P2027)
);

maxpool maxpool_346(
				.clk(clk),
				.rstn(rstn),
				.a0(A1067),
				.a1(A1077),
				.a2(A1167),
				.a3(A1177),
				.p(P2037)
);

maxpool maxpool_347(
				.clk(clk),
				.rstn(rstn),
				.a0(A1087),
				.a1(A1097),
				.a2(A1187),
				.a3(A1197),
				.p(P2047)
);

maxpool maxpool_348(
				.clk(clk),
				.rstn(rstn),
				.a0(A10A7),
				.a1(A10B7),
				.a2(A11A7),
				.a3(A11B7),
				.p(P2057)
);

maxpool maxpool_349(
				.clk(clk),
				.rstn(rstn),
				.a0(A10C7),
				.a1(A10D7),
				.a2(A11C7),
				.a3(A11D7),
				.p(P2067)
);

maxpool maxpool_350(
				.clk(clk),
				.rstn(rstn),
				.a0(A1207),
				.a1(A1217),
				.a2(A1307),
				.a3(A1317),
				.p(P2107)
);

maxpool maxpool_351(
				.clk(clk),
				.rstn(rstn),
				.a0(A1227),
				.a1(A1237),
				.a2(A1327),
				.a3(A1337),
				.p(P2117)
);

maxpool maxpool_352(
				.clk(clk),
				.rstn(rstn),
				.a0(A1247),
				.a1(A1257),
				.a2(A1347),
				.a3(A1357),
				.p(P2127)
);

maxpool maxpool_353(
				.clk(clk),
				.rstn(rstn),
				.a0(A1267),
				.a1(A1277),
				.a2(A1367),
				.a3(A1377),
				.p(P2137)
);

maxpool maxpool_354(
				.clk(clk),
				.rstn(rstn),
				.a0(A1287),
				.a1(A1297),
				.a2(A1387),
				.a3(A1397),
				.p(P2147)
);

maxpool maxpool_355(
				.clk(clk),
				.rstn(rstn),
				.a0(A12A7),
				.a1(A12B7),
				.a2(A13A7),
				.a3(A13B7),
				.p(P2157)
);

maxpool maxpool_356(
				.clk(clk),
				.rstn(rstn),
				.a0(A12C7),
				.a1(A12D7),
				.a2(A13C7),
				.a3(A13D7),
				.p(P2167)
);

maxpool maxpool_357(
				.clk(clk),
				.rstn(rstn),
				.a0(A1407),
				.a1(A1417),
				.a2(A1507),
				.a3(A1517),
				.p(P2207)
);

maxpool maxpool_358(
				.clk(clk),
				.rstn(rstn),
				.a0(A1427),
				.a1(A1437),
				.a2(A1527),
				.a3(A1537),
				.p(P2217)
);

maxpool maxpool_359(
				.clk(clk),
				.rstn(rstn),
				.a0(A1447),
				.a1(A1457),
				.a2(A1547),
				.a3(A1557),
				.p(P2227)
);

maxpool maxpool_360(
				.clk(clk),
				.rstn(rstn),
				.a0(A1467),
				.a1(A1477),
				.a2(A1567),
				.a3(A1577),
				.p(P2237)
);

maxpool maxpool_361(
				.clk(clk),
				.rstn(rstn),
				.a0(A1487),
				.a1(A1497),
				.a2(A1587),
				.a3(A1597),
				.p(P2247)
);

maxpool maxpool_362(
				.clk(clk),
				.rstn(rstn),
				.a0(A14A7),
				.a1(A14B7),
				.a2(A15A7),
				.a3(A15B7),
				.p(P2257)
);

maxpool maxpool_363(
				.clk(clk),
				.rstn(rstn),
				.a0(A14C7),
				.a1(A14D7),
				.a2(A15C7),
				.a3(A15D7),
				.p(P2267)
);

maxpool maxpool_364(
				.clk(clk),
				.rstn(rstn),
				.a0(A1607),
				.a1(A1617),
				.a2(A1707),
				.a3(A1717),
				.p(P2307)
);

maxpool maxpool_365(
				.clk(clk),
				.rstn(rstn),
				.a0(A1627),
				.a1(A1637),
				.a2(A1727),
				.a3(A1737),
				.p(P2317)
);

maxpool maxpool_366(
				.clk(clk),
				.rstn(rstn),
				.a0(A1647),
				.a1(A1657),
				.a2(A1747),
				.a3(A1757),
				.p(P2327)
);

maxpool maxpool_367(
				.clk(clk),
				.rstn(rstn),
				.a0(A1667),
				.a1(A1677),
				.a2(A1767),
				.a3(A1777),
				.p(P2337)
);

maxpool maxpool_368(
				.clk(clk),
				.rstn(rstn),
				.a0(A1687),
				.a1(A1697),
				.a2(A1787),
				.a3(A1797),
				.p(P2347)
);

maxpool maxpool_369(
				.clk(clk),
				.rstn(rstn),
				.a0(A16A7),
				.a1(A16B7),
				.a2(A17A7),
				.a3(A17B7),
				.p(P2357)
);

maxpool maxpool_370(
				.clk(clk),
				.rstn(rstn),
				.a0(A16C7),
				.a1(A16D7),
				.a2(A17C7),
				.a3(A17D7),
				.p(P2367)
);

maxpool maxpool_371(
				.clk(clk),
				.rstn(rstn),
				.a0(A1807),
				.a1(A1817),
				.a2(A1907),
				.a3(A1917),
				.p(P2407)
);

maxpool maxpool_372(
				.clk(clk),
				.rstn(rstn),
				.a0(A1827),
				.a1(A1837),
				.a2(A1927),
				.a3(A1937),
				.p(P2417)
);

maxpool maxpool_373(
				.clk(clk),
				.rstn(rstn),
				.a0(A1847),
				.a1(A1857),
				.a2(A1947),
				.a3(A1957),
				.p(P2427)
);

maxpool maxpool_374(
				.clk(clk),
				.rstn(rstn),
				.a0(A1867),
				.a1(A1877),
				.a2(A1967),
				.a3(A1977),
				.p(P2437)
);

maxpool maxpool_375(
				.clk(clk),
				.rstn(rstn),
				.a0(A1887),
				.a1(A1897),
				.a2(A1987),
				.a3(A1997),
				.p(P2447)
);

maxpool maxpool_376(
				.clk(clk),
				.rstn(rstn),
				.a0(A18A7),
				.a1(A18B7),
				.a2(A19A7),
				.a3(A19B7),
				.p(P2457)
);

maxpool maxpool_377(
				.clk(clk),
				.rstn(rstn),
				.a0(A18C7),
				.a1(A18D7),
				.a2(A19C7),
				.a3(A19D7),
				.p(P2467)
);

maxpool maxpool_378(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A07),
				.a1(A1A17),
				.a2(A1B07),
				.a3(A1B17),
				.p(P2507)
);

maxpool maxpool_379(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A27),
				.a1(A1A37),
				.a2(A1B27),
				.a3(A1B37),
				.p(P2517)
);

maxpool maxpool_380(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A47),
				.a1(A1A57),
				.a2(A1B47),
				.a3(A1B57),
				.p(P2527)
);

maxpool maxpool_381(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A67),
				.a1(A1A77),
				.a2(A1B67),
				.a3(A1B77),
				.p(P2537)
);

maxpool maxpool_382(
				.clk(clk),
				.rstn(rstn),
				.a0(A1A87),
				.a1(A1A97),
				.a2(A1B87),
				.a3(A1B97),
				.p(P2547)
);

maxpool maxpool_383(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AA7),
				.a1(A1AB7),
				.a2(A1BA7),
				.a3(A1BB7),
				.p(P2557)
);

maxpool maxpool_384(
				.clk(clk),
				.rstn(rstn),
				.a0(A1AC7),
				.a1(A1AD7),
				.a2(A1BC7),
				.a3(A1BD7),
				.p(P2567)
);

maxpool maxpool_385(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C07),
				.a1(A1C17),
				.a2(A1D07),
				.a3(A1D17),
				.p(P2607)
);

maxpool maxpool_386(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C27),
				.a1(A1C37),
				.a2(A1D27),
				.a3(A1D37),
				.p(P2617)
);

maxpool maxpool_387(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C47),
				.a1(A1C57),
				.a2(A1D47),
				.a3(A1D57),
				.p(P2627)
);

maxpool maxpool_388(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C67),
				.a1(A1C77),
				.a2(A1D67),
				.a3(A1D77),
				.p(P2637)
);

maxpool maxpool_389(
				.clk(clk),
				.rstn(rstn),
				.a0(A1C87),
				.a1(A1C97),
				.a2(A1D87),
				.a3(A1D97),
				.p(P2647)
);

maxpool maxpool_390(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CA7),
				.a1(A1CB7),
				.a2(A1DA7),
				.a3(A1DB7),
				.p(P2657)
);

maxpool maxpool_391(
				.clk(clk),
				.rstn(rstn),
				.a0(A1CC7),
				.a1(A1CD7),
				.a2(A1DC7),
				.a3(A1DD7),
				.p(P2667)
);

endmodule