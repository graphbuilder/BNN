module test_layer_all(
clk, 
rstn
);
input clk;
input rstn;

(*DONT_TOUCH="true"*) wire P2000;
(*DONT_TOUCH="true"*) wire P2010;
(*DONT_TOUCH="true"*) wire P2020;
(*DONT_TOUCH="true"*) wire P2030;
(*DONT_TOUCH="true"*) wire P2040;
(*DONT_TOUCH="true"*) wire P2050;
(*DONT_TOUCH="true"*) wire P2060;
(*DONT_TOUCH="true"*) wire P2100;
(*DONT_TOUCH="true"*) wire P2110;
(*DONT_TOUCH="true"*) wire P2120;
(*DONT_TOUCH="true"*) wire P2130;
(*DONT_TOUCH="true"*) wire P2140;
(*DONT_TOUCH="true"*) wire P2150;
(*DONT_TOUCH="true"*) wire P2160;
(*DONT_TOUCH="true"*) wire P2200;
(*DONT_TOUCH="true"*) wire P2210;
(*DONT_TOUCH="true"*) wire P2220;
(*DONT_TOUCH="true"*) wire P2230;
(*DONT_TOUCH="true"*) wire P2240;
(*DONT_TOUCH="true"*) wire P2250;
(*DONT_TOUCH="true"*) wire P2260;
(*DONT_TOUCH="true"*) wire P2300;
(*DONT_TOUCH="true"*) wire P2310;
(*DONT_TOUCH="true"*) wire P2320;
(*DONT_TOUCH="true"*) wire P2330;
(*DONT_TOUCH="true"*) wire P2340;
(*DONT_TOUCH="true"*) wire P2350;
(*DONT_TOUCH="true"*) wire P2360;
(*DONT_TOUCH="true"*) wire P2400;
(*DONT_TOUCH="true"*) wire P2410;
(*DONT_TOUCH="true"*) wire P2420;
(*DONT_TOUCH="true"*) wire P2430;
(*DONT_TOUCH="true"*) wire P2440;
(*DONT_TOUCH="true"*) wire P2450;
(*DONT_TOUCH="true"*) wire P2460;
(*DONT_TOUCH="true"*) wire P2500;
(*DONT_TOUCH="true"*) wire P2510;
(*DONT_TOUCH="true"*) wire P2520;
(*DONT_TOUCH="true"*) wire P2530;
(*DONT_TOUCH="true"*) wire P2540;
(*DONT_TOUCH="true"*) wire P2550;
(*DONT_TOUCH="true"*) wire P2560;
(*DONT_TOUCH="true"*) wire P2600;
(*DONT_TOUCH="true"*) wire P2610;
(*DONT_TOUCH="true"*) wire P2620;
(*DONT_TOUCH="true"*) wire P2630;
(*DONT_TOUCH="true"*) wire P2640;
(*DONT_TOUCH="true"*) wire P2650;
(*DONT_TOUCH="true"*) wire P2660;
(*DONT_TOUCH="true"*) wire P2001;
(*DONT_TOUCH="true"*) wire P2011;
(*DONT_TOUCH="true"*) wire P2021;
(*DONT_TOUCH="true"*) wire P2031;
(*DONT_TOUCH="true"*) wire P2041;
(*DONT_TOUCH="true"*) wire P2051;
(*DONT_TOUCH="true"*) wire P2061;
(*DONT_TOUCH="true"*) wire P2101;
(*DONT_TOUCH="true"*) wire P2111;
(*DONT_TOUCH="true"*) wire P2121;
(*DONT_TOUCH="true"*) wire P2131;
(*DONT_TOUCH="true"*) wire P2141;
(*DONT_TOUCH="true"*) wire P2151;
(*DONT_TOUCH="true"*) wire P2161;
(*DONT_TOUCH="true"*) wire P2201;
(*DONT_TOUCH="true"*) wire P2211;
(*DONT_TOUCH="true"*) wire P2221;
(*DONT_TOUCH="true"*) wire P2231;
(*DONT_TOUCH="true"*) wire P2241;
(*DONT_TOUCH="true"*) wire P2251;
(*DONT_TOUCH="true"*) wire P2261;
(*DONT_TOUCH="true"*) wire P2301;
(*DONT_TOUCH="true"*) wire P2311;
(*DONT_TOUCH="true"*) wire P2321;
(*DONT_TOUCH="true"*) wire P2331;
(*DONT_TOUCH="true"*) wire P2341;
(*DONT_TOUCH="true"*) wire P2351;
(*DONT_TOUCH="true"*) wire P2361;
(*DONT_TOUCH="true"*) wire P2401;
(*DONT_TOUCH="true"*) wire P2411;
(*DONT_TOUCH="true"*) wire P2421;
(*DONT_TOUCH="true"*) wire P2431;
(*DONT_TOUCH="true"*) wire P2441;
(*DONT_TOUCH="true"*) wire P2451;
(*DONT_TOUCH="true"*) wire P2461;
(*DONT_TOUCH="true"*) wire P2501;
(*DONT_TOUCH="true"*) wire P2511;
(*DONT_TOUCH="true"*) wire P2521;
(*DONT_TOUCH="true"*) wire P2531;
(*DONT_TOUCH="true"*) wire P2541;
(*DONT_TOUCH="true"*) wire P2551;
(*DONT_TOUCH="true"*) wire P2561;
(*DONT_TOUCH="true"*) wire P2601;
(*DONT_TOUCH="true"*) wire P2611;
(*DONT_TOUCH="true"*) wire P2621;
(*DONT_TOUCH="true"*) wire P2631;
(*DONT_TOUCH="true"*) wire P2641;
(*DONT_TOUCH="true"*) wire P2651;
(*DONT_TOUCH="true"*) wire P2661;
(*DONT_TOUCH="true"*) wire P2002;
(*DONT_TOUCH="true"*) wire P2012;
(*DONT_TOUCH="true"*) wire P2022;
(*DONT_TOUCH="true"*) wire P2032;
(*DONT_TOUCH="true"*) wire P2042;
(*DONT_TOUCH="true"*) wire P2052;
(*DONT_TOUCH="true"*) wire P2062;
(*DONT_TOUCH="true"*) wire P2102;
(*DONT_TOUCH="true"*) wire P2112;
(*DONT_TOUCH="true"*) wire P2122;
(*DONT_TOUCH="true"*) wire P2132;
(*DONT_TOUCH="true"*) wire P2142;
(*DONT_TOUCH="true"*) wire P2152;
(*DONT_TOUCH="true"*) wire P2162;
(*DONT_TOUCH="true"*) wire P2202;
(*DONT_TOUCH="true"*) wire P2212;
(*DONT_TOUCH="true"*) wire P2222;
(*DONT_TOUCH="true"*) wire P2232;
(*DONT_TOUCH="true"*) wire P2242;
(*DONT_TOUCH="true"*) wire P2252;
(*DONT_TOUCH="true"*) wire P2262;
(*DONT_TOUCH="true"*) wire P2302;
(*DONT_TOUCH="true"*) wire P2312;
(*DONT_TOUCH="true"*) wire P2322;
(*DONT_TOUCH="true"*) wire P2332;
(*DONT_TOUCH="true"*) wire P2342;
(*DONT_TOUCH="true"*) wire P2352;
(*DONT_TOUCH="true"*) wire P2362;
(*DONT_TOUCH="true"*) wire P2402;
(*DONT_TOUCH="true"*) wire P2412;
(*DONT_TOUCH="true"*) wire P2422;
(*DONT_TOUCH="true"*) wire P2432;
(*DONT_TOUCH="true"*) wire P2442;
(*DONT_TOUCH="true"*) wire P2452;
(*DONT_TOUCH="true"*) wire P2462;
(*DONT_TOUCH="true"*) wire P2502;
(*DONT_TOUCH="true"*) wire P2512;
(*DONT_TOUCH="true"*) wire P2522;
(*DONT_TOUCH="true"*) wire P2532;
(*DONT_TOUCH="true"*) wire P2542;
(*DONT_TOUCH="true"*) wire P2552;
(*DONT_TOUCH="true"*) wire P2562;
(*DONT_TOUCH="true"*) wire P2602;
(*DONT_TOUCH="true"*) wire P2612;
(*DONT_TOUCH="true"*) wire P2622;
(*DONT_TOUCH="true"*) wire P2632;
(*DONT_TOUCH="true"*) wire P2642;
(*DONT_TOUCH="true"*) wire P2652;
(*DONT_TOUCH="true"*) wire P2662;
(*DONT_TOUCH="true"*) wire P2003;
(*DONT_TOUCH="true"*) wire P2013;
(*DONT_TOUCH="true"*) wire P2023;
(*DONT_TOUCH="true"*) wire P2033;
(*DONT_TOUCH="true"*) wire P2043;
(*DONT_TOUCH="true"*) wire P2053;
(*DONT_TOUCH="true"*) wire P2063;
(*DONT_TOUCH="true"*) wire P2103;
(*DONT_TOUCH="true"*) wire P2113;
(*DONT_TOUCH="true"*) wire P2123;
(*DONT_TOUCH="true"*) wire P2133;
(*DONT_TOUCH="true"*) wire P2143;
(*DONT_TOUCH="true"*) wire P2153;
(*DONT_TOUCH="true"*) wire P2163;
(*DONT_TOUCH="true"*) wire P2203;
(*DONT_TOUCH="true"*) wire P2213;
(*DONT_TOUCH="true"*) wire P2223;
(*DONT_TOUCH="true"*) wire P2233;
(*DONT_TOUCH="true"*) wire P2243;
(*DONT_TOUCH="true"*) wire P2253;
(*DONT_TOUCH="true"*) wire P2263;
(*DONT_TOUCH="true"*) wire P2303;
(*DONT_TOUCH="true"*) wire P2313;
(*DONT_TOUCH="true"*) wire P2323;
(*DONT_TOUCH="true"*) wire P2333;
(*DONT_TOUCH="true"*) wire P2343;
(*DONT_TOUCH="true"*) wire P2353;
(*DONT_TOUCH="true"*) wire P2363;
(*DONT_TOUCH="true"*) wire P2403;
(*DONT_TOUCH="true"*) wire P2413;
(*DONT_TOUCH="true"*) wire P2423;
(*DONT_TOUCH="true"*) wire P2433;
(*DONT_TOUCH="true"*) wire P2443;
(*DONT_TOUCH="true"*) wire P2453;
(*DONT_TOUCH="true"*) wire P2463;
(*DONT_TOUCH="true"*) wire P2503;
(*DONT_TOUCH="true"*) wire P2513;
(*DONT_TOUCH="true"*) wire P2523;
(*DONT_TOUCH="true"*) wire P2533;
(*DONT_TOUCH="true"*) wire P2543;
(*DONT_TOUCH="true"*) wire P2553;
(*DONT_TOUCH="true"*) wire P2563;
(*DONT_TOUCH="true"*) wire P2603;
(*DONT_TOUCH="true"*) wire P2613;
(*DONT_TOUCH="true"*) wire P2623;
(*DONT_TOUCH="true"*) wire P2633;
(*DONT_TOUCH="true"*) wire P2643;
(*DONT_TOUCH="true"*) wire P2653;
(*DONT_TOUCH="true"*) wire P2663;
(*DONT_TOUCH="true"*) wire P2004;
(*DONT_TOUCH="true"*) wire P2014;
(*DONT_TOUCH="true"*) wire P2024;
(*DONT_TOUCH="true"*) wire P2034;
(*DONT_TOUCH="true"*) wire P2044;
(*DONT_TOUCH="true"*) wire P2054;
(*DONT_TOUCH="true"*) wire P2064;
(*DONT_TOUCH="true"*) wire P2104;
(*DONT_TOUCH="true"*) wire P2114;
(*DONT_TOUCH="true"*) wire P2124;
(*DONT_TOUCH="true"*) wire P2134;
(*DONT_TOUCH="true"*) wire P2144;
(*DONT_TOUCH="true"*) wire P2154;
(*DONT_TOUCH="true"*) wire P2164;
(*DONT_TOUCH="true"*) wire P2204;
(*DONT_TOUCH="true"*) wire P2214;
(*DONT_TOUCH="true"*) wire P2224;
(*DONT_TOUCH="true"*) wire P2234;
(*DONT_TOUCH="true"*) wire P2244;
(*DONT_TOUCH="true"*) wire P2254;
(*DONT_TOUCH="true"*) wire P2264;
(*DONT_TOUCH="true"*) wire P2304;
(*DONT_TOUCH="true"*) wire P2314;
(*DONT_TOUCH="true"*) wire P2324;
(*DONT_TOUCH="true"*) wire P2334;
(*DONT_TOUCH="true"*) wire P2344;
(*DONT_TOUCH="true"*) wire P2354;
(*DONT_TOUCH="true"*) wire P2364;
(*DONT_TOUCH="true"*) wire P2404;
(*DONT_TOUCH="true"*) wire P2414;
(*DONT_TOUCH="true"*) wire P2424;
(*DONT_TOUCH="true"*) wire P2434;
(*DONT_TOUCH="true"*) wire P2444;
(*DONT_TOUCH="true"*) wire P2454;
(*DONT_TOUCH="true"*) wire P2464;
(*DONT_TOUCH="true"*) wire P2504;
(*DONT_TOUCH="true"*) wire P2514;
(*DONT_TOUCH="true"*) wire P2524;
(*DONT_TOUCH="true"*) wire P2534;
(*DONT_TOUCH="true"*) wire P2544;
(*DONT_TOUCH="true"*) wire P2554;
(*DONT_TOUCH="true"*) wire P2564;
(*DONT_TOUCH="true"*) wire P2604;
(*DONT_TOUCH="true"*) wire P2614;
(*DONT_TOUCH="true"*) wire P2624;
(*DONT_TOUCH="true"*) wire P2634;
(*DONT_TOUCH="true"*) wire P2644;
(*DONT_TOUCH="true"*) wire P2654;
(*DONT_TOUCH="true"*) wire P2664;
(*DONT_TOUCH="true"*) wire P2005;
(*DONT_TOUCH="true"*) wire P2015;
(*DONT_TOUCH="true"*) wire P2025;
(*DONT_TOUCH="true"*) wire P2035;
(*DONT_TOUCH="true"*) wire P2045;
(*DONT_TOUCH="true"*) wire P2055;
(*DONT_TOUCH="true"*) wire P2065;
(*DONT_TOUCH="true"*) wire P2105;
(*DONT_TOUCH="true"*) wire P2115;
(*DONT_TOUCH="true"*) wire P2125;
(*DONT_TOUCH="true"*) wire P2135;
(*DONT_TOUCH="true"*) wire P2145;
(*DONT_TOUCH="true"*) wire P2155;
(*DONT_TOUCH="true"*) wire P2165;
(*DONT_TOUCH="true"*) wire P2205;
(*DONT_TOUCH="true"*) wire P2215;
(*DONT_TOUCH="true"*) wire P2225;
(*DONT_TOUCH="true"*) wire P2235;
(*DONT_TOUCH="true"*) wire P2245;
(*DONT_TOUCH="true"*) wire P2255;
(*DONT_TOUCH="true"*) wire P2265;
(*DONT_TOUCH="true"*) wire P2305;
(*DONT_TOUCH="true"*) wire P2315;
(*DONT_TOUCH="true"*) wire P2325;
(*DONT_TOUCH="true"*) wire P2335;
(*DONT_TOUCH="true"*) wire P2345;
(*DONT_TOUCH="true"*) wire P2355;
(*DONT_TOUCH="true"*) wire P2365;
(*DONT_TOUCH="true"*) wire P2405;
(*DONT_TOUCH="true"*) wire P2415;
(*DONT_TOUCH="true"*) wire P2425;
(*DONT_TOUCH="true"*) wire P2435;
(*DONT_TOUCH="true"*) wire P2445;
(*DONT_TOUCH="true"*) wire P2455;
(*DONT_TOUCH="true"*) wire P2465;
(*DONT_TOUCH="true"*) wire P2505;
(*DONT_TOUCH="true"*) wire P2515;
(*DONT_TOUCH="true"*) wire P2525;
(*DONT_TOUCH="true"*) wire P2535;
(*DONT_TOUCH="true"*) wire P2545;
(*DONT_TOUCH="true"*) wire P2555;
(*DONT_TOUCH="true"*) wire P2565;
(*DONT_TOUCH="true"*) wire P2605;
(*DONT_TOUCH="true"*) wire P2615;
(*DONT_TOUCH="true"*) wire P2625;
(*DONT_TOUCH="true"*) wire P2635;
(*DONT_TOUCH="true"*) wire P2645;
(*DONT_TOUCH="true"*) wire P2655;
(*DONT_TOUCH="true"*) wire P2665;
(*DONT_TOUCH="true"*) wire P2006;
(*DONT_TOUCH="true"*) wire P2016;
(*DONT_TOUCH="true"*) wire P2026;
(*DONT_TOUCH="true"*) wire P2036;
(*DONT_TOUCH="true"*) wire P2046;
(*DONT_TOUCH="true"*) wire P2056;
(*DONT_TOUCH="true"*) wire P2066;
(*DONT_TOUCH="true"*) wire P2106;
(*DONT_TOUCH="true"*) wire P2116;
(*DONT_TOUCH="true"*) wire P2126;
(*DONT_TOUCH="true"*) wire P2136;
(*DONT_TOUCH="true"*) wire P2146;
(*DONT_TOUCH="true"*) wire P2156;
(*DONT_TOUCH="true"*) wire P2166;
(*DONT_TOUCH="true"*) wire P2206;
(*DONT_TOUCH="true"*) wire P2216;
(*DONT_TOUCH="true"*) wire P2226;
(*DONT_TOUCH="true"*) wire P2236;
(*DONT_TOUCH="true"*) wire P2246;
(*DONT_TOUCH="true"*) wire P2256;
(*DONT_TOUCH="true"*) wire P2266;
(*DONT_TOUCH="true"*) wire P2306;
(*DONT_TOUCH="true"*) wire P2316;
(*DONT_TOUCH="true"*) wire P2326;
(*DONT_TOUCH="true"*) wire P2336;
(*DONT_TOUCH="true"*) wire P2346;
(*DONT_TOUCH="true"*) wire P2356;
(*DONT_TOUCH="true"*) wire P2366;
(*DONT_TOUCH="true"*) wire P2406;
(*DONT_TOUCH="true"*) wire P2416;
(*DONT_TOUCH="true"*) wire P2426;
(*DONT_TOUCH="true"*) wire P2436;
(*DONT_TOUCH="true"*) wire P2446;
(*DONT_TOUCH="true"*) wire P2456;
(*DONT_TOUCH="true"*) wire P2466;
(*DONT_TOUCH="true"*) wire P2506;
(*DONT_TOUCH="true"*) wire P2516;
(*DONT_TOUCH="true"*) wire P2526;
(*DONT_TOUCH="true"*) wire P2536;
(*DONT_TOUCH="true"*) wire P2546;
(*DONT_TOUCH="true"*) wire P2556;
(*DONT_TOUCH="true"*) wire P2566;
(*DONT_TOUCH="true"*) wire P2606;
(*DONT_TOUCH="true"*) wire P2616;
(*DONT_TOUCH="true"*) wire P2626;
(*DONT_TOUCH="true"*) wire P2636;
(*DONT_TOUCH="true"*) wire P2646;
(*DONT_TOUCH="true"*) wire P2656;
(*DONT_TOUCH="true"*) wire P2666;
(*DONT_TOUCH="true"*) wire P2007;
(*DONT_TOUCH="true"*) wire P2017;
(*DONT_TOUCH="true"*) wire P2027;
(*DONT_TOUCH="true"*) wire P2037;
(*DONT_TOUCH="true"*) wire P2047;
(*DONT_TOUCH="true"*) wire P2057;
(*DONT_TOUCH="true"*) wire P2067;
(*DONT_TOUCH="true"*) wire P2107;
(*DONT_TOUCH="true"*) wire P2117;
(*DONT_TOUCH="true"*) wire P2127;
(*DONT_TOUCH="true"*) wire P2137;
(*DONT_TOUCH="true"*) wire P2147;
(*DONT_TOUCH="true"*) wire P2157;
(*DONT_TOUCH="true"*) wire P2167;
(*DONT_TOUCH="true"*) wire P2207;
(*DONT_TOUCH="true"*) wire P2217;
(*DONT_TOUCH="true"*) wire P2227;
(*DONT_TOUCH="true"*) wire P2237;
(*DONT_TOUCH="true"*) wire P2247;
(*DONT_TOUCH="true"*) wire P2257;
(*DONT_TOUCH="true"*) wire P2267;
(*DONT_TOUCH="true"*) wire P2307;
(*DONT_TOUCH="true"*) wire P2317;
(*DONT_TOUCH="true"*) wire P2327;
(*DONT_TOUCH="true"*) wire P2337;
(*DONT_TOUCH="true"*) wire P2347;
(*DONT_TOUCH="true"*) wire P2357;
(*DONT_TOUCH="true"*) wire P2367;
(*DONT_TOUCH="true"*) wire P2407;
(*DONT_TOUCH="true"*) wire P2417;
(*DONT_TOUCH="true"*) wire P2427;
(*DONT_TOUCH="true"*) wire P2437;
(*DONT_TOUCH="true"*) wire P2447;
(*DONT_TOUCH="true"*) wire P2457;
(*DONT_TOUCH="true"*) wire P2467;
(*DONT_TOUCH="true"*) wire P2507;
(*DONT_TOUCH="true"*) wire P2517;
(*DONT_TOUCH="true"*) wire P2527;
(*DONT_TOUCH="true"*) wire P2537;
(*DONT_TOUCH="true"*) wire P2547;
(*DONT_TOUCH="true"*) wire P2557;
(*DONT_TOUCH="true"*) wire P2567;
(*DONT_TOUCH="true"*) wire P2607;
(*DONT_TOUCH="true"*) wire P2617;
(*DONT_TOUCH="true"*) wire P2627;
(*DONT_TOUCH="true"*) wire P2637;
(*DONT_TOUCH="true"*) wire P2647;
(*DONT_TOUCH="true"*) wire P2657;
(*DONT_TOUCH="true"*) wire P2667;
(*DONT_TOUCH="true"*) wire P3000;
(*DONT_TOUCH="true"*) wire P3010;
(*DONT_TOUCH="true"*) wire P3020;
(*DONT_TOUCH="true"*) wire P3030;
(*DONT_TOUCH="true"*) wire P3040;
(*DONT_TOUCH="true"*) wire P3100;
(*DONT_TOUCH="true"*) wire P3110;
(*DONT_TOUCH="true"*) wire P3120;
(*DONT_TOUCH="true"*) wire P3130;
(*DONT_TOUCH="true"*) wire P3140;
(*DONT_TOUCH="true"*) wire P3200;
(*DONT_TOUCH="true"*) wire P3210;
(*DONT_TOUCH="true"*) wire P3220;
(*DONT_TOUCH="true"*) wire P3230;
(*DONT_TOUCH="true"*) wire P3240;
(*DONT_TOUCH="true"*) wire P3300;
(*DONT_TOUCH="true"*) wire P3310;
(*DONT_TOUCH="true"*) wire P3320;
(*DONT_TOUCH="true"*) wire P3330;
(*DONT_TOUCH="true"*) wire P3340;
(*DONT_TOUCH="true"*) wire P3400;
(*DONT_TOUCH="true"*) wire P3410;
(*DONT_TOUCH="true"*) wire P3420;
(*DONT_TOUCH="true"*) wire P3430;
(*DONT_TOUCH="true"*) wire P3440;
(*DONT_TOUCH="true"*) wire P3001;
(*DONT_TOUCH="true"*) wire P3011;
(*DONT_TOUCH="true"*) wire P3021;
(*DONT_TOUCH="true"*) wire P3031;
(*DONT_TOUCH="true"*) wire P3041;
(*DONT_TOUCH="true"*) wire P3101;
(*DONT_TOUCH="true"*) wire P3111;
(*DONT_TOUCH="true"*) wire P3121;
(*DONT_TOUCH="true"*) wire P3131;
(*DONT_TOUCH="true"*) wire P3141;
(*DONT_TOUCH="true"*) wire P3201;
(*DONT_TOUCH="true"*) wire P3211;
(*DONT_TOUCH="true"*) wire P3221;
(*DONT_TOUCH="true"*) wire P3231;
(*DONT_TOUCH="true"*) wire P3241;
(*DONT_TOUCH="true"*) wire P3301;
(*DONT_TOUCH="true"*) wire P3311;
(*DONT_TOUCH="true"*) wire P3321;
(*DONT_TOUCH="true"*) wire P3331;
(*DONT_TOUCH="true"*) wire P3341;
(*DONT_TOUCH="true"*) wire P3401;
(*DONT_TOUCH="true"*) wire P3411;
(*DONT_TOUCH="true"*) wire P3421;
(*DONT_TOUCH="true"*) wire P3431;
(*DONT_TOUCH="true"*) wire P3441;
(*DONT_TOUCH="true"*) wire P3002;
(*DONT_TOUCH="true"*) wire P3012;
(*DONT_TOUCH="true"*) wire P3022;
(*DONT_TOUCH="true"*) wire P3032;
(*DONT_TOUCH="true"*) wire P3042;
(*DONT_TOUCH="true"*) wire P3102;
(*DONT_TOUCH="true"*) wire P3112;
(*DONT_TOUCH="true"*) wire P3122;
(*DONT_TOUCH="true"*) wire P3132;
(*DONT_TOUCH="true"*) wire P3142;
(*DONT_TOUCH="true"*) wire P3202;
(*DONT_TOUCH="true"*) wire P3212;
(*DONT_TOUCH="true"*) wire P3222;
(*DONT_TOUCH="true"*) wire P3232;
(*DONT_TOUCH="true"*) wire P3242;
(*DONT_TOUCH="true"*) wire P3302;
(*DONT_TOUCH="true"*) wire P3312;
(*DONT_TOUCH="true"*) wire P3322;
(*DONT_TOUCH="true"*) wire P3332;
(*DONT_TOUCH="true"*) wire P3342;
(*DONT_TOUCH="true"*) wire P3402;
(*DONT_TOUCH="true"*) wire P3412;
(*DONT_TOUCH="true"*) wire P3422;
(*DONT_TOUCH="true"*) wire P3432;
(*DONT_TOUCH="true"*) wire P3442;
(*DONT_TOUCH="true"*) wire P3003;
(*DONT_TOUCH="true"*) wire P3013;
(*DONT_TOUCH="true"*) wire P3023;
(*DONT_TOUCH="true"*) wire P3033;
(*DONT_TOUCH="true"*) wire P3043;
(*DONT_TOUCH="true"*) wire P3103;
(*DONT_TOUCH="true"*) wire P3113;
(*DONT_TOUCH="true"*) wire P3123;
(*DONT_TOUCH="true"*) wire P3133;
(*DONT_TOUCH="true"*) wire P3143;
(*DONT_TOUCH="true"*) wire P3203;
(*DONT_TOUCH="true"*) wire P3213;
(*DONT_TOUCH="true"*) wire P3223;
(*DONT_TOUCH="true"*) wire P3233;
(*DONT_TOUCH="true"*) wire P3243;
(*DONT_TOUCH="true"*) wire P3303;
(*DONT_TOUCH="true"*) wire P3313;
(*DONT_TOUCH="true"*) wire P3323;
(*DONT_TOUCH="true"*) wire P3333;
(*DONT_TOUCH="true"*) wire P3343;
(*DONT_TOUCH="true"*) wire P3403;
(*DONT_TOUCH="true"*) wire P3413;
(*DONT_TOUCH="true"*) wire P3423;
(*DONT_TOUCH="true"*) wire P3433;
(*DONT_TOUCH="true"*) wire P3443;
(*DONT_TOUCH="true"*) wire P3004;
(*DONT_TOUCH="true"*) wire P3014;
(*DONT_TOUCH="true"*) wire P3024;
(*DONT_TOUCH="true"*) wire P3034;
(*DONT_TOUCH="true"*) wire P3044;
(*DONT_TOUCH="true"*) wire P3104;
(*DONT_TOUCH="true"*) wire P3114;
(*DONT_TOUCH="true"*) wire P3124;
(*DONT_TOUCH="true"*) wire P3134;
(*DONT_TOUCH="true"*) wire P3144;
(*DONT_TOUCH="true"*) wire P3204;
(*DONT_TOUCH="true"*) wire P3214;
(*DONT_TOUCH="true"*) wire P3224;
(*DONT_TOUCH="true"*) wire P3234;
(*DONT_TOUCH="true"*) wire P3244;
(*DONT_TOUCH="true"*) wire P3304;
(*DONT_TOUCH="true"*) wire P3314;
(*DONT_TOUCH="true"*) wire P3324;
(*DONT_TOUCH="true"*) wire P3334;
(*DONT_TOUCH="true"*) wire P3344;
(*DONT_TOUCH="true"*) wire P3404;
(*DONT_TOUCH="true"*) wire P3414;
(*DONT_TOUCH="true"*) wire P3424;
(*DONT_TOUCH="true"*) wire P3434;
(*DONT_TOUCH="true"*) wire P3444;
(*DONT_TOUCH="true"*) wire P3005;
(*DONT_TOUCH="true"*) wire P3015;
(*DONT_TOUCH="true"*) wire P3025;
(*DONT_TOUCH="true"*) wire P3035;
(*DONT_TOUCH="true"*) wire P3045;
(*DONT_TOUCH="true"*) wire P3105;
(*DONT_TOUCH="true"*) wire P3115;
(*DONT_TOUCH="true"*) wire P3125;
(*DONT_TOUCH="true"*) wire P3135;
(*DONT_TOUCH="true"*) wire P3145;
(*DONT_TOUCH="true"*) wire P3205;
(*DONT_TOUCH="true"*) wire P3215;
(*DONT_TOUCH="true"*) wire P3225;
(*DONT_TOUCH="true"*) wire P3235;
(*DONT_TOUCH="true"*) wire P3245;
(*DONT_TOUCH="true"*) wire P3305;
(*DONT_TOUCH="true"*) wire P3315;
(*DONT_TOUCH="true"*) wire P3325;
(*DONT_TOUCH="true"*) wire P3335;
(*DONT_TOUCH="true"*) wire P3345;
(*DONT_TOUCH="true"*) wire P3405;
(*DONT_TOUCH="true"*) wire P3415;
(*DONT_TOUCH="true"*) wire P3425;
(*DONT_TOUCH="true"*) wire P3435;
(*DONT_TOUCH="true"*) wire P3445;
(*DONT_TOUCH="true"*) wire P3006;
(*DONT_TOUCH="true"*) wire P3016;
(*DONT_TOUCH="true"*) wire P3026;
(*DONT_TOUCH="true"*) wire P3036;
(*DONT_TOUCH="true"*) wire P3046;
(*DONT_TOUCH="true"*) wire P3106;
(*DONT_TOUCH="true"*) wire P3116;
(*DONT_TOUCH="true"*) wire P3126;
(*DONT_TOUCH="true"*) wire P3136;
(*DONT_TOUCH="true"*) wire P3146;
(*DONT_TOUCH="true"*) wire P3206;
(*DONT_TOUCH="true"*) wire P3216;
(*DONT_TOUCH="true"*) wire P3226;
(*DONT_TOUCH="true"*) wire P3236;
(*DONT_TOUCH="true"*) wire P3246;
(*DONT_TOUCH="true"*) wire P3306;
(*DONT_TOUCH="true"*) wire P3316;
(*DONT_TOUCH="true"*) wire P3326;
(*DONT_TOUCH="true"*) wire P3336;
(*DONT_TOUCH="true"*) wire P3346;
(*DONT_TOUCH="true"*) wire P3406;
(*DONT_TOUCH="true"*) wire P3416;
(*DONT_TOUCH="true"*) wire P3426;
(*DONT_TOUCH="true"*) wire P3436;
(*DONT_TOUCH="true"*) wire P3446;
(*DONT_TOUCH="true"*) wire P3007;
(*DONT_TOUCH="true"*) wire P3017;
(*DONT_TOUCH="true"*) wire P3027;
(*DONT_TOUCH="true"*) wire P3037;
(*DONT_TOUCH="true"*) wire P3047;
(*DONT_TOUCH="true"*) wire P3107;
(*DONT_TOUCH="true"*) wire P3117;
(*DONT_TOUCH="true"*) wire P3127;
(*DONT_TOUCH="true"*) wire P3137;
(*DONT_TOUCH="true"*) wire P3147;
(*DONT_TOUCH="true"*) wire P3207;
(*DONT_TOUCH="true"*) wire P3217;
(*DONT_TOUCH="true"*) wire P3227;
(*DONT_TOUCH="true"*) wire P3237;
(*DONT_TOUCH="true"*) wire P3247;
(*DONT_TOUCH="true"*) wire P3307;
(*DONT_TOUCH="true"*) wire P3317;
(*DONT_TOUCH="true"*) wire P3327;
(*DONT_TOUCH="true"*) wire P3337;
(*DONT_TOUCH="true"*) wire P3347;
(*DONT_TOUCH="true"*) wire P3407;
(*DONT_TOUCH="true"*) wire P3417;
(*DONT_TOUCH="true"*) wire P3427;
(*DONT_TOUCH="true"*) wire P3437;
(*DONT_TOUCH="true"*) wire P3447;
(*DONT_TOUCH="true"*) wire P3008;
(*DONT_TOUCH="true"*) wire P3018;
(*DONT_TOUCH="true"*) wire P3028;
(*DONT_TOUCH="true"*) wire P3038;
(*DONT_TOUCH="true"*) wire P3048;
(*DONT_TOUCH="true"*) wire P3108;
(*DONT_TOUCH="true"*) wire P3118;
(*DONT_TOUCH="true"*) wire P3128;
(*DONT_TOUCH="true"*) wire P3138;
(*DONT_TOUCH="true"*) wire P3148;
(*DONT_TOUCH="true"*) wire P3208;
(*DONT_TOUCH="true"*) wire P3218;
(*DONT_TOUCH="true"*) wire P3228;
(*DONT_TOUCH="true"*) wire P3238;
(*DONT_TOUCH="true"*) wire P3248;
(*DONT_TOUCH="true"*) wire P3308;
(*DONT_TOUCH="true"*) wire P3318;
(*DONT_TOUCH="true"*) wire P3328;
(*DONT_TOUCH="true"*) wire P3338;
(*DONT_TOUCH="true"*) wire P3348;
(*DONT_TOUCH="true"*) wire P3408;
(*DONT_TOUCH="true"*) wire P3418;
(*DONT_TOUCH="true"*) wire P3428;
(*DONT_TOUCH="true"*) wire P3438;
(*DONT_TOUCH="true"*) wire P3448;
(*DONT_TOUCH="true"*) wire P3009;
(*DONT_TOUCH="true"*) wire P3019;
(*DONT_TOUCH="true"*) wire P3029;
(*DONT_TOUCH="true"*) wire P3039;
(*DONT_TOUCH="true"*) wire P3049;
(*DONT_TOUCH="true"*) wire P3109;
(*DONT_TOUCH="true"*) wire P3119;
(*DONT_TOUCH="true"*) wire P3129;
(*DONT_TOUCH="true"*) wire P3139;
(*DONT_TOUCH="true"*) wire P3149;
(*DONT_TOUCH="true"*) wire P3209;
(*DONT_TOUCH="true"*) wire P3219;
(*DONT_TOUCH="true"*) wire P3229;
(*DONT_TOUCH="true"*) wire P3239;
(*DONT_TOUCH="true"*) wire P3249;
(*DONT_TOUCH="true"*) wire P3309;
(*DONT_TOUCH="true"*) wire P3319;
(*DONT_TOUCH="true"*) wire P3329;
(*DONT_TOUCH="true"*) wire P3339;
(*DONT_TOUCH="true"*) wire P3349;
(*DONT_TOUCH="true"*) wire P3409;
(*DONT_TOUCH="true"*) wire P3419;
(*DONT_TOUCH="true"*) wire P3429;
(*DONT_TOUCH="true"*) wire P3439;
(*DONT_TOUCH="true"*) wire P3449;
(*DONT_TOUCH="true"*) wire P300A;
(*DONT_TOUCH="true"*) wire P301A;
(*DONT_TOUCH="true"*) wire P302A;
(*DONT_TOUCH="true"*) wire P303A;
(*DONT_TOUCH="true"*) wire P304A;
(*DONT_TOUCH="true"*) wire P310A;
(*DONT_TOUCH="true"*) wire P311A;
(*DONT_TOUCH="true"*) wire P312A;
(*DONT_TOUCH="true"*) wire P313A;
(*DONT_TOUCH="true"*) wire P314A;
(*DONT_TOUCH="true"*) wire P320A;
(*DONT_TOUCH="true"*) wire P321A;
(*DONT_TOUCH="true"*) wire P322A;
(*DONT_TOUCH="true"*) wire P323A;
(*DONT_TOUCH="true"*) wire P324A;
(*DONT_TOUCH="true"*) wire P330A;
(*DONT_TOUCH="true"*) wire P331A;
(*DONT_TOUCH="true"*) wire P332A;
(*DONT_TOUCH="true"*) wire P333A;
(*DONT_TOUCH="true"*) wire P334A;
(*DONT_TOUCH="true"*) wire P340A;
(*DONT_TOUCH="true"*) wire P341A;
(*DONT_TOUCH="true"*) wire P342A;
(*DONT_TOUCH="true"*) wire P343A;
(*DONT_TOUCH="true"*) wire P344A;
(*DONT_TOUCH="true"*) wire P300B;
(*DONT_TOUCH="true"*) wire P301B;
(*DONT_TOUCH="true"*) wire P302B;
(*DONT_TOUCH="true"*) wire P303B;
(*DONT_TOUCH="true"*) wire P304B;
(*DONT_TOUCH="true"*) wire P310B;
(*DONT_TOUCH="true"*) wire P311B;
(*DONT_TOUCH="true"*) wire P312B;
(*DONT_TOUCH="true"*) wire P313B;
(*DONT_TOUCH="true"*) wire P314B;
(*DONT_TOUCH="true"*) wire P320B;
(*DONT_TOUCH="true"*) wire P321B;
(*DONT_TOUCH="true"*) wire P322B;
(*DONT_TOUCH="true"*) wire P323B;
(*DONT_TOUCH="true"*) wire P324B;
(*DONT_TOUCH="true"*) wire P330B;
(*DONT_TOUCH="true"*) wire P331B;
(*DONT_TOUCH="true"*) wire P332B;
(*DONT_TOUCH="true"*) wire P333B;
(*DONT_TOUCH="true"*) wire P334B;
(*DONT_TOUCH="true"*) wire P340B;
(*DONT_TOUCH="true"*) wire P341B;
(*DONT_TOUCH="true"*) wire P342B;
(*DONT_TOUCH="true"*) wire P343B;
(*DONT_TOUCH="true"*) wire P344B;
(*DONT_TOUCH="true"*) wire P300C;
(*DONT_TOUCH="true"*) wire P301C;
(*DONT_TOUCH="true"*) wire P302C;
(*DONT_TOUCH="true"*) wire P303C;
(*DONT_TOUCH="true"*) wire P304C;
(*DONT_TOUCH="true"*) wire P310C;
(*DONT_TOUCH="true"*) wire P311C;
(*DONT_TOUCH="true"*) wire P312C;
(*DONT_TOUCH="true"*) wire P313C;
(*DONT_TOUCH="true"*) wire P314C;
(*DONT_TOUCH="true"*) wire P320C;
(*DONT_TOUCH="true"*) wire P321C;
(*DONT_TOUCH="true"*) wire P322C;
(*DONT_TOUCH="true"*) wire P323C;
(*DONT_TOUCH="true"*) wire P324C;
(*DONT_TOUCH="true"*) wire P330C;
(*DONT_TOUCH="true"*) wire P331C;
(*DONT_TOUCH="true"*) wire P332C;
(*DONT_TOUCH="true"*) wire P333C;
(*DONT_TOUCH="true"*) wire P334C;
(*DONT_TOUCH="true"*) wire P340C;
(*DONT_TOUCH="true"*) wire P341C;
(*DONT_TOUCH="true"*) wire P342C;
(*DONT_TOUCH="true"*) wire P343C;
(*DONT_TOUCH="true"*) wire P344C;
(*DONT_TOUCH="true"*) wire P300D;
(*DONT_TOUCH="true"*) wire P301D;
(*DONT_TOUCH="true"*) wire P302D;
(*DONT_TOUCH="true"*) wire P303D;
(*DONT_TOUCH="true"*) wire P304D;
(*DONT_TOUCH="true"*) wire P310D;
(*DONT_TOUCH="true"*) wire P311D;
(*DONT_TOUCH="true"*) wire P312D;
(*DONT_TOUCH="true"*) wire P313D;
(*DONT_TOUCH="true"*) wire P314D;
(*DONT_TOUCH="true"*) wire P320D;
(*DONT_TOUCH="true"*) wire P321D;
(*DONT_TOUCH="true"*) wire P322D;
(*DONT_TOUCH="true"*) wire P323D;
(*DONT_TOUCH="true"*) wire P324D;
(*DONT_TOUCH="true"*) wire P330D;
(*DONT_TOUCH="true"*) wire P331D;
(*DONT_TOUCH="true"*) wire P332D;
(*DONT_TOUCH="true"*) wire P333D;
(*DONT_TOUCH="true"*) wire P334D;
(*DONT_TOUCH="true"*) wire P340D;
(*DONT_TOUCH="true"*) wire P341D;
(*DONT_TOUCH="true"*) wire P342D;
(*DONT_TOUCH="true"*) wire P343D;
(*DONT_TOUCH="true"*) wire P344D;
(*DONT_TOUCH="true"*) wire P300E;
(*DONT_TOUCH="true"*) wire P301E;
(*DONT_TOUCH="true"*) wire P302E;
(*DONT_TOUCH="true"*) wire P303E;
(*DONT_TOUCH="true"*) wire P304E;
(*DONT_TOUCH="true"*) wire P310E;
(*DONT_TOUCH="true"*) wire P311E;
(*DONT_TOUCH="true"*) wire P312E;
(*DONT_TOUCH="true"*) wire P313E;
(*DONT_TOUCH="true"*) wire P314E;
(*DONT_TOUCH="true"*) wire P320E;
(*DONT_TOUCH="true"*) wire P321E;
(*DONT_TOUCH="true"*) wire P322E;
(*DONT_TOUCH="true"*) wire P323E;
(*DONT_TOUCH="true"*) wire P324E;
(*DONT_TOUCH="true"*) wire P330E;
(*DONT_TOUCH="true"*) wire P331E;
(*DONT_TOUCH="true"*) wire P332E;
(*DONT_TOUCH="true"*) wire P333E;
(*DONT_TOUCH="true"*) wire P334E;
(*DONT_TOUCH="true"*) wire P340E;
(*DONT_TOUCH="true"*) wire P341E;
(*DONT_TOUCH="true"*) wire P342E;
(*DONT_TOUCH="true"*) wire P343E;
(*DONT_TOUCH="true"*) wire P344E;
(*DONT_TOUCH="true"*) wire P300F;
(*DONT_TOUCH="true"*) wire P301F;
(*DONT_TOUCH="true"*) wire P302F;
(*DONT_TOUCH="true"*) wire P303F;
(*DONT_TOUCH="true"*) wire P304F;
(*DONT_TOUCH="true"*) wire P310F;
(*DONT_TOUCH="true"*) wire P311F;
(*DONT_TOUCH="true"*) wire P312F;
(*DONT_TOUCH="true"*) wire P313F;
(*DONT_TOUCH="true"*) wire P314F;
(*DONT_TOUCH="true"*) wire P320F;
(*DONT_TOUCH="true"*) wire P321F;
(*DONT_TOUCH="true"*) wire P322F;
(*DONT_TOUCH="true"*) wire P323F;
(*DONT_TOUCH="true"*) wire P324F;
(*DONT_TOUCH="true"*) wire P330F;
(*DONT_TOUCH="true"*) wire P331F;
(*DONT_TOUCH="true"*) wire P332F;
(*DONT_TOUCH="true"*) wire P333F;
(*DONT_TOUCH="true"*) wire P334F;
(*DONT_TOUCH="true"*) wire P340F;
(*DONT_TOUCH="true"*) wire P341F;
(*DONT_TOUCH="true"*) wire P342F;
(*DONT_TOUCH="true"*) wire P343F;
(*DONT_TOUCH="true"*) wire P344F;
(*DONT_TOUCH="true"*) wire W20000,W20010,W20020,W20100,W20110,W20120,W20200,W20210,W20220;
(*DONT_TOUCH="true"*) wire W20001,W20011,W20021,W20101,W20111,W20121,W20201,W20211,W20221;
(*DONT_TOUCH="true"*) wire W20002,W20012,W20022,W20102,W20112,W20122,W20202,W20212,W20222;
(*DONT_TOUCH="true"*) wire W20003,W20013,W20023,W20103,W20113,W20123,W20203,W20213,W20223;
(*DONT_TOUCH="true"*) wire W20004,W20014,W20024,W20104,W20114,W20124,W20204,W20214,W20224;
(*DONT_TOUCH="true"*) wire W20005,W20015,W20025,W20105,W20115,W20125,W20205,W20215,W20225;
(*DONT_TOUCH="true"*) wire W20006,W20016,W20026,W20106,W20116,W20126,W20206,W20216,W20226;
(*DONT_TOUCH="true"*) wire W20007,W20017,W20027,W20107,W20117,W20127,W20207,W20217,W20227;
(*DONT_TOUCH="true"*) wire W21000,W21010,W21020,W21100,W21110,W21120,W21200,W21210,W21220;
(*DONT_TOUCH="true"*) wire W21001,W21011,W21021,W21101,W21111,W21121,W21201,W21211,W21221;
(*DONT_TOUCH="true"*) wire W21002,W21012,W21022,W21102,W21112,W21122,W21202,W21212,W21222;
(*DONT_TOUCH="true"*) wire W21003,W21013,W21023,W21103,W21113,W21123,W21203,W21213,W21223;
(*DONT_TOUCH="true"*) wire W21004,W21014,W21024,W21104,W21114,W21124,W21204,W21214,W21224;
(*DONT_TOUCH="true"*) wire W21005,W21015,W21025,W21105,W21115,W21125,W21205,W21215,W21225;
(*DONT_TOUCH="true"*) wire W21006,W21016,W21026,W21106,W21116,W21126,W21206,W21216,W21226;
(*DONT_TOUCH="true"*) wire W21007,W21017,W21027,W21107,W21117,W21127,W21207,W21217,W21227;
(*DONT_TOUCH="true"*) wire W22000,W22010,W22020,W22100,W22110,W22120,W22200,W22210,W22220;
(*DONT_TOUCH="true"*) wire W22001,W22011,W22021,W22101,W22111,W22121,W22201,W22211,W22221;
(*DONT_TOUCH="true"*) wire W22002,W22012,W22022,W22102,W22112,W22122,W22202,W22212,W22222;
(*DONT_TOUCH="true"*) wire W22003,W22013,W22023,W22103,W22113,W22123,W22203,W22213,W22223;
(*DONT_TOUCH="true"*) wire W22004,W22014,W22024,W22104,W22114,W22124,W22204,W22214,W22224;
(*DONT_TOUCH="true"*) wire W22005,W22015,W22025,W22105,W22115,W22125,W22205,W22215,W22225;
(*DONT_TOUCH="true"*) wire W22006,W22016,W22026,W22106,W22116,W22126,W22206,W22216,W22226;
(*DONT_TOUCH="true"*) wire W22007,W22017,W22027,W22107,W22117,W22127,W22207,W22217,W22227;
(*DONT_TOUCH="true"*) wire W23000,W23010,W23020,W23100,W23110,W23120,W23200,W23210,W23220;
(*DONT_TOUCH="true"*) wire W23001,W23011,W23021,W23101,W23111,W23121,W23201,W23211,W23221;
(*DONT_TOUCH="true"*) wire W23002,W23012,W23022,W23102,W23112,W23122,W23202,W23212,W23222;
(*DONT_TOUCH="true"*) wire W23003,W23013,W23023,W23103,W23113,W23123,W23203,W23213,W23223;
(*DONT_TOUCH="true"*) wire W23004,W23014,W23024,W23104,W23114,W23124,W23204,W23214,W23224;
(*DONT_TOUCH="true"*) wire W23005,W23015,W23025,W23105,W23115,W23125,W23205,W23215,W23225;
(*DONT_TOUCH="true"*) wire W23006,W23016,W23026,W23106,W23116,W23126,W23206,W23216,W23226;
(*DONT_TOUCH="true"*) wire W23007,W23017,W23027,W23107,W23117,W23127,W23207,W23217,W23227;
(*DONT_TOUCH="true"*) wire W24000,W24010,W24020,W24100,W24110,W24120,W24200,W24210,W24220;
(*DONT_TOUCH="true"*) wire W24001,W24011,W24021,W24101,W24111,W24121,W24201,W24211,W24221;
(*DONT_TOUCH="true"*) wire W24002,W24012,W24022,W24102,W24112,W24122,W24202,W24212,W24222;
(*DONT_TOUCH="true"*) wire W24003,W24013,W24023,W24103,W24113,W24123,W24203,W24213,W24223;
(*DONT_TOUCH="true"*) wire W24004,W24014,W24024,W24104,W24114,W24124,W24204,W24214,W24224;
(*DONT_TOUCH="true"*) wire W24005,W24015,W24025,W24105,W24115,W24125,W24205,W24215,W24225;
(*DONT_TOUCH="true"*) wire W24006,W24016,W24026,W24106,W24116,W24126,W24206,W24216,W24226;
(*DONT_TOUCH="true"*) wire W24007,W24017,W24027,W24107,W24117,W24127,W24207,W24217,W24227;
(*DONT_TOUCH="true"*) wire W25000,W25010,W25020,W25100,W25110,W25120,W25200,W25210,W25220;
(*DONT_TOUCH="true"*) wire W25001,W25011,W25021,W25101,W25111,W25121,W25201,W25211,W25221;
(*DONT_TOUCH="true"*) wire W25002,W25012,W25022,W25102,W25112,W25122,W25202,W25212,W25222;
(*DONT_TOUCH="true"*) wire W25003,W25013,W25023,W25103,W25113,W25123,W25203,W25213,W25223;
(*DONT_TOUCH="true"*) wire W25004,W25014,W25024,W25104,W25114,W25124,W25204,W25214,W25224;
(*DONT_TOUCH="true"*) wire W25005,W25015,W25025,W25105,W25115,W25125,W25205,W25215,W25225;
(*DONT_TOUCH="true"*) wire W25006,W25016,W25026,W25106,W25116,W25126,W25206,W25216,W25226;
(*DONT_TOUCH="true"*) wire W25007,W25017,W25027,W25107,W25117,W25127,W25207,W25217,W25227;
(*DONT_TOUCH="true"*) wire W26000,W26010,W26020,W26100,W26110,W26120,W26200,W26210,W26220;
(*DONT_TOUCH="true"*) wire W26001,W26011,W26021,W26101,W26111,W26121,W26201,W26211,W26221;
(*DONT_TOUCH="true"*) wire W26002,W26012,W26022,W26102,W26112,W26122,W26202,W26212,W26222;
(*DONT_TOUCH="true"*) wire W26003,W26013,W26023,W26103,W26113,W26123,W26203,W26213,W26223;
(*DONT_TOUCH="true"*) wire W26004,W26014,W26024,W26104,W26114,W26124,W26204,W26214,W26224;
(*DONT_TOUCH="true"*) wire W26005,W26015,W26025,W26105,W26115,W26125,W26205,W26215,W26225;
(*DONT_TOUCH="true"*) wire W26006,W26016,W26026,W26106,W26116,W26126,W26206,W26216,W26226;
(*DONT_TOUCH="true"*) wire W26007,W26017,W26027,W26107,W26117,W26127,W26207,W26217,W26227;
(*DONT_TOUCH="true"*) wire W27000,W27010,W27020,W27100,W27110,W27120,W27200,W27210,W27220;
(*DONT_TOUCH="true"*) wire W27001,W27011,W27021,W27101,W27111,W27121,W27201,W27211,W27221;
(*DONT_TOUCH="true"*) wire W27002,W27012,W27022,W27102,W27112,W27122,W27202,W27212,W27222;
(*DONT_TOUCH="true"*) wire W27003,W27013,W27023,W27103,W27113,W27123,W27203,W27213,W27223;
(*DONT_TOUCH="true"*) wire W27004,W27014,W27024,W27104,W27114,W27124,W27204,W27214,W27224;
(*DONT_TOUCH="true"*) wire W27005,W27015,W27025,W27105,W27115,W27125,W27205,W27215,W27225;
(*DONT_TOUCH="true"*) wire W27006,W27016,W27026,W27106,W27116,W27126,W27206,W27216,W27226;
(*DONT_TOUCH="true"*) wire W27007,W27017,W27027,W27107,W27117,W27127,W27207,W27217,W27227;
(*DONT_TOUCH="true"*) wire W28000,W28010,W28020,W28100,W28110,W28120,W28200,W28210,W28220;
(*DONT_TOUCH="true"*) wire W28001,W28011,W28021,W28101,W28111,W28121,W28201,W28211,W28221;
(*DONT_TOUCH="true"*) wire W28002,W28012,W28022,W28102,W28112,W28122,W28202,W28212,W28222;
(*DONT_TOUCH="true"*) wire W28003,W28013,W28023,W28103,W28113,W28123,W28203,W28213,W28223;
(*DONT_TOUCH="true"*) wire W28004,W28014,W28024,W28104,W28114,W28124,W28204,W28214,W28224;
(*DONT_TOUCH="true"*) wire W28005,W28015,W28025,W28105,W28115,W28125,W28205,W28215,W28225;
(*DONT_TOUCH="true"*) wire W28006,W28016,W28026,W28106,W28116,W28126,W28206,W28216,W28226;
(*DONT_TOUCH="true"*) wire W28007,W28017,W28027,W28107,W28117,W28127,W28207,W28217,W28227;
(*DONT_TOUCH="true"*) wire W29000,W29010,W29020,W29100,W29110,W29120,W29200,W29210,W29220;
(*DONT_TOUCH="true"*) wire W29001,W29011,W29021,W29101,W29111,W29121,W29201,W29211,W29221;
(*DONT_TOUCH="true"*) wire W29002,W29012,W29022,W29102,W29112,W29122,W29202,W29212,W29222;
(*DONT_TOUCH="true"*) wire W29003,W29013,W29023,W29103,W29113,W29123,W29203,W29213,W29223;
(*DONT_TOUCH="true"*) wire W29004,W29014,W29024,W29104,W29114,W29124,W29204,W29214,W29224;
(*DONT_TOUCH="true"*) wire W29005,W29015,W29025,W29105,W29115,W29125,W29205,W29215,W29225;
(*DONT_TOUCH="true"*) wire W29006,W29016,W29026,W29106,W29116,W29126,W29206,W29216,W29226;
(*DONT_TOUCH="true"*) wire W29007,W29017,W29027,W29107,W29117,W29127,W29207,W29217,W29227;
(*DONT_TOUCH="true"*) wire W2A000,W2A010,W2A020,W2A100,W2A110,W2A120,W2A200,W2A210,W2A220;
(*DONT_TOUCH="true"*) wire W2A001,W2A011,W2A021,W2A101,W2A111,W2A121,W2A201,W2A211,W2A221;
(*DONT_TOUCH="true"*) wire W2A002,W2A012,W2A022,W2A102,W2A112,W2A122,W2A202,W2A212,W2A222;
(*DONT_TOUCH="true"*) wire W2A003,W2A013,W2A023,W2A103,W2A113,W2A123,W2A203,W2A213,W2A223;
(*DONT_TOUCH="true"*) wire W2A004,W2A014,W2A024,W2A104,W2A114,W2A124,W2A204,W2A214,W2A224;
(*DONT_TOUCH="true"*) wire W2A005,W2A015,W2A025,W2A105,W2A115,W2A125,W2A205,W2A215,W2A225;
(*DONT_TOUCH="true"*) wire W2A006,W2A016,W2A026,W2A106,W2A116,W2A126,W2A206,W2A216,W2A226;
(*DONT_TOUCH="true"*) wire W2A007,W2A017,W2A027,W2A107,W2A117,W2A127,W2A207,W2A217,W2A227;
(*DONT_TOUCH="true"*) wire W2B000,W2B010,W2B020,W2B100,W2B110,W2B120,W2B200,W2B210,W2B220;
(*DONT_TOUCH="true"*) wire W2B001,W2B011,W2B021,W2B101,W2B111,W2B121,W2B201,W2B211,W2B221;
(*DONT_TOUCH="true"*) wire W2B002,W2B012,W2B022,W2B102,W2B112,W2B122,W2B202,W2B212,W2B222;
(*DONT_TOUCH="true"*) wire W2B003,W2B013,W2B023,W2B103,W2B113,W2B123,W2B203,W2B213,W2B223;
(*DONT_TOUCH="true"*) wire W2B004,W2B014,W2B024,W2B104,W2B114,W2B124,W2B204,W2B214,W2B224;
(*DONT_TOUCH="true"*) wire W2B005,W2B015,W2B025,W2B105,W2B115,W2B125,W2B205,W2B215,W2B225;
(*DONT_TOUCH="true"*) wire W2B006,W2B016,W2B026,W2B106,W2B116,W2B126,W2B206,W2B216,W2B226;
(*DONT_TOUCH="true"*) wire W2B007,W2B017,W2B027,W2B107,W2B117,W2B127,W2B207,W2B217,W2B227;
(*DONT_TOUCH="true"*) wire W2C000,W2C010,W2C020,W2C100,W2C110,W2C120,W2C200,W2C210,W2C220;
(*DONT_TOUCH="true"*) wire W2C001,W2C011,W2C021,W2C101,W2C111,W2C121,W2C201,W2C211,W2C221;
(*DONT_TOUCH="true"*) wire W2C002,W2C012,W2C022,W2C102,W2C112,W2C122,W2C202,W2C212,W2C222;
(*DONT_TOUCH="true"*) wire W2C003,W2C013,W2C023,W2C103,W2C113,W2C123,W2C203,W2C213,W2C223;
(*DONT_TOUCH="true"*) wire W2C004,W2C014,W2C024,W2C104,W2C114,W2C124,W2C204,W2C214,W2C224;
(*DONT_TOUCH="true"*) wire W2C005,W2C015,W2C025,W2C105,W2C115,W2C125,W2C205,W2C215,W2C225;
(*DONT_TOUCH="true"*) wire W2C006,W2C016,W2C026,W2C106,W2C116,W2C126,W2C206,W2C216,W2C226;
(*DONT_TOUCH="true"*) wire W2C007,W2C017,W2C027,W2C107,W2C117,W2C127,W2C207,W2C217,W2C227;
(*DONT_TOUCH="true"*) wire W2D000,W2D010,W2D020,W2D100,W2D110,W2D120,W2D200,W2D210,W2D220;
(*DONT_TOUCH="true"*) wire W2D001,W2D011,W2D021,W2D101,W2D111,W2D121,W2D201,W2D211,W2D221;
(*DONT_TOUCH="true"*) wire W2D002,W2D012,W2D022,W2D102,W2D112,W2D122,W2D202,W2D212,W2D222;
(*DONT_TOUCH="true"*) wire W2D003,W2D013,W2D023,W2D103,W2D113,W2D123,W2D203,W2D213,W2D223;
(*DONT_TOUCH="true"*) wire W2D004,W2D014,W2D024,W2D104,W2D114,W2D124,W2D204,W2D214,W2D224;
(*DONT_TOUCH="true"*) wire W2D005,W2D015,W2D025,W2D105,W2D115,W2D125,W2D205,W2D215,W2D225;
(*DONT_TOUCH="true"*) wire W2D006,W2D016,W2D026,W2D106,W2D116,W2D126,W2D206,W2D216,W2D226;
(*DONT_TOUCH="true"*) wire W2D007,W2D017,W2D027,W2D107,W2D117,W2D127,W2D207,W2D217,W2D227;
(*DONT_TOUCH="true"*) wire W2E000,W2E010,W2E020,W2E100,W2E110,W2E120,W2E200,W2E210,W2E220;
(*DONT_TOUCH="true"*) wire W2E001,W2E011,W2E021,W2E101,W2E111,W2E121,W2E201,W2E211,W2E221;
(*DONT_TOUCH="true"*) wire W2E002,W2E012,W2E022,W2E102,W2E112,W2E122,W2E202,W2E212,W2E222;
(*DONT_TOUCH="true"*) wire W2E003,W2E013,W2E023,W2E103,W2E113,W2E123,W2E203,W2E213,W2E223;
(*DONT_TOUCH="true"*) wire W2E004,W2E014,W2E024,W2E104,W2E114,W2E124,W2E204,W2E214,W2E224;
(*DONT_TOUCH="true"*) wire W2E005,W2E015,W2E025,W2E105,W2E115,W2E125,W2E205,W2E215,W2E225;
(*DONT_TOUCH="true"*) wire W2E006,W2E016,W2E026,W2E106,W2E116,W2E126,W2E206,W2E216,W2E226;
(*DONT_TOUCH="true"*) wire W2E007,W2E017,W2E027,W2E107,W2E117,W2E127,W2E207,W2E217,W2E227;
(*DONT_TOUCH="true"*) wire W2F000,W2F010,W2F020,W2F100,W2F110,W2F120,W2F200,W2F210,W2F220;
(*DONT_TOUCH="true"*) wire W2F001,W2F011,W2F021,W2F101,W2F111,W2F121,W2F201,W2F211,W2F221;
(*DONT_TOUCH="true"*) wire W2F002,W2F012,W2F022,W2F102,W2F112,W2F122,W2F202,W2F212,W2F222;
(*DONT_TOUCH="true"*) wire W2F003,W2F013,W2F023,W2F103,W2F113,W2F123,W2F203,W2F213,W2F223;
(*DONT_TOUCH="true"*) wire W2F004,W2F014,W2F024,W2F104,W2F114,W2F124,W2F204,W2F214,W2F224;
(*DONT_TOUCH="true"*) wire W2F005,W2F015,W2F025,W2F105,W2F115,W2F125,W2F205,W2F215,W2F225;
(*DONT_TOUCH="true"*) wire W2F006,W2F016,W2F026,W2F106,W2F116,W2F126,W2F206,W2F216,W2F226;
(*DONT_TOUCH="true"*) wire W2F007,W2F017,W2F027,W2F107,W2F117,W2F127,W2F207,W2F217,W2F227;
(*DONT_TOUCH="true"*) wire signed [4:0] c20000,c21000,c22000,c23000,c24000,c25000,c26000,c27000;
(*DONT_TOUCH="true"*) wire signed [4:0] c20010,c21010,c22010,c23010,c24010,c25010,c26010,c27010;
(*DONT_TOUCH="true"*) wire signed [4:0] c20020,c21020,c22020,c23020,c24020,c25020,c26020,c27020;
(*DONT_TOUCH="true"*) wire signed [4:0] c20030,c21030,c22030,c23030,c24030,c25030,c26030,c27030;
(*DONT_TOUCH="true"*) wire signed [4:0] c20040,c21040,c22040,c23040,c24040,c25040,c26040,c27040;
(*DONT_TOUCH="true"*) wire signed [4:0] c20100,c21100,c22100,c23100,c24100,c25100,c26100,c27100;
(*DONT_TOUCH="true"*) wire signed [4:0] c20110,c21110,c22110,c23110,c24110,c25110,c26110,c27110;
(*DONT_TOUCH="true"*) wire signed [4:0] c20120,c21120,c22120,c23120,c24120,c25120,c26120,c27120;
(*DONT_TOUCH="true"*) wire signed [4:0] c20130,c21130,c22130,c23130,c24130,c25130,c26130,c27130;
(*DONT_TOUCH="true"*) wire signed [4:0] c20140,c21140,c22140,c23140,c24140,c25140,c26140,c27140;
(*DONT_TOUCH="true"*) wire signed [4:0] c20200,c21200,c22200,c23200,c24200,c25200,c26200,c27200;
(*DONT_TOUCH="true"*) wire signed [4:0] c20210,c21210,c22210,c23210,c24210,c25210,c26210,c27210;
(*DONT_TOUCH="true"*) wire signed [4:0] c20220,c21220,c22220,c23220,c24220,c25220,c26220,c27220;
(*DONT_TOUCH="true"*) wire signed [4:0] c20230,c21230,c22230,c23230,c24230,c25230,c26230,c27230;
(*DONT_TOUCH="true"*) wire signed [4:0] c20240,c21240,c22240,c23240,c24240,c25240,c26240,c27240;
(*DONT_TOUCH="true"*) wire signed [4:0] c20300,c21300,c22300,c23300,c24300,c25300,c26300,c27300;
(*DONT_TOUCH="true"*) wire signed [4:0] c20310,c21310,c22310,c23310,c24310,c25310,c26310,c27310;
(*DONT_TOUCH="true"*) wire signed [4:0] c20320,c21320,c22320,c23320,c24320,c25320,c26320,c27320;
(*DONT_TOUCH="true"*) wire signed [4:0] c20330,c21330,c22330,c23330,c24330,c25330,c26330,c27330;
(*DONT_TOUCH="true"*) wire signed [4:0] c20340,c21340,c22340,c23340,c24340,c25340,c26340,c27340;
(*DONT_TOUCH="true"*) wire signed [4:0] c20400,c21400,c22400,c23400,c24400,c25400,c26400,c27400;
(*DONT_TOUCH="true"*) wire signed [4:0] c20410,c21410,c22410,c23410,c24410,c25410,c26410,c27410;
(*DONT_TOUCH="true"*) wire signed [4:0] c20420,c21420,c22420,c23420,c24420,c25420,c26420,c27420;
(*DONT_TOUCH="true"*) wire signed [4:0] c20430,c21430,c22430,c23430,c24430,c25430,c26430,c27430;
(*DONT_TOUCH="true"*) wire signed [4:0] c20440,c21440,c22440,c23440,c24440,c25440,c26440,c27440;
(*DONT_TOUCH="true"*) wire signed [4:0] c20001,c21001,c22001,c23001,c24001,c25001,c26001,c27001;
(*DONT_TOUCH="true"*) wire signed [4:0] c20011,c21011,c22011,c23011,c24011,c25011,c26011,c27011;
(*DONT_TOUCH="true"*) wire signed [4:0] c20021,c21021,c22021,c23021,c24021,c25021,c26021,c27021;
(*DONT_TOUCH="true"*) wire signed [4:0] c20031,c21031,c22031,c23031,c24031,c25031,c26031,c27031;
(*DONT_TOUCH="true"*) wire signed [4:0] c20041,c21041,c22041,c23041,c24041,c25041,c26041,c27041;
(*DONT_TOUCH="true"*) wire signed [4:0] c20101,c21101,c22101,c23101,c24101,c25101,c26101,c27101;
(*DONT_TOUCH="true"*) wire signed [4:0] c20111,c21111,c22111,c23111,c24111,c25111,c26111,c27111;
(*DONT_TOUCH="true"*) wire signed [4:0] c20121,c21121,c22121,c23121,c24121,c25121,c26121,c27121;
(*DONT_TOUCH="true"*) wire signed [4:0] c20131,c21131,c22131,c23131,c24131,c25131,c26131,c27131;
(*DONT_TOUCH="true"*) wire signed [4:0] c20141,c21141,c22141,c23141,c24141,c25141,c26141,c27141;
(*DONT_TOUCH="true"*) wire signed [4:0] c20201,c21201,c22201,c23201,c24201,c25201,c26201,c27201;
(*DONT_TOUCH="true"*) wire signed [4:0] c20211,c21211,c22211,c23211,c24211,c25211,c26211,c27211;
(*DONT_TOUCH="true"*) wire signed [4:0] c20221,c21221,c22221,c23221,c24221,c25221,c26221,c27221;
(*DONT_TOUCH="true"*) wire signed [4:0] c20231,c21231,c22231,c23231,c24231,c25231,c26231,c27231;
(*DONT_TOUCH="true"*) wire signed [4:0] c20241,c21241,c22241,c23241,c24241,c25241,c26241,c27241;
(*DONT_TOUCH="true"*) wire signed [4:0] c20301,c21301,c22301,c23301,c24301,c25301,c26301,c27301;
(*DONT_TOUCH="true"*) wire signed [4:0] c20311,c21311,c22311,c23311,c24311,c25311,c26311,c27311;
(*DONT_TOUCH="true"*) wire signed [4:0] c20321,c21321,c22321,c23321,c24321,c25321,c26321,c27321;
(*DONT_TOUCH="true"*) wire signed [4:0] c20331,c21331,c22331,c23331,c24331,c25331,c26331,c27331;
(*DONT_TOUCH="true"*) wire signed [4:0] c20341,c21341,c22341,c23341,c24341,c25341,c26341,c27341;
(*DONT_TOUCH="true"*) wire signed [4:0] c20401,c21401,c22401,c23401,c24401,c25401,c26401,c27401;
(*DONT_TOUCH="true"*) wire signed [4:0] c20411,c21411,c22411,c23411,c24411,c25411,c26411,c27411;
(*DONT_TOUCH="true"*) wire signed [4:0] c20421,c21421,c22421,c23421,c24421,c25421,c26421,c27421;
(*DONT_TOUCH="true"*) wire signed [4:0] c20431,c21431,c22431,c23431,c24431,c25431,c26431,c27431;
(*DONT_TOUCH="true"*) wire signed [4:0] c20441,c21441,c22441,c23441,c24441,c25441,c26441,c27441;
(*DONT_TOUCH="true"*) wire signed [4:0] c20002,c21002,c22002,c23002,c24002,c25002,c26002,c27002;
(*DONT_TOUCH="true"*) wire signed [4:0] c20012,c21012,c22012,c23012,c24012,c25012,c26012,c27012;
(*DONT_TOUCH="true"*) wire signed [4:0] c20022,c21022,c22022,c23022,c24022,c25022,c26022,c27022;
(*DONT_TOUCH="true"*) wire signed [4:0] c20032,c21032,c22032,c23032,c24032,c25032,c26032,c27032;
(*DONT_TOUCH="true"*) wire signed [4:0] c20042,c21042,c22042,c23042,c24042,c25042,c26042,c27042;
(*DONT_TOUCH="true"*) wire signed [4:0] c20102,c21102,c22102,c23102,c24102,c25102,c26102,c27102;
(*DONT_TOUCH="true"*) wire signed [4:0] c20112,c21112,c22112,c23112,c24112,c25112,c26112,c27112;
(*DONT_TOUCH="true"*) wire signed [4:0] c20122,c21122,c22122,c23122,c24122,c25122,c26122,c27122;
(*DONT_TOUCH="true"*) wire signed [4:0] c20132,c21132,c22132,c23132,c24132,c25132,c26132,c27132;
(*DONT_TOUCH="true"*) wire signed [4:0] c20142,c21142,c22142,c23142,c24142,c25142,c26142,c27142;
(*DONT_TOUCH="true"*) wire signed [4:0] c20202,c21202,c22202,c23202,c24202,c25202,c26202,c27202;
(*DONT_TOUCH="true"*) wire signed [4:0] c20212,c21212,c22212,c23212,c24212,c25212,c26212,c27212;
(*DONT_TOUCH="true"*) wire signed [4:0] c20222,c21222,c22222,c23222,c24222,c25222,c26222,c27222;
(*DONT_TOUCH="true"*) wire signed [4:0] c20232,c21232,c22232,c23232,c24232,c25232,c26232,c27232;
(*DONT_TOUCH="true"*) wire signed [4:0] c20242,c21242,c22242,c23242,c24242,c25242,c26242,c27242;
(*DONT_TOUCH="true"*) wire signed [4:0] c20302,c21302,c22302,c23302,c24302,c25302,c26302,c27302;
(*DONT_TOUCH="true"*) wire signed [4:0] c20312,c21312,c22312,c23312,c24312,c25312,c26312,c27312;
(*DONT_TOUCH="true"*) wire signed [4:0] c20322,c21322,c22322,c23322,c24322,c25322,c26322,c27322;
(*DONT_TOUCH="true"*) wire signed [4:0] c20332,c21332,c22332,c23332,c24332,c25332,c26332,c27332;
(*DONT_TOUCH="true"*) wire signed [4:0] c20342,c21342,c22342,c23342,c24342,c25342,c26342,c27342;
(*DONT_TOUCH="true"*) wire signed [4:0] c20402,c21402,c22402,c23402,c24402,c25402,c26402,c27402;
(*DONT_TOUCH="true"*) wire signed [4:0] c20412,c21412,c22412,c23412,c24412,c25412,c26412,c27412;
(*DONT_TOUCH="true"*) wire signed [4:0] c20422,c21422,c22422,c23422,c24422,c25422,c26422,c27422;
(*DONT_TOUCH="true"*) wire signed [4:0] c20432,c21432,c22432,c23432,c24432,c25432,c26432,c27432;
(*DONT_TOUCH="true"*) wire signed [4:0] c20442,c21442,c22442,c23442,c24442,c25442,c26442,c27442;
(*DONT_TOUCH="true"*) wire signed [4:0] c20003,c21003,c22003,c23003,c24003,c25003,c26003,c27003;
(*DONT_TOUCH="true"*) wire signed [4:0] c20013,c21013,c22013,c23013,c24013,c25013,c26013,c27013;
(*DONT_TOUCH="true"*) wire signed [4:0] c20023,c21023,c22023,c23023,c24023,c25023,c26023,c27023;
(*DONT_TOUCH="true"*) wire signed [4:0] c20033,c21033,c22033,c23033,c24033,c25033,c26033,c27033;
(*DONT_TOUCH="true"*) wire signed [4:0] c20043,c21043,c22043,c23043,c24043,c25043,c26043,c27043;
(*DONT_TOUCH="true"*) wire signed [4:0] c20103,c21103,c22103,c23103,c24103,c25103,c26103,c27103;
(*DONT_TOUCH="true"*) wire signed [4:0] c20113,c21113,c22113,c23113,c24113,c25113,c26113,c27113;
(*DONT_TOUCH="true"*) wire signed [4:0] c20123,c21123,c22123,c23123,c24123,c25123,c26123,c27123;
(*DONT_TOUCH="true"*) wire signed [4:0] c20133,c21133,c22133,c23133,c24133,c25133,c26133,c27133;
(*DONT_TOUCH="true"*) wire signed [4:0] c20143,c21143,c22143,c23143,c24143,c25143,c26143,c27143;
(*DONT_TOUCH="true"*) wire signed [4:0] c20203,c21203,c22203,c23203,c24203,c25203,c26203,c27203;
(*DONT_TOUCH="true"*) wire signed [4:0] c20213,c21213,c22213,c23213,c24213,c25213,c26213,c27213;
(*DONT_TOUCH="true"*) wire signed [4:0] c20223,c21223,c22223,c23223,c24223,c25223,c26223,c27223;
(*DONT_TOUCH="true"*) wire signed [4:0] c20233,c21233,c22233,c23233,c24233,c25233,c26233,c27233;
(*DONT_TOUCH="true"*) wire signed [4:0] c20243,c21243,c22243,c23243,c24243,c25243,c26243,c27243;
(*DONT_TOUCH="true"*) wire signed [4:0] c20303,c21303,c22303,c23303,c24303,c25303,c26303,c27303;
(*DONT_TOUCH="true"*) wire signed [4:0] c20313,c21313,c22313,c23313,c24313,c25313,c26313,c27313;
(*DONT_TOUCH="true"*) wire signed [4:0] c20323,c21323,c22323,c23323,c24323,c25323,c26323,c27323;
(*DONT_TOUCH="true"*) wire signed [4:0] c20333,c21333,c22333,c23333,c24333,c25333,c26333,c27333;
(*DONT_TOUCH="true"*) wire signed [4:0] c20343,c21343,c22343,c23343,c24343,c25343,c26343,c27343;
(*DONT_TOUCH="true"*) wire signed [4:0] c20403,c21403,c22403,c23403,c24403,c25403,c26403,c27403;
(*DONT_TOUCH="true"*) wire signed [4:0] c20413,c21413,c22413,c23413,c24413,c25413,c26413,c27413;
(*DONT_TOUCH="true"*) wire signed [4:0] c20423,c21423,c22423,c23423,c24423,c25423,c26423,c27423;
(*DONT_TOUCH="true"*) wire signed [4:0] c20433,c21433,c22433,c23433,c24433,c25433,c26433,c27433;
(*DONT_TOUCH="true"*) wire signed [4:0] c20443,c21443,c22443,c23443,c24443,c25443,c26443,c27443;
(*DONT_TOUCH="true"*) wire signed [4:0] c20004,c21004,c22004,c23004,c24004,c25004,c26004,c27004;
(*DONT_TOUCH="true"*) wire signed [4:0] c20014,c21014,c22014,c23014,c24014,c25014,c26014,c27014;
(*DONT_TOUCH="true"*) wire signed [4:0] c20024,c21024,c22024,c23024,c24024,c25024,c26024,c27024;
(*DONT_TOUCH="true"*) wire signed [4:0] c20034,c21034,c22034,c23034,c24034,c25034,c26034,c27034;
(*DONT_TOUCH="true"*) wire signed [4:0] c20044,c21044,c22044,c23044,c24044,c25044,c26044,c27044;
(*DONT_TOUCH="true"*) wire signed [4:0] c20104,c21104,c22104,c23104,c24104,c25104,c26104,c27104;
(*DONT_TOUCH="true"*) wire signed [4:0] c20114,c21114,c22114,c23114,c24114,c25114,c26114,c27114;
(*DONT_TOUCH="true"*) wire signed [4:0] c20124,c21124,c22124,c23124,c24124,c25124,c26124,c27124;
(*DONT_TOUCH="true"*) wire signed [4:0] c20134,c21134,c22134,c23134,c24134,c25134,c26134,c27134;
(*DONT_TOUCH="true"*) wire signed [4:0] c20144,c21144,c22144,c23144,c24144,c25144,c26144,c27144;
(*DONT_TOUCH="true"*) wire signed [4:0] c20204,c21204,c22204,c23204,c24204,c25204,c26204,c27204;
(*DONT_TOUCH="true"*) wire signed [4:0] c20214,c21214,c22214,c23214,c24214,c25214,c26214,c27214;
(*DONT_TOUCH="true"*) wire signed [4:0] c20224,c21224,c22224,c23224,c24224,c25224,c26224,c27224;
(*DONT_TOUCH="true"*) wire signed [4:0] c20234,c21234,c22234,c23234,c24234,c25234,c26234,c27234;
(*DONT_TOUCH="true"*) wire signed [4:0] c20244,c21244,c22244,c23244,c24244,c25244,c26244,c27244;
(*DONT_TOUCH="true"*) wire signed [4:0] c20304,c21304,c22304,c23304,c24304,c25304,c26304,c27304;
(*DONT_TOUCH="true"*) wire signed [4:0] c20314,c21314,c22314,c23314,c24314,c25314,c26314,c27314;
(*DONT_TOUCH="true"*) wire signed [4:0] c20324,c21324,c22324,c23324,c24324,c25324,c26324,c27324;
(*DONT_TOUCH="true"*) wire signed [4:0] c20334,c21334,c22334,c23334,c24334,c25334,c26334,c27334;
(*DONT_TOUCH="true"*) wire signed [4:0] c20344,c21344,c22344,c23344,c24344,c25344,c26344,c27344;
(*DONT_TOUCH="true"*) wire signed [4:0] c20404,c21404,c22404,c23404,c24404,c25404,c26404,c27404;
(*DONT_TOUCH="true"*) wire signed [4:0] c20414,c21414,c22414,c23414,c24414,c25414,c26414,c27414;
(*DONT_TOUCH="true"*) wire signed [4:0] c20424,c21424,c22424,c23424,c24424,c25424,c26424,c27424;
(*DONT_TOUCH="true"*) wire signed [4:0] c20434,c21434,c22434,c23434,c24434,c25434,c26434,c27434;
(*DONT_TOUCH="true"*) wire signed [4:0] c20444,c21444,c22444,c23444,c24444,c25444,c26444,c27444;
(*DONT_TOUCH="true"*) wire signed [4:0] c20005,c21005,c22005,c23005,c24005,c25005,c26005,c27005;
(*DONT_TOUCH="true"*) wire signed [4:0] c20015,c21015,c22015,c23015,c24015,c25015,c26015,c27015;
(*DONT_TOUCH="true"*) wire signed [4:0] c20025,c21025,c22025,c23025,c24025,c25025,c26025,c27025;
(*DONT_TOUCH="true"*) wire signed [4:0] c20035,c21035,c22035,c23035,c24035,c25035,c26035,c27035;
(*DONT_TOUCH="true"*) wire signed [4:0] c20045,c21045,c22045,c23045,c24045,c25045,c26045,c27045;
(*DONT_TOUCH="true"*) wire signed [4:0] c20105,c21105,c22105,c23105,c24105,c25105,c26105,c27105;
(*DONT_TOUCH="true"*) wire signed [4:0] c20115,c21115,c22115,c23115,c24115,c25115,c26115,c27115;
(*DONT_TOUCH="true"*) wire signed [4:0] c20125,c21125,c22125,c23125,c24125,c25125,c26125,c27125;
(*DONT_TOUCH="true"*) wire signed [4:0] c20135,c21135,c22135,c23135,c24135,c25135,c26135,c27135;
(*DONT_TOUCH="true"*) wire signed [4:0] c20145,c21145,c22145,c23145,c24145,c25145,c26145,c27145;
(*DONT_TOUCH="true"*) wire signed [4:0] c20205,c21205,c22205,c23205,c24205,c25205,c26205,c27205;
(*DONT_TOUCH="true"*) wire signed [4:0] c20215,c21215,c22215,c23215,c24215,c25215,c26215,c27215;
(*DONT_TOUCH="true"*) wire signed [4:0] c20225,c21225,c22225,c23225,c24225,c25225,c26225,c27225;
(*DONT_TOUCH="true"*) wire signed [4:0] c20235,c21235,c22235,c23235,c24235,c25235,c26235,c27235;
(*DONT_TOUCH="true"*) wire signed [4:0] c20245,c21245,c22245,c23245,c24245,c25245,c26245,c27245;
(*DONT_TOUCH="true"*) wire signed [4:0] c20305,c21305,c22305,c23305,c24305,c25305,c26305,c27305;
(*DONT_TOUCH="true"*) wire signed [4:0] c20315,c21315,c22315,c23315,c24315,c25315,c26315,c27315;
(*DONT_TOUCH="true"*) wire signed [4:0] c20325,c21325,c22325,c23325,c24325,c25325,c26325,c27325;
(*DONT_TOUCH="true"*) wire signed [4:0] c20335,c21335,c22335,c23335,c24335,c25335,c26335,c27335;
(*DONT_TOUCH="true"*) wire signed [4:0] c20345,c21345,c22345,c23345,c24345,c25345,c26345,c27345;
(*DONT_TOUCH="true"*) wire signed [4:0] c20405,c21405,c22405,c23405,c24405,c25405,c26405,c27405;
(*DONT_TOUCH="true"*) wire signed [4:0] c20415,c21415,c22415,c23415,c24415,c25415,c26415,c27415;
(*DONT_TOUCH="true"*) wire signed [4:0] c20425,c21425,c22425,c23425,c24425,c25425,c26425,c27425;
(*DONT_TOUCH="true"*) wire signed [4:0] c20435,c21435,c22435,c23435,c24435,c25435,c26435,c27435;
(*DONT_TOUCH="true"*) wire signed [4:0] c20445,c21445,c22445,c23445,c24445,c25445,c26445,c27445;
(*DONT_TOUCH="true"*) wire signed [4:0] c20006,c21006,c22006,c23006,c24006,c25006,c26006,c27006;
(*DONT_TOUCH="true"*) wire signed [4:0] c20016,c21016,c22016,c23016,c24016,c25016,c26016,c27016;
(*DONT_TOUCH="true"*) wire signed [4:0] c20026,c21026,c22026,c23026,c24026,c25026,c26026,c27026;
(*DONT_TOUCH="true"*) wire signed [4:0] c20036,c21036,c22036,c23036,c24036,c25036,c26036,c27036;
(*DONT_TOUCH="true"*) wire signed [4:0] c20046,c21046,c22046,c23046,c24046,c25046,c26046,c27046;
(*DONT_TOUCH="true"*) wire signed [4:0] c20106,c21106,c22106,c23106,c24106,c25106,c26106,c27106;
(*DONT_TOUCH="true"*) wire signed [4:0] c20116,c21116,c22116,c23116,c24116,c25116,c26116,c27116;
(*DONT_TOUCH="true"*) wire signed [4:0] c20126,c21126,c22126,c23126,c24126,c25126,c26126,c27126;
(*DONT_TOUCH="true"*) wire signed [4:0] c20136,c21136,c22136,c23136,c24136,c25136,c26136,c27136;
(*DONT_TOUCH="true"*) wire signed [4:0] c20146,c21146,c22146,c23146,c24146,c25146,c26146,c27146;
(*DONT_TOUCH="true"*) wire signed [4:0] c20206,c21206,c22206,c23206,c24206,c25206,c26206,c27206;
(*DONT_TOUCH="true"*) wire signed [4:0] c20216,c21216,c22216,c23216,c24216,c25216,c26216,c27216;
(*DONT_TOUCH="true"*) wire signed [4:0] c20226,c21226,c22226,c23226,c24226,c25226,c26226,c27226;
(*DONT_TOUCH="true"*) wire signed [4:0] c20236,c21236,c22236,c23236,c24236,c25236,c26236,c27236;
(*DONT_TOUCH="true"*) wire signed [4:0] c20246,c21246,c22246,c23246,c24246,c25246,c26246,c27246;
(*DONT_TOUCH="true"*) wire signed [4:0] c20306,c21306,c22306,c23306,c24306,c25306,c26306,c27306;
(*DONT_TOUCH="true"*) wire signed [4:0] c20316,c21316,c22316,c23316,c24316,c25316,c26316,c27316;
(*DONT_TOUCH="true"*) wire signed [4:0] c20326,c21326,c22326,c23326,c24326,c25326,c26326,c27326;
(*DONT_TOUCH="true"*) wire signed [4:0] c20336,c21336,c22336,c23336,c24336,c25336,c26336,c27336;
(*DONT_TOUCH="true"*) wire signed [4:0] c20346,c21346,c22346,c23346,c24346,c25346,c26346,c27346;
(*DONT_TOUCH="true"*) wire signed [4:0] c20406,c21406,c22406,c23406,c24406,c25406,c26406,c27406;
(*DONT_TOUCH="true"*) wire signed [4:0] c20416,c21416,c22416,c23416,c24416,c25416,c26416,c27416;
(*DONT_TOUCH="true"*) wire signed [4:0] c20426,c21426,c22426,c23426,c24426,c25426,c26426,c27426;
(*DONT_TOUCH="true"*) wire signed [4:0] c20436,c21436,c22436,c23436,c24436,c25436,c26436,c27436;
(*DONT_TOUCH="true"*) wire signed [4:0] c20446,c21446,c22446,c23446,c24446,c25446,c26446,c27446;
(*DONT_TOUCH="true"*) wire signed [4:0] c20007,c21007,c22007,c23007,c24007,c25007,c26007,c27007;
(*DONT_TOUCH="true"*) wire signed [4:0] c20017,c21017,c22017,c23017,c24017,c25017,c26017,c27017;
(*DONT_TOUCH="true"*) wire signed [4:0] c20027,c21027,c22027,c23027,c24027,c25027,c26027,c27027;
(*DONT_TOUCH="true"*) wire signed [4:0] c20037,c21037,c22037,c23037,c24037,c25037,c26037,c27037;
(*DONT_TOUCH="true"*) wire signed [4:0] c20047,c21047,c22047,c23047,c24047,c25047,c26047,c27047;
(*DONT_TOUCH="true"*) wire signed [4:0] c20107,c21107,c22107,c23107,c24107,c25107,c26107,c27107;
(*DONT_TOUCH="true"*) wire signed [4:0] c20117,c21117,c22117,c23117,c24117,c25117,c26117,c27117;
(*DONT_TOUCH="true"*) wire signed [4:0] c20127,c21127,c22127,c23127,c24127,c25127,c26127,c27127;
(*DONT_TOUCH="true"*) wire signed [4:0] c20137,c21137,c22137,c23137,c24137,c25137,c26137,c27137;
(*DONT_TOUCH="true"*) wire signed [4:0] c20147,c21147,c22147,c23147,c24147,c25147,c26147,c27147;
(*DONT_TOUCH="true"*) wire signed [4:0] c20207,c21207,c22207,c23207,c24207,c25207,c26207,c27207;
(*DONT_TOUCH="true"*) wire signed [4:0] c20217,c21217,c22217,c23217,c24217,c25217,c26217,c27217;
(*DONT_TOUCH="true"*) wire signed [4:0] c20227,c21227,c22227,c23227,c24227,c25227,c26227,c27227;
(*DONT_TOUCH="true"*) wire signed [4:0] c20237,c21237,c22237,c23237,c24237,c25237,c26237,c27237;
(*DONT_TOUCH="true"*) wire signed [4:0] c20247,c21247,c22247,c23247,c24247,c25247,c26247,c27247;
(*DONT_TOUCH="true"*) wire signed [4:0] c20307,c21307,c22307,c23307,c24307,c25307,c26307,c27307;
(*DONT_TOUCH="true"*) wire signed [4:0] c20317,c21317,c22317,c23317,c24317,c25317,c26317,c27317;
(*DONT_TOUCH="true"*) wire signed [4:0] c20327,c21327,c22327,c23327,c24327,c25327,c26327,c27327;
(*DONT_TOUCH="true"*) wire signed [4:0] c20337,c21337,c22337,c23337,c24337,c25337,c26337,c27337;
(*DONT_TOUCH="true"*) wire signed [4:0] c20347,c21347,c22347,c23347,c24347,c25347,c26347,c27347;
(*DONT_TOUCH="true"*) wire signed [4:0] c20407,c21407,c22407,c23407,c24407,c25407,c26407,c27407;
(*DONT_TOUCH="true"*) wire signed [4:0] c20417,c21417,c22417,c23417,c24417,c25417,c26417,c27417;
(*DONT_TOUCH="true"*) wire signed [4:0] c20427,c21427,c22427,c23427,c24427,c25427,c26427,c27427;
(*DONT_TOUCH="true"*) wire signed [4:0] c20437,c21437,c22437,c23437,c24437,c25437,c26437,c27437;
(*DONT_TOUCH="true"*) wire signed [4:0] c20447,c21447,c22447,c23447,c24447,c25447,c26447,c27447;
(*DONT_TOUCH="true"*) wire signed [4:0] c20008,c21008,c22008,c23008,c24008,c25008,c26008,c27008;
(*DONT_TOUCH="true"*) wire signed [4:0] c20018,c21018,c22018,c23018,c24018,c25018,c26018,c27018;
(*DONT_TOUCH="true"*) wire signed [4:0] c20028,c21028,c22028,c23028,c24028,c25028,c26028,c27028;
(*DONT_TOUCH="true"*) wire signed [4:0] c20038,c21038,c22038,c23038,c24038,c25038,c26038,c27038;
(*DONT_TOUCH="true"*) wire signed [4:0] c20048,c21048,c22048,c23048,c24048,c25048,c26048,c27048;
(*DONT_TOUCH="true"*) wire signed [4:0] c20108,c21108,c22108,c23108,c24108,c25108,c26108,c27108;
(*DONT_TOUCH="true"*) wire signed [4:0] c20118,c21118,c22118,c23118,c24118,c25118,c26118,c27118;
(*DONT_TOUCH="true"*) wire signed [4:0] c20128,c21128,c22128,c23128,c24128,c25128,c26128,c27128;
(*DONT_TOUCH="true"*) wire signed [4:0] c20138,c21138,c22138,c23138,c24138,c25138,c26138,c27138;
(*DONT_TOUCH="true"*) wire signed [4:0] c20148,c21148,c22148,c23148,c24148,c25148,c26148,c27148;
(*DONT_TOUCH="true"*) wire signed [4:0] c20208,c21208,c22208,c23208,c24208,c25208,c26208,c27208;
(*DONT_TOUCH="true"*) wire signed [4:0] c20218,c21218,c22218,c23218,c24218,c25218,c26218,c27218;
(*DONT_TOUCH="true"*) wire signed [4:0] c20228,c21228,c22228,c23228,c24228,c25228,c26228,c27228;
(*DONT_TOUCH="true"*) wire signed [4:0] c20238,c21238,c22238,c23238,c24238,c25238,c26238,c27238;
(*DONT_TOUCH="true"*) wire signed [4:0] c20248,c21248,c22248,c23248,c24248,c25248,c26248,c27248;
(*DONT_TOUCH="true"*) wire signed [4:0] c20308,c21308,c22308,c23308,c24308,c25308,c26308,c27308;
(*DONT_TOUCH="true"*) wire signed [4:0] c20318,c21318,c22318,c23318,c24318,c25318,c26318,c27318;
(*DONT_TOUCH="true"*) wire signed [4:0] c20328,c21328,c22328,c23328,c24328,c25328,c26328,c27328;
(*DONT_TOUCH="true"*) wire signed [4:0] c20338,c21338,c22338,c23338,c24338,c25338,c26338,c27338;
(*DONT_TOUCH="true"*) wire signed [4:0] c20348,c21348,c22348,c23348,c24348,c25348,c26348,c27348;
(*DONT_TOUCH="true"*) wire signed [4:0] c20408,c21408,c22408,c23408,c24408,c25408,c26408,c27408;
(*DONT_TOUCH="true"*) wire signed [4:0] c20418,c21418,c22418,c23418,c24418,c25418,c26418,c27418;
(*DONT_TOUCH="true"*) wire signed [4:0] c20428,c21428,c22428,c23428,c24428,c25428,c26428,c27428;
(*DONT_TOUCH="true"*) wire signed [4:0] c20438,c21438,c22438,c23438,c24438,c25438,c26438,c27438;
(*DONT_TOUCH="true"*) wire signed [4:0] c20448,c21448,c22448,c23448,c24448,c25448,c26448,c27448;
(*DONT_TOUCH="true"*) wire signed [4:0] c20009,c21009,c22009,c23009,c24009,c25009,c26009,c27009;
(*DONT_TOUCH="true"*) wire signed [4:0] c20019,c21019,c22019,c23019,c24019,c25019,c26019,c27019;
(*DONT_TOUCH="true"*) wire signed [4:0] c20029,c21029,c22029,c23029,c24029,c25029,c26029,c27029;
(*DONT_TOUCH="true"*) wire signed [4:0] c20039,c21039,c22039,c23039,c24039,c25039,c26039,c27039;
(*DONT_TOUCH="true"*) wire signed [4:0] c20049,c21049,c22049,c23049,c24049,c25049,c26049,c27049;
(*DONT_TOUCH="true"*) wire signed [4:0] c20109,c21109,c22109,c23109,c24109,c25109,c26109,c27109;
(*DONT_TOUCH="true"*) wire signed [4:0] c20119,c21119,c22119,c23119,c24119,c25119,c26119,c27119;
(*DONT_TOUCH="true"*) wire signed [4:0] c20129,c21129,c22129,c23129,c24129,c25129,c26129,c27129;
(*DONT_TOUCH="true"*) wire signed [4:0] c20139,c21139,c22139,c23139,c24139,c25139,c26139,c27139;
(*DONT_TOUCH="true"*) wire signed [4:0] c20149,c21149,c22149,c23149,c24149,c25149,c26149,c27149;
(*DONT_TOUCH="true"*) wire signed [4:0] c20209,c21209,c22209,c23209,c24209,c25209,c26209,c27209;
(*DONT_TOUCH="true"*) wire signed [4:0] c20219,c21219,c22219,c23219,c24219,c25219,c26219,c27219;
(*DONT_TOUCH="true"*) wire signed [4:0] c20229,c21229,c22229,c23229,c24229,c25229,c26229,c27229;
(*DONT_TOUCH="true"*) wire signed [4:0] c20239,c21239,c22239,c23239,c24239,c25239,c26239,c27239;
(*DONT_TOUCH="true"*) wire signed [4:0] c20249,c21249,c22249,c23249,c24249,c25249,c26249,c27249;
(*DONT_TOUCH="true"*) wire signed [4:0] c20309,c21309,c22309,c23309,c24309,c25309,c26309,c27309;
(*DONT_TOUCH="true"*) wire signed [4:0] c20319,c21319,c22319,c23319,c24319,c25319,c26319,c27319;
(*DONT_TOUCH="true"*) wire signed [4:0] c20329,c21329,c22329,c23329,c24329,c25329,c26329,c27329;
(*DONT_TOUCH="true"*) wire signed [4:0] c20339,c21339,c22339,c23339,c24339,c25339,c26339,c27339;
(*DONT_TOUCH="true"*) wire signed [4:0] c20349,c21349,c22349,c23349,c24349,c25349,c26349,c27349;
(*DONT_TOUCH="true"*) wire signed [4:0] c20409,c21409,c22409,c23409,c24409,c25409,c26409,c27409;
(*DONT_TOUCH="true"*) wire signed [4:0] c20419,c21419,c22419,c23419,c24419,c25419,c26419,c27419;
(*DONT_TOUCH="true"*) wire signed [4:0] c20429,c21429,c22429,c23429,c24429,c25429,c26429,c27429;
(*DONT_TOUCH="true"*) wire signed [4:0] c20439,c21439,c22439,c23439,c24439,c25439,c26439,c27439;
(*DONT_TOUCH="true"*) wire signed [4:0] c20449,c21449,c22449,c23449,c24449,c25449,c26449,c27449;
(*DONT_TOUCH="true"*) wire signed [4:0] c2000A,c2100A,c2200A,c2300A,c2400A,c2500A,c2600A,c2700A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2001A,c2101A,c2201A,c2301A,c2401A,c2501A,c2601A,c2701A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2002A,c2102A,c2202A,c2302A,c2402A,c2502A,c2602A,c2702A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2003A,c2103A,c2203A,c2303A,c2403A,c2503A,c2603A,c2703A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2004A,c2104A,c2204A,c2304A,c2404A,c2504A,c2604A,c2704A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2010A,c2110A,c2210A,c2310A,c2410A,c2510A,c2610A,c2710A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2011A,c2111A,c2211A,c2311A,c2411A,c2511A,c2611A,c2711A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2012A,c2112A,c2212A,c2312A,c2412A,c2512A,c2612A,c2712A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2013A,c2113A,c2213A,c2313A,c2413A,c2513A,c2613A,c2713A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2014A,c2114A,c2214A,c2314A,c2414A,c2514A,c2614A,c2714A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2020A,c2120A,c2220A,c2320A,c2420A,c2520A,c2620A,c2720A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2021A,c2121A,c2221A,c2321A,c2421A,c2521A,c2621A,c2721A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2022A,c2122A,c2222A,c2322A,c2422A,c2522A,c2622A,c2722A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2023A,c2123A,c2223A,c2323A,c2423A,c2523A,c2623A,c2723A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2024A,c2124A,c2224A,c2324A,c2424A,c2524A,c2624A,c2724A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2030A,c2130A,c2230A,c2330A,c2430A,c2530A,c2630A,c2730A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2031A,c2131A,c2231A,c2331A,c2431A,c2531A,c2631A,c2731A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2032A,c2132A,c2232A,c2332A,c2432A,c2532A,c2632A,c2732A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2033A,c2133A,c2233A,c2333A,c2433A,c2533A,c2633A,c2733A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2034A,c2134A,c2234A,c2334A,c2434A,c2534A,c2634A,c2734A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2040A,c2140A,c2240A,c2340A,c2440A,c2540A,c2640A,c2740A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2041A,c2141A,c2241A,c2341A,c2441A,c2541A,c2641A,c2741A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2042A,c2142A,c2242A,c2342A,c2442A,c2542A,c2642A,c2742A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2043A,c2143A,c2243A,c2343A,c2443A,c2543A,c2643A,c2743A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2044A,c2144A,c2244A,c2344A,c2444A,c2544A,c2644A,c2744A;
(*DONT_TOUCH="true"*) wire signed [4:0] c2000B,c2100B,c2200B,c2300B,c2400B,c2500B,c2600B,c2700B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2001B,c2101B,c2201B,c2301B,c2401B,c2501B,c2601B,c2701B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2002B,c2102B,c2202B,c2302B,c2402B,c2502B,c2602B,c2702B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2003B,c2103B,c2203B,c2303B,c2403B,c2503B,c2603B,c2703B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2004B,c2104B,c2204B,c2304B,c2404B,c2504B,c2604B,c2704B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2010B,c2110B,c2210B,c2310B,c2410B,c2510B,c2610B,c2710B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2011B,c2111B,c2211B,c2311B,c2411B,c2511B,c2611B,c2711B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2012B,c2112B,c2212B,c2312B,c2412B,c2512B,c2612B,c2712B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2013B,c2113B,c2213B,c2313B,c2413B,c2513B,c2613B,c2713B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2014B,c2114B,c2214B,c2314B,c2414B,c2514B,c2614B,c2714B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2020B,c2120B,c2220B,c2320B,c2420B,c2520B,c2620B,c2720B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2021B,c2121B,c2221B,c2321B,c2421B,c2521B,c2621B,c2721B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2022B,c2122B,c2222B,c2322B,c2422B,c2522B,c2622B,c2722B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2023B,c2123B,c2223B,c2323B,c2423B,c2523B,c2623B,c2723B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2024B,c2124B,c2224B,c2324B,c2424B,c2524B,c2624B,c2724B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2030B,c2130B,c2230B,c2330B,c2430B,c2530B,c2630B,c2730B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2031B,c2131B,c2231B,c2331B,c2431B,c2531B,c2631B,c2731B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2032B,c2132B,c2232B,c2332B,c2432B,c2532B,c2632B,c2732B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2033B,c2133B,c2233B,c2333B,c2433B,c2533B,c2633B,c2733B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2034B,c2134B,c2234B,c2334B,c2434B,c2534B,c2634B,c2734B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2040B,c2140B,c2240B,c2340B,c2440B,c2540B,c2640B,c2740B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2041B,c2141B,c2241B,c2341B,c2441B,c2541B,c2641B,c2741B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2042B,c2142B,c2242B,c2342B,c2442B,c2542B,c2642B,c2742B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2043B,c2143B,c2243B,c2343B,c2443B,c2543B,c2643B,c2743B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2044B,c2144B,c2244B,c2344B,c2444B,c2544B,c2644B,c2744B;
(*DONT_TOUCH="true"*) wire signed [4:0] c2000C,c2100C,c2200C,c2300C,c2400C,c2500C,c2600C,c2700C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2001C,c2101C,c2201C,c2301C,c2401C,c2501C,c2601C,c2701C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2002C,c2102C,c2202C,c2302C,c2402C,c2502C,c2602C,c2702C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2003C,c2103C,c2203C,c2303C,c2403C,c2503C,c2603C,c2703C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2004C,c2104C,c2204C,c2304C,c2404C,c2504C,c2604C,c2704C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2010C,c2110C,c2210C,c2310C,c2410C,c2510C,c2610C,c2710C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2011C,c2111C,c2211C,c2311C,c2411C,c2511C,c2611C,c2711C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2012C,c2112C,c2212C,c2312C,c2412C,c2512C,c2612C,c2712C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2013C,c2113C,c2213C,c2313C,c2413C,c2513C,c2613C,c2713C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2014C,c2114C,c2214C,c2314C,c2414C,c2514C,c2614C,c2714C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2020C,c2120C,c2220C,c2320C,c2420C,c2520C,c2620C,c2720C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2021C,c2121C,c2221C,c2321C,c2421C,c2521C,c2621C,c2721C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2022C,c2122C,c2222C,c2322C,c2422C,c2522C,c2622C,c2722C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2023C,c2123C,c2223C,c2323C,c2423C,c2523C,c2623C,c2723C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2024C,c2124C,c2224C,c2324C,c2424C,c2524C,c2624C,c2724C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2030C,c2130C,c2230C,c2330C,c2430C,c2530C,c2630C,c2730C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2031C,c2131C,c2231C,c2331C,c2431C,c2531C,c2631C,c2731C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2032C,c2132C,c2232C,c2332C,c2432C,c2532C,c2632C,c2732C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2033C,c2133C,c2233C,c2333C,c2433C,c2533C,c2633C,c2733C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2034C,c2134C,c2234C,c2334C,c2434C,c2534C,c2634C,c2734C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2040C,c2140C,c2240C,c2340C,c2440C,c2540C,c2640C,c2740C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2041C,c2141C,c2241C,c2341C,c2441C,c2541C,c2641C,c2741C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2042C,c2142C,c2242C,c2342C,c2442C,c2542C,c2642C,c2742C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2043C,c2143C,c2243C,c2343C,c2443C,c2543C,c2643C,c2743C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2044C,c2144C,c2244C,c2344C,c2444C,c2544C,c2644C,c2744C;
(*DONT_TOUCH="true"*) wire signed [4:0] c2000D,c2100D,c2200D,c2300D,c2400D,c2500D,c2600D,c2700D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2001D,c2101D,c2201D,c2301D,c2401D,c2501D,c2601D,c2701D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2002D,c2102D,c2202D,c2302D,c2402D,c2502D,c2602D,c2702D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2003D,c2103D,c2203D,c2303D,c2403D,c2503D,c2603D,c2703D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2004D,c2104D,c2204D,c2304D,c2404D,c2504D,c2604D,c2704D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2010D,c2110D,c2210D,c2310D,c2410D,c2510D,c2610D,c2710D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2011D,c2111D,c2211D,c2311D,c2411D,c2511D,c2611D,c2711D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2012D,c2112D,c2212D,c2312D,c2412D,c2512D,c2612D,c2712D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2013D,c2113D,c2213D,c2313D,c2413D,c2513D,c2613D,c2713D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2014D,c2114D,c2214D,c2314D,c2414D,c2514D,c2614D,c2714D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2020D,c2120D,c2220D,c2320D,c2420D,c2520D,c2620D,c2720D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2021D,c2121D,c2221D,c2321D,c2421D,c2521D,c2621D,c2721D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2022D,c2122D,c2222D,c2322D,c2422D,c2522D,c2622D,c2722D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2023D,c2123D,c2223D,c2323D,c2423D,c2523D,c2623D,c2723D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2024D,c2124D,c2224D,c2324D,c2424D,c2524D,c2624D,c2724D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2030D,c2130D,c2230D,c2330D,c2430D,c2530D,c2630D,c2730D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2031D,c2131D,c2231D,c2331D,c2431D,c2531D,c2631D,c2731D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2032D,c2132D,c2232D,c2332D,c2432D,c2532D,c2632D,c2732D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2033D,c2133D,c2233D,c2333D,c2433D,c2533D,c2633D,c2733D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2034D,c2134D,c2234D,c2334D,c2434D,c2534D,c2634D,c2734D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2040D,c2140D,c2240D,c2340D,c2440D,c2540D,c2640D,c2740D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2041D,c2141D,c2241D,c2341D,c2441D,c2541D,c2641D,c2741D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2042D,c2142D,c2242D,c2342D,c2442D,c2542D,c2642D,c2742D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2043D,c2143D,c2243D,c2343D,c2443D,c2543D,c2643D,c2743D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2044D,c2144D,c2244D,c2344D,c2444D,c2544D,c2644D,c2744D;
(*DONT_TOUCH="true"*) wire signed [4:0] c2000E,c2100E,c2200E,c2300E,c2400E,c2500E,c2600E,c2700E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2001E,c2101E,c2201E,c2301E,c2401E,c2501E,c2601E,c2701E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2002E,c2102E,c2202E,c2302E,c2402E,c2502E,c2602E,c2702E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2003E,c2103E,c2203E,c2303E,c2403E,c2503E,c2603E,c2703E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2004E,c2104E,c2204E,c2304E,c2404E,c2504E,c2604E,c2704E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2010E,c2110E,c2210E,c2310E,c2410E,c2510E,c2610E,c2710E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2011E,c2111E,c2211E,c2311E,c2411E,c2511E,c2611E,c2711E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2012E,c2112E,c2212E,c2312E,c2412E,c2512E,c2612E,c2712E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2013E,c2113E,c2213E,c2313E,c2413E,c2513E,c2613E,c2713E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2014E,c2114E,c2214E,c2314E,c2414E,c2514E,c2614E,c2714E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2020E,c2120E,c2220E,c2320E,c2420E,c2520E,c2620E,c2720E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2021E,c2121E,c2221E,c2321E,c2421E,c2521E,c2621E,c2721E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2022E,c2122E,c2222E,c2322E,c2422E,c2522E,c2622E,c2722E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2023E,c2123E,c2223E,c2323E,c2423E,c2523E,c2623E,c2723E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2024E,c2124E,c2224E,c2324E,c2424E,c2524E,c2624E,c2724E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2030E,c2130E,c2230E,c2330E,c2430E,c2530E,c2630E,c2730E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2031E,c2131E,c2231E,c2331E,c2431E,c2531E,c2631E,c2731E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2032E,c2132E,c2232E,c2332E,c2432E,c2532E,c2632E,c2732E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2033E,c2133E,c2233E,c2333E,c2433E,c2533E,c2633E,c2733E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2034E,c2134E,c2234E,c2334E,c2434E,c2534E,c2634E,c2734E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2040E,c2140E,c2240E,c2340E,c2440E,c2540E,c2640E,c2740E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2041E,c2141E,c2241E,c2341E,c2441E,c2541E,c2641E,c2741E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2042E,c2142E,c2242E,c2342E,c2442E,c2542E,c2642E,c2742E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2043E,c2143E,c2243E,c2343E,c2443E,c2543E,c2643E,c2743E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2044E,c2144E,c2244E,c2344E,c2444E,c2544E,c2644E,c2744E;
(*DONT_TOUCH="true"*) wire signed [4:0] c2000F,c2100F,c2200F,c2300F,c2400F,c2500F,c2600F,c2700F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2001F,c2101F,c2201F,c2301F,c2401F,c2501F,c2601F,c2701F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2002F,c2102F,c2202F,c2302F,c2402F,c2502F,c2602F,c2702F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2003F,c2103F,c2203F,c2303F,c2403F,c2503F,c2603F,c2703F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2004F,c2104F,c2204F,c2304F,c2404F,c2504F,c2604F,c2704F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2010F,c2110F,c2210F,c2310F,c2410F,c2510F,c2610F,c2710F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2011F,c2111F,c2211F,c2311F,c2411F,c2511F,c2611F,c2711F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2012F,c2112F,c2212F,c2312F,c2412F,c2512F,c2612F,c2712F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2013F,c2113F,c2213F,c2313F,c2413F,c2513F,c2613F,c2713F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2014F,c2114F,c2214F,c2314F,c2414F,c2514F,c2614F,c2714F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2020F,c2120F,c2220F,c2320F,c2420F,c2520F,c2620F,c2720F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2021F,c2121F,c2221F,c2321F,c2421F,c2521F,c2621F,c2721F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2022F,c2122F,c2222F,c2322F,c2422F,c2522F,c2622F,c2722F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2023F,c2123F,c2223F,c2323F,c2423F,c2523F,c2623F,c2723F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2024F,c2124F,c2224F,c2324F,c2424F,c2524F,c2624F,c2724F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2030F,c2130F,c2230F,c2330F,c2430F,c2530F,c2630F,c2730F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2031F,c2131F,c2231F,c2331F,c2431F,c2531F,c2631F,c2731F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2032F,c2132F,c2232F,c2332F,c2432F,c2532F,c2632F,c2732F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2033F,c2133F,c2233F,c2333F,c2433F,c2533F,c2633F,c2733F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2034F,c2134F,c2234F,c2334F,c2434F,c2534F,c2634F,c2734F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2040F,c2140F,c2240F,c2340F,c2440F,c2540F,c2640F,c2740F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2041F,c2141F,c2241F,c2341F,c2441F,c2541F,c2641F,c2741F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2042F,c2142F,c2242F,c2342F,c2442F,c2542F,c2642F,c2742F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2043F,c2143F,c2243F,c2343F,c2443F,c2543F,c2643F,c2743F;
(*DONT_TOUCH="true"*) wire signed [4:0] c2044F,c2144F,c2244F,c2344F,c2444F,c2544F,c2644F,c2744F;
(*DONT_TOUCH="true"*) wire signed [7:0] C2000;
(*DONT_TOUCH="true"*) wire A2000;
(*DONT_TOUCH="true"*) wire signed [7:0] C2010;
(*DONT_TOUCH="true"*) wire A2010;
(*DONT_TOUCH="true"*) wire signed [7:0] C2020;
(*DONT_TOUCH="true"*) wire A2020;
(*DONT_TOUCH="true"*) wire signed [7:0] C2030;
(*DONT_TOUCH="true"*) wire A2030;
(*DONT_TOUCH="true"*) wire signed [7:0] C2040;
(*DONT_TOUCH="true"*) wire A2040;
(*DONT_TOUCH="true"*) wire signed [7:0] C2100;
(*DONT_TOUCH="true"*) wire A2100;
(*DONT_TOUCH="true"*) wire signed [7:0] C2110;
(*DONT_TOUCH="true"*) wire A2110;
(*DONT_TOUCH="true"*) wire signed [7:0] C2120;
(*DONT_TOUCH="true"*) wire A2120;
(*DONT_TOUCH="true"*) wire signed [7:0] C2130;
(*DONT_TOUCH="true"*) wire A2130;
(*DONT_TOUCH="true"*) wire signed [7:0] C2140;
(*DONT_TOUCH="true"*) wire A2140;
(*DONT_TOUCH="true"*) wire signed [7:0] C2200;
(*DONT_TOUCH="true"*) wire A2200;
(*DONT_TOUCH="true"*) wire signed [7:0] C2210;
(*DONT_TOUCH="true"*) wire A2210;
(*DONT_TOUCH="true"*) wire signed [7:0] C2220;
(*DONT_TOUCH="true"*) wire A2220;
(*DONT_TOUCH="true"*) wire signed [7:0] C2230;
(*DONT_TOUCH="true"*) wire A2230;
(*DONT_TOUCH="true"*) wire signed [7:0] C2240;
(*DONT_TOUCH="true"*) wire A2240;
(*DONT_TOUCH="true"*) wire signed [7:0] C2300;
(*DONT_TOUCH="true"*) wire A2300;
(*DONT_TOUCH="true"*) wire signed [7:0] C2310;
(*DONT_TOUCH="true"*) wire A2310;
(*DONT_TOUCH="true"*) wire signed [7:0] C2320;
(*DONT_TOUCH="true"*) wire A2320;
(*DONT_TOUCH="true"*) wire signed [7:0] C2330;
(*DONT_TOUCH="true"*) wire A2330;
(*DONT_TOUCH="true"*) wire signed [7:0] C2340;
(*DONT_TOUCH="true"*) wire A2340;
(*DONT_TOUCH="true"*) wire signed [7:0] C2400;
(*DONT_TOUCH="true"*) wire A2400;
(*DONT_TOUCH="true"*) wire signed [7:0] C2410;
(*DONT_TOUCH="true"*) wire A2410;
(*DONT_TOUCH="true"*) wire signed [7:0] C2420;
(*DONT_TOUCH="true"*) wire A2420;
(*DONT_TOUCH="true"*) wire signed [7:0] C2430;
(*DONT_TOUCH="true"*) wire A2430;
(*DONT_TOUCH="true"*) wire signed [7:0] C2440;
(*DONT_TOUCH="true"*) wire A2440;
(*DONT_TOUCH="true"*) wire signed [7:0] C2001;
(*DONT_TOUCH="true"*) wire A2001;
(*DONT_TOUCH="true"*) wire signed [7:0] C2011;
(*DONT_TOUCH="true"*) wire A2011;
(*DONT_TOUCH="true"*) wire signed [7:0] C2021;
(*DONT_TOUCH="true"*) wire A2021;
(*DONT_TOUCH="true"*) wire signed [7:0] C2031;
(*DONT_TOUCH="true"*) wire A2031;
(*DONT_TOUCH="true"*) wire signed [7:0] C2041;
(*DONT_TOUCH="true"*) wire A2041;
(*DONT_TOUCH="true"*) wire signed [7:0] C2101;
(*DONT_TOUCH="true"*) wire A2101;
(*DONT_TOUCH="true"*) wire signed [7:0] C2111;
(*DONT_TOUCH="true"*) wire A2111;
(*DONT_TOUCH="true"*) wire signed [7:0] C2121;
(*DONT_TOUCH="true"*) wire A2121;
(*DONT_TOUCH="true"*) wire signed [7:0] C2131;
(*DONT_TOUCH="true"*) wire A2131;
(*DONT_TOUCH="true"*) wire signed [7:0] C2141;
(*DONT_TOUCH="true"*) wire A2141;
(*DONT_TOUCH="true"*) wire signed [7:0] C2201;
(*DONT_TOUCH="true"*) wire A2201;
(*DONT_TOUCH="true"*) wire signed [7:0] C2211;
(*DONT_TOUCH="true"*) wire A2211;
(*DONT_TOUCH="true"*) wire signed [7:0] C2221;
(*DONT_TOUCH="true"*) wire A2221;
(*DONT_TOUCH="true"*) wire signed [7:0] C2231;
(*DONT_TOUCH="true"*) wire A2231;
(*DONT_TOUCH="true"*) wire signed [7:0] C2241;
(*DONT_TOUCH="true"*) wire A2241;
(*DONT_TOUCH="true"*) wire signed [7:0] C2301;
(*DONT_TOUCH="true"*) wire A2301;
(*DONT_TOUCH="true"*) wire signed [7:0] C2311;
(*DONT_TOUCH="true"*) wire A2311;
(*DONT_TOUCH="true"*) wire signed [7:0] C2321;
(*DONT_TOUCH="true"*) wire A2321;
(*DONT_TOUCH="true"*) wire signed [7:0] C2331;
(*DONT_TOUCH="true"*) wire A2331;
(*DONT_TOUCH="true"*) wire signed [7:0] C2341;
(*DONT_TOUCH="true"*) wire A2341;
(*DONT_TOUCH="true"*) wire signed [7:0] C2401;
(*DONT_TOUCH="true"*) wire A2401;
(*DONT_TOUCH="true"*) wire signed [7:0] C2411;
(*DONT_TOUCH="true"*) wire A2411;
(*DONT_TOUCH="true"*) wire signed [7:0] C2421;
(*DONT_TOUCH="true"*) wire A2421;
(*DONT_TOUCH="true"*) wire signed [7:0] C2431;
(*DONT_TOUCH="true"*) wire A2431;
(*DONT_TOUCH="true"*) wire signed [7:0] C2441;
(*DONT_TOUCH="true"*) wire A2441;
(*DONT_TOUCH="true"*) wire signed [7:0] C2002;
(*DONT_TOUCH="true"*) wire A2002;
(*DONT_TOUCH="true"*) wire signed [7:0] C2012;
(*DONT_TOUCH="true"*) wire A2012;
(*DONT_TOUCH="true"*) wire signed [7:0] C2022;
(*DONT_TOUCH="true"*) wire A2022;
(*DONT_TOUCH="true"*) wire signed [7:0] C2032;
(*DONT_TOUCH="true"*) wire A2032;
(*DONT_TOUCH="true"*) wire signed [7:0] C2042;
(*DONT_TOUCH="true"*) wire A2042;
(*DONT_TOUCH="true"*) wire signed [7:0] C2102;
(*DONT_TOUCH="true"*) wire A2102;
(*DONT_TOUCH="true"*) wire signed [7:0] C2112;
(*DONT_TOUCH="true"*) wire A2112;
(*DONT_TOUCH="true"*) wire signed [7:0] C2122;
(*DONT_TOUCH="true"*) wire A2122;
(*DONT_TOUCH="true"*) wire signed [7:0] C2132;
(*DONT_TOUCH="true"*) wire A2132;
(*DONT_TOUCH="true"*) wire signed [7:0] C2142;
(*DONT_TOUCH="true"*) wire A2142;
(*DONT_TOUCH="true"*) wire signed [7:0] C2202;
(*DONT_TOUCH="true"*) wire A2202;
(*DONT_TOUCH="true"*) wire signed [7:0] C2212;
(*DONT_TOUCH="true"*) wire A2212;
(*DONT_TOUCH="true"*) wire signed [7:0] C2222;
(*DONT_TOUCH="true"*) wire A2222;
(*DONT_TOUCH="true"*) wire signed [7:0] C2232;
(*DONT_TOUCH="true"*) wire A2232;
(*DONT_TOUCH="true"*) wire signed [7:0] C2242;
(*DONT_TOUCH="true"*) wire A2242;
(*DONT_TOUCH="true"*) wire signed [7:0] C2302;
(*DONT_TOUCH="true"*) wire A2302;
(*DONT_TOUCH="true"*) wire signed [7:0] C2312;
(*DONT_TOUCH="true"*) wire A2312;
(*DONT_TOUCH="true"*) wire signed [7:0] C2322;
(*DONT_TOUCH="true"*) wire A2322;
(*DONT_TOUCH="true"*) wire signed [7:0] C2332;
(*DONT_TOUCH="true"*) wire A2332;
(*DONT_TOUCH="true"*) wire signed [7:0] C2342;
(*DONT_TOUCH="true"*) wire A2342;
(*DONT_TOUCH="true"*) wire signed [7:0] C2402;
(*DONT_TOUCH="true"*) wire A2402;
(*DONT_TOUCH="true"*) wire signed [7:0] C2412;
(*DONT_TOUCH="true"*) wire A2412;
(*DONT_TOUCH="true"*) wire signed [7:0] C2422;
(*DONT_TOUCH="true"*) wire A2422;
(*DONT_TOUCH="true"*) wire signed [7:0] C2432;
(*DONT_TOUCH="true"*) wire A2432;
(*DONT_TOUCH="true"*) wire signed [7:0] C2442;
(*DONT_TOUCH="true"*) wire A2442;
(*DONT_TOUCH="true"*) wire signed [7:0] C2003;
(*DONT_TOUCH="true"*) wire A2003;
(*DONT_TOUCH="true"*) wire signed [7:0] C2013;
(*DONT_TOUCH="true"*) wire A2013;
(*DONT_TOUCH="true"*) wire signed [7:0] C2023;
(*DONT_TOUCH="true"*) wire A2023;
(*DONT_TOUCH="true"*) wire signed [7:0] C2033;
(*DONT_TOUCH="true"*) wire A2033;
(*DONT_TOUCH="true"*) wire signed [7:0] C2043;
(*DONT_TOUCH="true"*) wire A2043;
(*DONT_TOUCH="true"*) wire signed [7:0] C2103;
(*DONT_TOUCH="true"*) wire A2103;
(*DONT_TOUCH="true"*) wire signed [7:0] C2113;
(*DONT_TOUCH="true"*) wire A2113;
(*DONT_TOUCH="true"*) wire signed [7:0] C2123;
(*DONT_TOUCH="true"*) wire A2123;
(*DONT_TOUCH="true"*) wire signed [7:0] C2133;
(*DONT_TOUCH="true"*) wire A2133;
(*DONT_TOUCH="true"*) wire signed [7:0] C2143;
(*DONT_TOUCH="true"*) wire A2143;
(*DONT_TOUCH="true"*) wire signed [7:0] C2203;
(*DONT_TOUCH="true"*) wire A2203;
(*DONT_TOUCH="true"*) wire signed [7:0] C2213;
(*DONT_TOUCH="true"*) wire A2213;
(*DONT_TOUCH="true"*) wire signed [7:0] C2223;
(*DONT_TOUCH="true"*) wire A2223;
(*DONT_TOUCH="true"*) wire signed [7:0] C2233;
(*DONT_TOUCH="true"*) wire A2233;
(*DONT_TOUCH="true"*) wire signed [7:0] C2243;
(*DONT_TOUCH="true"*) wire A2243;
(*DONT_TOUCH="true"*) wire signed [7:0] C2303;
(*DONT_TOUCH="true"*) wire A2303;
(*DONT_TOUCH="true"*) wire signed [7:0] C2313;
(*DONT_TOUCH="true"*) wire A2313;
(*DONT_TOUCH="true"*) wire signed [7:0] C2323;
(*DONT_TOUCH="true"*) wire A2323;
(*DONT_TOUCH="true"*) wire signed [7:0] C2333;
(*DONT_TOUCH="true"*) wire A2333;
(*DONT_TOUCH="true"*) wire signed [7:0] C2343;
(*DONT_TOUCH="true"*) wire A2343;
(*DONT_TOUCH="true"*) wire signed [7:0] C2403;
(*DONT_TOUCH="true"*) wire A2403;
(*DONT_TOUCH="true"*) wire signed [7:0] C2413;
(*DONT_TOUCH="true"*) wire A2413;
(*DONT_TOUCH="true"*) wire signed [7:0] C2423;
(*DONT_TOUCH="true"*) wire A2423;
(*DONT_TOUCH="true"*) wire signed [7:0] C2433;
(*DONT_TOUCH="true"*) wire A2433;
(*DONT_TOUCH="true"*) wire signed [7:0] C2443;
(*DONT_TOUCH="true"*) wire A2443;
(*DONT_TOUCH="true"*) wire signed [7:0] C2004;
(*DONT_TOUCH="true"*) wire A2004;
(*DONT_TOUCH="true"*) wire signed [7:0] C2014;
(*DONT_TOUCH="true"*) wire A2014;
(*DONT_TOUCH="true"*) wire signed [7:0] C2024;
(*DONT_TOUCH="true"*) wire A2024;
(*DONT_TOUCH="true"*) wire signed [7:0] C2034;
(*DONT_TOUCH="true"*) wire A2034;
(*DONT_TOUCH="true"*) wire signed [7:0] C2044;
(*DONT_TOUCH="true"*) wire A2044;
(*DONT_TOUCH="true"*) wire signed [7:0] C2104;
(*DONT_TOUCH="true"*) wire A2104;
(*DONT_TOUCH="true"*) wire signed [7:0] C2114;
(*DONT_TOUCH="true"*) wire A2114;
(*DONT_TOUCH="true"*) wire signed [7:0] C2124;
(*DONT_TOUCH="true"*) wire A2124;
(*DONT_TOUCH="true"*) wire signed [7:0] C2134;
(*DONT_TOUCH="true"*) wire A2134;
(*DONT_TOUCH="true"*) wire signed [7:0] C2144;
(*DONT_TOUCH="true"*) wire A2144;
(*DONT_TOUCH="true"*) wire signed [7:0] C2204;
(*DONT_TOUCH="true"*) wire A2204;
(*DONT_TOUCH="true"*) wire signed [7:0] C2214;
(*DONT_TOUCH="true"*) wire A2214;
(*DONT_TOUCH="true"*) wire signed [7:0] C2224;
(*DONT_TOUCH="true"*) wire A2224;
(*DONT_TOUCH="true"*) wire signed [7:0] C2234;
(*DONT_TOUCH="true"*) wire A2234;
(*DONT_TOUCH="true"*) wire signed [7:0] C2244;
(*DONT_TOUCH="true"*) wire A2244;
(*DONT_TOUCH="true"*) wire signed [7:0] C2304;
(*DONT_TOUCH="true"*) wire A2304;
(*DONT_TOUCH="true"*) wire signed [7:0] C2314;
(*DONT_TOUCH="true"*) wire A2314;
(*DONT_TOUCH="true"*) wire signed [7:0] C2324;
(*DONT_TOUCH="true"*) wire A2324;
(*DONT_TOUCH="true"*) wire signed [7:0] C2334;
(*DONT_TOUCH="true"*) wire A2334;
(*DONT_TOUCH="true"*) wire signed [7:0] C2344;
(*DONT_TOUCH="true"*) wire A2344;
(*DONT_TOUCH="true"*) wire signed [7:0] C2404;
(*DONT_TOUCH="true"*) wire A2404;
(*DONT_TOUCH="true"*) wire signed [7:0] C2414;
(*DONT_TOUCH="true"*) wire A2414;
(*DONT_TOUCH="true"*) wire signed [7:0] C2424;
(*DONT_TOUCH="true"*) wire A2424;
(*DONT_TOUCH="true"*) wire signed [7:0] C2434;
(*DONT_TOUCH="true"*) wire A2434;
(*DONT_TOUCH="true"*) wire signed [7:0] C2444;
(*DONT_TOUCH="true"*) wire A2444;
(*DONT_TOUCH="true"*) wire signed [7:0] C2005;
(*DONT_TOUCH="true"*) wire A2005;
(*DONT_TOUCH="true"*) wire signed [7:0] C2015;
(*DONT_TOUCH="true"*) wire A2015;
(*DONT_TOUCH="true"*) wire signed [7:0] C2025;
(*DONT_TOUCH="true"*) wire A2025;
(*DONT_TOUCH="true"*) wire signed [7:0] C2035;
(*DONT_TOUCH="true"*) wire A2035;
(*DONT_TOUCH="true"*) wire signed [7:0] C2045;
(*DONT_TOUCH="true"*) wire A2045;
(*DONT_TOUCH="true"*) wire signed [7:0] C2105;
(*DONT_TOUCH="true"*) wire A2105;
(*DONT_TOUCH="true"*) wire signed [7:0] C2115;
(*DONT_TOUCH="true"*) wire A2115;
(*DONT_TOUCH="true"*) wire signed [7:0] C2125;
(*DONT_TOUCH="true"*) wire A2125;
(*DONT_TOUCH="true"*) wire signed [7:0] C2135;
(*DONT_TOUCH="true"*) wire A2135;
(*DONT_TOUCH="true"*) wire signed [7:0] C2145;
(*DONT_TOUCH="true"*) wire A2145;
(*DONT_TOUCH="true"*) wire signed [7:0] C2205;
(*DONT_TOUCH="true"*) wire A2205;
(*DONT_TOUCH="true"*) wire signed [7:0] C2215;
(*DONT_TOUCH="true"*) wire A2215;
(*DONT_TOUCH="true"*) wire signed [7:0] C2225;
(*DONT_TOUCH="true"*) wire A2225;
(*DONT_TOUCH="true"*) wire signed [7:0] C2235;
(*DONT_TOUCH="true"*) wire A2235;
(*DONT_TOUCH="true"*) wire signed [7:0] C2245;
(*DONT_TOUCH="true"*) wire A2245;
(*DONT_TOUCH="true"*) wire signed [7:0] C2305;
(*DONT_TOUCH="true"*) wire A2305;
(*DONT_TOUCH="true"*) wire signed [7:0] C2315;
(*DONT_TOUCH="true"*) wire A2315;
(*DONT_TOUCH="true"*) wire signed [7:0] C2325;
(*DONT_TOUCH="true"*) wire A2325;
(*DONT_TOUCH="true"*) wire signed [7:0] C2335;
(*DONT_TOUCH="true"*) wire A2335;
(*DONT_TOUCH="true"*) wire signed [7:0] C2345;
(*DONT_TOUCH="true"*) wire A2345;
(*DONT_TOUCH="true"*) wire signed [7:0] C2405;
(*DONT_TOUCH="true"*) wire A2405;
(*DONT_TOUCH="true"*) wire signed [7:0] C2415;
(*DONT_TOUCH="true"*) wire A2415;
(*DONT_TOUCH="true"*) wire signed [7:0] C2425;
(*DONT_TOUCH="true"*) wire A2425;
(*DONT_TOUCH="true"*) wire signed [7:0] C2435;
(*DONT_TOUCH="true"*) wire A2435;
(*DONT_TOUCH="true"*) wire signed [7:0] C2445;
(*DONT_TOUCH="true"*) wire A2445;
(*DONT_TOUCH="true"*) wire signed [7:0] C2006;
(*DONT_TOUCH="true"*) wire A2006;
(*DONT_TOUCH="true"*) wire signed [7:0] C2016;
(*DONT_TOUCH="true"*) wire A2016;
(*DONT_TOUCH="true"*) wire signed [7:0] C2026;
(*DONT_TOUCH="true"*) wire A2026;
(*DONT_TOUCH="true"*) wire signed [7:0] C2036;
(*DONT_TOUCH="true"*) wire A2036;
(*DONT_TOUCH="true"*) wire signed [7:0] C2046;
(*DONT_TOUCH="true"*) wire A2046;
(*DONT_TOUCH="true"*) wire signed [7:0] C2106;
(*DONT_TOUCH="true"*) wire A2106;
(*DONT_TOUCH="true"*) wire signed [7:0] C2116;
(*DONT_TOUCH="true"*) wire A2116;
(*DONT_TOUCH="true"*) wire signed [7:0] C2126;
(*DONT_TOUCH="true"*) wire A2126;
(*DONT_TOUCH="true"*) wire signed [7:0] C2136;
(*DONT_TOUCH="true"*) wire A2136;
(*DONT_TOUCH="true"*) wire signed [7:0] C2146;
(*DONT_TOUCH="true"*) wire A2146;
(*DONT_TOUCH="true"*) wire signed [7:0] C2206;
(*DONT_TOUCH="true"*) wire A2206;
(*DONT_TOUCH="true"*) wire signed [7:0] C2216;
(*DONT_TOUCH="true"*) wire A2216;
(*DONT_TOUCH="true"*) wire signed [7:0] C2226;
(*DONT_TOUCH="true"*) wire A2226;
(*DONT_TOUCH="true"*) wire signed [7:0] C2236;
(*DONT_TOUCH="true"*) wire A2236;
(*DONT_TOUCH="true"*) wire signed [7:0] C2246;
(*DONT_TOUCH="true"*) wire A2246;
(*DONT_TOUCH="true"*) wire signed [7:0] C2306;
(*DONT_TOUCH="true"*) wire A2306;
(*DONT_TOUCH="true"*) wire signed [7:0] C2316;
(*DONT_TOUCH="true"*) wire A2316;
(*DONT_TOUCH="true"*) wire signed [7:0] C2326;
(*DONT_TOUCH="true"*) wire A2326;
(*DONT_TOUCH="true"*) wire signed [7:0] C2336;
(*DONT_TOUCH="true"*) wire A2336;
(*DONT_TOUCH="true"*) wire signed [7:0] C2346;
(*DONT_TOUCH="true"*) wire A2346;
(*DONT_TOUCH="true"*) wire signed [7:0] C2406;
(*DONT_TOUCH="true"*) wire A2406;
(*DONT_TOUCH="true"*) wire signed [7:0] C2416;
(*DONT_TOUCH="true"*) wire A2416;
(*DONT_TOUCH="true"*) wire signed [7:0] C2426;
(*DONT_TOUCH="true"*) wire A2426;
(*DONT_TOUCH="true"*) wire signed [7:0] C2436;
(*DONT_TOUCH="true"*) wire A2436;
(*DONT_TOUCH="true"*) wire signed [7:0] C2446;
(*DONT_TOUCH="true"*) wire A2446;
(*DONT_TOUCH="true"*) wire signed [7:0] C2007;
(*DONT_TOUCH="true"*) wire A2007;
(*DONT_TOUCH="true"*) wire signed [7:0] C2017;
(*DONT_TOUCH="true"*) wire A2017;
(*DONT_TOUCH="true"*) wire signed [7:0] C2027;
(*DONT_TOUCH="true"*) wire A2027;
(*DONT_TOUCH="true"*) wire signed [7:0] C2037;
(*DONT_TOUCH="true"*) wire A2037;
(*DONT_TOUCH="true"*) wire signed [7:0] C2047;
(*DONT_TOUCH="true"*) wire A2047;
(*DONT_TOUCH="true"*) wire signed [7:0] C2107;
(*DONT_TOUCH="true"*) wire A2107;
(*DONT_TOUCH="true"*) wire signed [7:0] C2117;
(*DONT_TOUCH="true"*) wire A2117;
(*DONT_TOUCH="true"*) wire signed [7:0] C2127;
(*DONT_TOUCH="true"*) wire A2127;
(*DONT_TOUCH="true"*) wire signed [7:0] C2137;
(*DONT_TOUCH="true"*) wire A2137;
(*DONT_TOUCH="true"*) wire signed [7:0] C2147;
(*DONT_TOUCH="true"*) wire A2147;
(*DONT_TOUCH="true"*) wire signed [7:0] C2207;
(*DONT_TOUCH="true"*) wire A2207;
(*DONT_TOUCH="true"*) wire signed [7:0] C2217;
(*DONT_TOUCH="true"*) wire A2217;
(*DONT_TOUCH="true"*) wire signed [7:0] C2227;
(*DONT_TOUCH="true"*) wire A2227;
(*DONT_TOUCH="true"*) wire signed [7:0] C2237;
(*DONT_TOUCH="true"*) wire A2237;
(*DONT_TOUCH="true"*) wire signed [7:0] C2247;
(*DONT_TOUCH="true"*) wire A2247;
(*DONT_TOUCH="true"*) wire signed [7:0] C2307;
(*DONT_TOUCH="true"*) wire A2307;
(*DONT_TOUCH="true"*) wire signed [7:0] C2317;
(*DONT_TOUCH="true"*) wire A2317;
(*DONT_TOUCH="true"*) wire signed [7:0] C2327;
(*DONT_TOUCH="true"*) wire A2327;
(*DONT_TOUCH="true"*) wire signed [7:0] C2337;
(*DONT_TOUCH="true"*) wire A2337;
(*DONT_TOUCH="true"*) wire signed [7:0] C2347;
(*DONT_TOUCH="true"*) wire A2347;
(*DONT_TOUCH="true"*) wire signed [7:0] C2407;
(*DONT_TOUCH="true"*) wire A2407;
(*DONT_TOUCH="true"*) wire signed [7:0] C2417;
(*DONT_TOUCH="true"*) wire A2417;
(*DONT_TOUCH="true"*) wire signed [7:0] C2427;
(*DONT_TOUCH="true"*) wire A2427;
(*DONT_TOUCH="true"*) wire signed [7:0] C2437;
(*DONT_TOUCH="true"*) wire A2437;
(*DONT_TOUCH="true"*) wire signed [7:0] C2447;
(*DONT_TOUCH="true"*) wire A2447;
(*DONT_TOUCH="true"*) wire signed [7:0] C2008;
(*DONT_TOUCH="true"*) wire A2008;
(*DONT_TOUCH="true"*) wire signed [7:0] C2018;
(*DONT_TOUCH="true"*) wire A2018;
(*DONT_TOUCH="true"*) wire signed [7:0] C2028;
(*DONT_TOUCH="true"*) wire A2028;
(*DONT_TOUCH="true"*) wire signed [7:0] C2038;
(*DONT_TOUCH="true"*) wire A2038;
(*DONT_TOUCH="true"*) wire signed [7:0] C2048;
(*DONT_TOUCH="true"*) wire A2048;
(*DONT_TOUCH="true"*) wire signed [7:0] C2108;
(*DONT_TOUCH="true"*) wire A2108;
(*DONT_TOUCH="true"*) wire signed [7:0] C2118;
(*DONT_TOUCH="true"*) wire A2118;
(*DONT_TOUCH="true"*) wire signed [7:0] C2128;
(*DONT_TOUCH="true"*) wire A2128;
(*DONT_TOUCH="true"*) wire signed [7:0] C2138;
(*DONT_TOUCH="true"*) wire A2138;
(*DONT_TOUCH="true"*) wire signed [7:0] C2148;
(*DONT_TOUCH="true"*) wire A2148;
(*DONT_TOUCH="true"*) wire signed [7:0] C2208;
(*DONT_TOUCH="true"*) wire A2208;
(*DONT_TOUCH="true"*) wire signed [7:0] C2218;
(*DONT_TOUCH="true"*) wire A2218;
(*DONT_TOUCH="true"*) wire signed [7:0] C2228;
(*DONT_TOUCH="true"*) wire A2228;
(*DONT_TOUCH="true"*) wire signed [7:0] C2238;
(*DONT_TOUCH="true"*) wire A2238;
(*DONT_TOUCH="true"*) wire signed [7:0] C2248;
(*DONT_TOUCH="true"*) wire A2248;
(*DONT_TOUCH="true"*) wire signed [7:0] C2308;
(*DONT_TOUCH="true"*) wire A2308;
(*DONT_TOUCH="true"*) wire signed [7:0] C2318;
(*DONT_TOUCH="true"*) wire A2318;
(*DONT_TOUCH="true"*) wire signed [7:0] C2328;
(*DONT_TOUCH="true"*) wire A2328;
(*DONT_TOUCH="true"*) wire signed [7:0] C2338;
(*DONT_TOUCH="true"*) wire A2338;
(*DONT_TOUCH="true"*) wire signed [7:0] C2348;
(*DONT_TOUCH="true"*) wire A2348;
(*DONT_TOUCH="true"*) wire signed [7:0] C2408;
(*DONT_TOUCH="true"*) wire A2408;
(*DONT_TOUCH="true"*) wire signed [7:0] C2418;
(*DONT_TOUCH="true"*) wire A2418;
(*DONT_TOUCH="true"*) wire signed [7:0] C2428;
(*DONT_TOUCH="true"*) wire A2428;
(*DONT_TOUCH="true"*) wire signed [7:0] C2438;
(*DONT_TOUCH="true"*) wire A2438;
(*DONT_TOUCH="true"*) wire signed [7:0] C2448;
(*DONT_TOUCH="true"*) wire A2448;
(*DONT_TOUCH="true"*) wire signed [7:0] C2009;
(*DONT_TOUCH="true"*) wire A2009;
(*DONT_TOUCH="true"*) wire signed [7:0] C2019;
(*DONT_TOUCH="true"*) wire A2019;
(*DONT_TOUCH="true"*) wire signed [7:0] C2029;
(*DONT_TOUCH="true"*) wire A2029;
(*DONT_TOUCH="true"*) wire signed [7:0] C2039;
(*DONT_TOUCH="true"*) wire A2039;
(*DONT_TOUCH="true"*) wire signed [7:0] C2049;
(*DONT_TOUCH="true"*) wire A2049;
(*DONT_TOUCH="true"*) wire signed [7:0] C2109;
(*DONT_TOUCH="true"*) wire A2109;
(*DONT_TOUCH="true"*) wire signed [7:0] C2119;
(*DONT_TOUCH="true"*) wire A2119;
(*DONT_TOUCH="true"*) wire signed [7:0] C2129;
(*DONT_TOUCH="true"*) wire A2129;
(*DONT_TOUCH="true"*) wire signed [7:0] C2139;
(*DONT_TOUCH="true"*) wire A2139;
(*DONT_TOUCH="true"*) wire signed [7:0] C2149;
(*DONT_TOUCH="true"*) wire A2149;
(*DONT_TOUCH="true"*) wire signed [7:0] C2209;
(*DONT_TOUCH="true"*) wire A2209;
(*DONT_TOUCH="true"*) wire signed [7:0] C2219;
(*DONT_TOUCH="true"*) wire A2219;
(*DONT_TOUCH="true"*) wire signed [7:0] C2229;
(*DONT_TOUCH="true"*) wire A2229;
(*DONT_TOUCH="true"*) wire signed [7:0] C2239;
(*DONT_TOUCH="true"*) wire A2239;
(*DONT_TOUCH="true"*) wire signed [7:0] C2249;
(*DONT_TOUCH="true"*) wire A2249;
(*DONT_TOUCH="true"*) wire signed [7:0] C2309;
(*DONT_TOUCH="true"*) wire A2309;
(*DONT_TOUCH="true"*) wire signed [7:0] C2319;
(*DONT_TOUCH="true"*) wire A2319;
(*DONT_TOUCH="true"*) wire signed [7:0] C2329;
(*DONT_TOUCH="true"*) wire A2329;
(*DONT_TOUCH="true"*) wire signed [7:0] C2339;
(*DONT_TOUCH="true"*) wire A2339;
(*DONT_TOUCH="true"*) wire signed [7:0] C2349;
(*DONT_TOUCH="true"*) wire A2349;
(*DONT_TOUCH="true"*) wire signed [7:0] C2409;
(*DONT_TOUCH="true"*) wire A2409;
(*DONT_TOUCH="true"*) wire signed [7:0] C2419;
(*DONT_TOUCH="true"*) wire A2419;
(*DONT_TOUCH="true"*) wire signed [7:0] C2429;
(*DONT_TOUCH="true"*) wire A2429;
(*DONT_TOUCH="true"*) wire signed [7:0] C2439;
(*DONT_TOUCH="true"*) wire A2439;
(*DONT_TOUCH="true"*) wire signed [7:0] C2449;
(*DONT_TOUCH="true"*) wire A2449;
(*DONT_TOUCH="true"*) wire signed [7:0] C200A;
(*DONT_TOUCH="true"*) wire A200A;
(*DONT_TOUCH="true"*) wire signed [7:0] C201A;
(*DONT_TOUCH="true"*) wire A201A;
(*DONT_TOUCH="true"*) wire signed [7:0] C202A;
(*DONT_TOUCH="true"*) wire A202A;
(*DONT_TOUCH="true"*) wire signed [7:0] C203A;
(*DONT_TOUCH="true"*) wire A203A;
(*DONT_TOUCH="true"*) wire signed [7:0] C204A;
(*DONT_TOUCH="true"*) wire A204A;
(*DONT_TOUCH="true"*) wire signed [7:0] C210A;
(*DONT_TOUCH="true"*) wire A210A;
(*DONT_TOUCH="true"*) wire signed [7:0] C211A;
(*DONT_TOUCH="true"*) wire A211A;
(*DONT_TOUCH="true"*) wire signed [7:0] C212A;
(*DONT_TOUCH="true"*) wire A212A;
(*DONT_TOUCH="true"*) wire signed [7:0] C213A;
(*DONT_TOUCH="true"*) wire A213A;
(*DONT_TOUCH="true"*) wire signed [7:0] C214A;
(*DONT_TOUCH="true"*) wire A214A;
(*DONT_TOUCH="true"*) wire signed [7:0] C220A;
(*DONT_TOUCH="true"*) wire A220A;
(*DONT_TOUCH="true"*) wire signed [7:0] C221A;
(*DONT_TOUCH="true"*) wire A221A;
(*DONT_TOUCH="true"*) wire signed [7:0] C222A;
(*DONT_TOUCH="true"*) wire A222A;
(*DONT_TOUCH="true"*) wire signed [7:0] C223A;
(*DONT_TOUCH="true"*) wire A223A;
(*DONT_TOUCH="true"*) wire signed [7:0] C224A;
(*DONT_TOUCH="true"*) wire A224A;
(*DONT_TOUCH="true"*) wire signed [7:0] C230A;
(*DONT_TOUCH="true"*) wire A230A;
(*DONT_TOUCH="true"*) wire signed [7:0] C231A;
(*DONT_TOUCH="true"*) wire A231A;
(*DONT_TOUCH="true"*) wire signed [7:0] C232A;
(*DONT_TOUCH="true"*) wire A232A;
(*DONT_TOUCH="true"*) wire signed [7:0] C233A;
(*DONT_TOUCH="true"*) wire A233A;
(*DONT_TOUCH="true"*) wire signed [7:0] C234A;
(*DONT_TOUCH="true"*) wire A234A;
(*DONT_TOUCH="true"*) wire signed [7:0] C240A;
(*DONT_TOUCH="true"*) wire A240A;
(*DONT_TOUCH="true"*) wire signed [7:0] C241A;
(*DONT_TOUCH="true"*) wire A241A;
(*DONT_TOUCH="true"*) wire signed [7:0] C242A;
(*DONT_TOUCH="true"*) wire A242A;
(*DONT_TOUCH="true"*) wire signed [7:0] C243A;
(*DONT_TOUCH="true"*) wire A243A;
(*DONT_TOUCH="true"*) wire signed [7:0] C244A;
(*DONT_TOUCH="true"*) wire A244A;
(*DONT_TOUCH="true"*) wire signed [7:0] C200B;
(*DONT_TOUCH="true"*) wire A200B;
(*DONT_TOUCH="true"*) wire signed [7:0] C201B;
(*DONT_TOUCH="true"*) wire A201B;
(*DONT_TOUCH="true"*) wire signed [7:0] C202B;
(*DONT_TOUCH="true"*) wire A202B;
(*DONT_TOUCH="true"*) wire signed [7:0] C203B;
(*DONT_TOUCH="true"*) wire A203B;
(*DONT_TOUCH="true"*) wire signed [7:0] C204B;
(*DONT_TOUCH="true"*) wire A204B;
(*DONT_TOUCH="true"*) wire signed [7:0] C210B;
(*DONT_TOUCH="true"*) wire A210B;
(*DONT_TOUCH="true"*) wire signed [7:0] C211B;
(*DONT_TOUCH="true"*) wire A211B;
(*DONT_TOUCH="true"*) wire signed [7:0] C212B;
(*DONT_TOUCH="true"*) wire A212B;
(*DONT_TOUCH="true"*) wire signed [7:0] C213B;
(*DONT_TOUCH="true"*) wire A213B;
(*DONT_TOUCH="true"*) wire signed [7:0] C214B;
(*DONT_TOUCH="true"*) wire A214B;
(*DONT_TOUCH="true"*) wire signed [7:0] C220B;
(*DONT_TOUCH="true"*) wire A220B;
(*DONT_TOUCH="true"*) wire signed [7:0] C221B;
(*DONT_TOUCH="true"*) wire A221B;
(*DONT_TOUCH="true"*) wire signed [7:0] C222B;
(*DONT_TOUCH="true"*) wire A222B;
(*DONT_TOUCH="true"*) wire signed [7:0] C223B;
(*DONT_TOUCH="true"*) wire A223B;
(*DONT_TOUCH="true"*) wire signed [7:0] C224B;
(*DONT_TOUCH="true"*) wire A224B;
(*DONT_TOUCH="true"*) wire signed [7:0] C230B;
(*DONT_TOUCH="true"*) wire A230B;
(*DONT_TOUCH="true"*) wire signed [7:0] C231B;
(*DONT_TOUCH="true"*) wire A231B;
(*DONT_TOUCH="true"*) wire signed [7:0] C232B;
(*DONT_TOUCH="true"*) wire A232B;
(*DONT_TOUCH="true"*) wire signed [7:0] C233B;
(*DONT_TOUCH="true"*) wire A233B;
(*DONT_TOUCH="true"*) wire signed [7:0] C234B;
(*DONT_TOUCH="true"*) wire A234B;
(*DONT_TOUCH="true"*) wire signed [7:0] C240B;
(*DONT_TOUCH="true"*) wire A240B;
(*DONT_TOUCH="true"*) wire signed [7:0] C241B;
(*DONT_TOUCH="true"*) wire A241B;
(*DONT_TOUCH="true"*) wire signed [7:0] C242B;
(*DONT_TOUCH="true"*) wire A242B;
(*DONT_TOUCH="true"*) wire signed [7:0] C243B;
(*DONT_TOUCH="true"*) wire A243B;
(*DONT_TOUCH="true"*) wire signed [7:0] C244B;
(*DONT_TOUCH="true"*) wire A244B;
(*DONT_TOUCH="true"*) wire signed [7:0] C200C;
(*DONT_TOUCH="true"*) wire A200C;
(*DONT_TOUCH="true"*) wire signed [7:0] C201C;
(*DONT_TOUCH="true"*) wire A201C;
(*DONT_TOUCH="true"*) wire signed [7:0] C202C;
(*DONT_TOUCH="true"*) wire A202C;
(*DONT_TOUCH="true"*) wire signed [7:0] C203C;
(*DONT_TOUCH="true"*) wire A203C;
(*DONT_TOUCH="true"*) wire signed [7:0] C204C;
(*DONT_TOUCH="true"*) wire A204C;
(*DONT_TOUCH="true"*) wire signed [7:0] C210C;
(*DONT_TOUCH="true"*) wire A210C;
(*DONT_TOUCH="true"*) wire signed [7:0] C211C;
(*DONT_TOUCH="true"*) wire A211C;
(*DONT_TOUCH="true"*) wire signed [7:0] C212C;
(*DONT_TOUCH="true"*) wire A212C;
(*DONT_TOUCH="true"*) wire signed [7:0] C213C;
(*DONT_TOUCH="true"*) wire A213C;
(*DONT_TOUCH="true"*) wire signed [7:0] C214C;
(*DONT_TOUCH="true"*) wire A214C;
(*DONT_TOUCH="true"*) wire signed [7:0] C220C;
(*DONT_TOUCH="true"*) wire A220C;
(*DONT_TOUCH="true"*) wire signed [7:0] C221C;
(*DONT_TOUCH="true"*) wire A221C;
(*DONT_TOUCH="true"*) wire signed [7:0] C222C;
(*DONT_TOUCH="true"*) wire A222C;
(*DONT_TOUCH="true"*) wire signed [7:0] C223C;
(*DONT_TOUCH="true"*) wire A223C;
(*DONT_TOUCH="true"*) wire signed [7:0] C224C;
(*DONT_TOUCH="true"*) wire A224C;
(*DONT_TOUCH="true"*) wire signed [7:0] C230C;
(*DONT_TOUCH="true"*) wire A230C;
(*DONT_TOUCH="true"*) wire signed [7:0] C231C;
(*DONT_TOUCH="true"*) wire A231C;
(*DONT_TOUCH="true"*) wire signed [7:0] C232C;
(*DONT_TOUCH="true"*) wire A232C;
(*DONT_TOUCH="true"*) wire signed [7:0] C233C;
(*DONT_TOUCH="true"*) wire A233C;
(*DONT_TOUCH="true"*) wire signed [7:0] C234C;
(*DONT_TOUCH="true"*) wire A234C;
(*DONT_TOUCH="true"*) wire signed [7:0] C240C;
(*DONT_TOUCH="true"*) wire A240C;
(*DONT_TOUCH="true"*) wire signed [7:0] C241C;
(*DONT_TOUCH="true"*) wire A241C;
(*DONT_TOUCH="true"*) wire signed [7:0] C242C;
(*DONT_TOUCH="true"*) wire A242C;
(*DONT_TOUCH="true"*) wire signed [7:0] C243C;
(*DONT_TOUCH="true"*) wire A243C;
(*DONT_TOUCH="true"*) wire signed [7:0] C244C;
(*DONT_TOUCH="true"*) wire A244C;
(*DONT_TOUCH="true"*) wire signed [7:0] C200D;
(*DONT_TOUCH="true"*) wire A200D;
(*DONT_TOUCH="true"*) wire signed [7:0] C201D;
(*DONT_TOUCH="true"*) wire A201D;
(*DONT_TOUCH="true"*) wire signed [7:0] C202D;
(*DONT_TOUCH="true"*) wire A202D;
(*DONT_TOUCH="true"*) wire signed [7:0] C203D;
(*DONT_TOUCH="true"*) wire A203D;
(*DONT_TOUCH="true"*) wire signed [7:0] C204D;
(*DONT_TOUCH="true"*) wire A204D;
(*DONT_TOUCH="true"*) wire signed [7:0] C210D;
(*DONT_TOUCH="true"*) wire A210D;
(*DONT_TOUCH="true"*) wire signed [7:0] C211D;
(*DONT_TOUCH="true"*) wire A211D;
(*DONT_TOUCH="true"*) wire signed [7:0] C212D;
(*DONT_TOUCH="true"*) wire A212D;
(*DONT_TOUCH="true"*) wire signed [7:0] C213D;
(*DONT_TOUCH="true"*) wire A213D;
(*DONT_TOUCH="true"*) wire signed [7:0] C214D;
(*DONT_TOUCH="true"*) wire A214D;
(*DONT_TOUCH="true"*) wire signed [7:0] C220D;
(*DONT_TOUCH="true"*) wire A220D;
(*DONT_TOUCH="true"*) wire signed [7:0] C221D;
(*DONT_TOUCH="true"*) wire A221D;
(*DONT_TOUCH="true"*) wire signed [7:0] C222D;
(*DONT_TOUCH="true"*) wire A222D;
(*DONT_TOUCH="true"*) wire signed [7:0] C223D;
(*DONT_TOUCH="true"*) wire A223D;
(*DONT_TOUCH="true"*) wire signed [7:0] C224D;
(*DONT_TOUCH="true"*) wire A224D;
(*DONT_TOUCH="true"*) wire signed [7:0] C230D;
(*DONT_TOUCH="true"*) wire A230D;
(*DONT_TOUCH="true"*) wire signed [7:0] C231D;
(*DONT_TOUCH="true"*) wire A231D;
(*DONT_TOUCH="true"*) wire signed [7:0] C232D;
(*DONT_TOUCH="true"*) wire A232D;
(*DONT_TOUCH="true"*) wire signed [7:0] C233D;
(*DONT_TOUCH="true"*) wire A233D;
(*DONT_TOUCH="true"*) wire signed [7:0] C234D;
(*DONT_TOUCH="true"*) wire A234D;
(*DONT_TOUCH="true"*) wire signed [7:0] C240D;
(*DONT_TOUCH="true"*) wire A240D;
(*DONT_TOUCH="true"*) wire signed [7:0] C241D;
(*DONT_TOUCH="true"*) wire A241D;
(*DONT_TOUCH="true"*) wire signed [7:0] C242D;
(*DONT_TOUCH="true"*) wire A242D;
(*DONT_TOUCH="true"*) wire signed [7:0] C243D;
(*DONT_TOUCH="true"*) wire A243D;
(*DONT_TOUCH="true"*) wire signed [7:0] C244D;
(*DONT_TOUCH="true"*) wire A244D;
(*DONT_TOUCH="true"*) wire signed [7:0] C200E;
(*DONT_TOUCH="true"*) wire A200E;
(*DONT_TOUCH="true"*) wire signed [7:0] C201E;
(*DONT_TOUCH="true"*) wire A201E;
(*DONT_TOUCH="true"*) wire signed [7:0] C202E;
(*DONT_TOUCH="true"*) wire A202E;
(*DONT_TOUCH="true"*) wire signed [7:0] C203E;
(*DONT_TOUCH="true"*) wire A203E;
(*DONT_TOUCH="true"*) wire signed [7:0] C204E;
(*DONT_TOUCH="true"*) wire A204E;
(*DONT_TOUCH="true"*) wire signed [7:0] C210E;
(*DONT_TOUCH="true"*) wire A210E;
(*DONT_TOUCH="true"*) wire signed [7:0] C211E;
(*DONT_TOUCH="true"*) wire A211E;
(*DONT_TOUCH="true"*) wire signed [7:0] C212E;
(*DONT_TOUCH="true"*) wire A212E;
(*DONT_TOUCH="true"*) wire signed [7:0] C213E;
(*DONT_TOUCH="true"*) wire A213E;
(*DONT_TOUCH="true"*) wire signed [7:0] C214E;
(*DONT_TOUCH="true"*) wire A214E;
(*DONT_TOUCH="true"*) wire signed [7:0] C220E;
(*DONT_TOUCH="true"*) wire A220E;
(*DONT_TOUCH="true"*) wire signed [7:0] C221E;
(*DONT_TOUCH="true"*) wire A221E;
(*DONT_TOUCH="true"*) wire signed [7:0] C222E;
(*DONT_TOUCH="true"*) wire A222E;
(*DONT_TOUCH="true"*) wire signed [7:0] C223E;
(*DONT_TOUCH="true"*) wire A223E;
(*DONT_TOUCH="true"*) wire signed [7:0] C224E;
(*DONT_TOUCH="true"*) wire A224E;
(*DONT_TOUCH="true"*) wire signed [7:0] C230E;
(*DONT_TOUCH="true"*) wire A230E;
(*DONT_TOUCH="true"*) wire signed [7:0] C231E;
(*DONT_TOUCH="true"*) wire A231E;
(*DONT_TOUCH="true"*) wire signed [7:0] C232E;
(*DONT_TOUCH="true"*) wire A232E;
(*DONT_TOUCH="true"*) wire signed [7:0] C233E;
(*DONT_TOUCH="true"*) wire A233E;
(*DONT_TOUCH="true"*) wire signed [7:0] C234E;
(*DONT_TOUCH="true"*) wire A234E;
(*DONT_TOUCH="true"*) wire signed [7:0] C240E;
(*DONT_TOUCH="true"*) wire A240E;
(*DONT_TOUCH="true"*) wire signed [7:0] C241E;
(*DONT_TOUCH="true"*) wire A241E;
(*DONT_TOUCH="true"*) wire signed [7:0] C242E;
(*DONT_TOUCH="true"*) wire A242E;
(*DONT_TOUCH="true"*) wire signed [7:0] C243E;
(*DONT_TOUCH="true"*) wire A243E;
(*DONT_TOUCH="true"*) wire signed [7:0] C244E;
(*DONT_TOUCH="true"*) wire A244E;
(*DONT_TOUCH="true"*) wire signed [7:0] C200F;
(*DONT_TOUCH="true"*) wire A200F;
(*DONT_TOUCH="true"*) wire signed [7:0] C201F;
(*DONT_TOUCH="true"*) wire A201F;
(*DONT_TOUCH="true"*) wire signed [7:0] C202F;
(*DONT_TOUCH="true"*) wire A202F;
(*DONT_TOUCH="true"*) wire signed [7:0] C203F;
(*DONT_TOUCH="true"*) wire A203F;
(*DONT_TOUCH="true"*) wire signed [7:0] C204F;
(*DONT_TOUCH="true"*) wire A204F;
(*DONT_TOUCH="true"*) wire signed [7:0] C210F;
(*DONT_TOUCH="true"*) wire A210F;
(*DONT_TOUCH="true"*) wire signed [7:0] C211F;
(*DONT_TOUCH="true"*) wire A211F;
(*DONT_TOUCH="true"*) wire signed [7:0] C212F;
(*DONT_TOUCH="true"*) wire A212F;
(*DONT_TOUCH="true"*) wire signed [7:0] C213F;
(*DONT_TOUCH="true"*) wire A213F;
(*DONT_TOUCH="true"*) wire signed [7:0] C214F;
(*DONT_TOUCH="true"*) wire A214F;
(*DONT_TOUCH="true"*) wire signed [7:0] C220F;
(*DONT_TOUCH="true"*) wire A220F;
(*DONT_TOUCH="true"*) wire signed [7:0] C221F;
(*DONT_TOUCH="true"*) wire A221F;
(*DONT_TOUCH="true"*) wire signed [7:0] C222F;
(*DONT_TOUCH="true"*) wire A222F;
(*DONT_TOUCH="true"*) wire signed [7:0] C223F;
(*DONT_TOUCH="true"*) wire A223F;
(*DONT_TOUCH="true"*) wire signed [7:0] C224F;
(*DONT_TOUCH="true"*) wire A224F;
(*DONT_TOUCH="true"*) wire signed [7:0] C230F;
(*DONT_TOUCH="true"*) wire A230F;
(*DONT_TOUCH="true"*) wire signed [7:0] C231F;
(*DONT_TOUCH="true"*) wire A231F;
(*DONT_TOUCH="true"*) wire signed [7:0] C232F;
(*DONT_TOUCH="true"*) wire A232F;
(*DONT_TOUCH="true"*) wire signed [7:0] C233F;
(*DONT_TOUCH="true"*) wire A233F;
(*DONT_TOUCH="true"*) wire signed [7:0] C234F;
(*DONT_TOUCH="true"*) wire A234F;
(*DONT_TOUCH="true"*) wire signed [7:0] C240F;
(*DONT_TOUCH="true"*) wire A240F;
(*DONT_TOUCH="true"*) wire signed [7:0] C241F;
(*DONT_TOUCH="true"*) wire A241F;
(*DONT_TOUCH="true"*) wire signed [7:0] C242F;
(*DONT_TOUCH="true"*) wire A242F;
(*DONT_TOUCH="true"*) wire signed [7:0] C243F;
(*DONT_TOUCH="true"*) wire A243F;
(*DONT_TOUCH="true"*) wire signed [7:0] C244F;
(*DONT_TOUCH="true"*) wire A244F;
DFF_save_fm DFF_P0(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2000));
DFF_save_fm DFF_P1(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2010));
DFF_save_fm DFF_P2(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2020));
DFF_save_fm DFF_P3(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2030));
DFF_save_fm DFF_P4(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2040));
DFF_save_fm DFF_P5(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2050));
DFF_save_fm DFF_P6(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2060));
DFF_save_fm DFF_P7(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2100));
DFF_save_fm DFF_P8(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2110));
DFF_save_fm DFF_P9(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2120));
DFF_save_fm DFF_P10(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2130));
DFF_save_fm DFF_P11(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2140));
DFF_save_fm DFF_P12(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2150));
DFF_save_fm DFF_P13(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2160));
DFF_save_fm DFF_P14(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2200));
DFF_save_fm DFF_P15(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2210));
DFF_save_fm DFF_P16(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2220));
DFF_save_fm DFF_P17(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2230));
DFF_save_fm DFF_P18(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2240));
DFF_save_fm DFF_P19(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2250));
DFF_save_fm DFF_P20(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2260));
DFF_save_fm DFF_P21(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2300));
DFF_save_fm DFF_P22(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2310));
DFF_save_fm DFF_P23(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2320));
DFF_save_fm DFF_P24(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2330));
DFF_save_fm DFF_P25(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2340));
DFF_save_fm DFF_P26(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2350));
DFF_save_fm DFF_P27(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2360));
DFF_save_fm DFF_P28(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2400));
DFF_save_fm DFF_P29(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2410));
DFF_save_fm DFF_P30(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2420));
DFF_save_fm DFF_P31(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2430));
DFF_save_fm DFF_P32(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2440));
DFF_save_fm DFF_P33(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2450));
DFF_save_fm DFF_P34(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2460));
DFF_save_fm DFF_P35(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2500));
DFF_save_fm DFF_P36(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2510));
DFF_save_fm DFF_P37(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2520));
DFF_save_fm DFF_P38(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2530));
DFF_save_fm DFF_P39(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2540));
DFF_save_fm DFF_P40(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2550));
DFF_save_fm DFF_P41(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2560));
DFF_save_fm DFF_P42(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2600));
DFF_save_fm DFF_P43(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2610));
DFF_save_fm DFF_P44(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2620));
DFF_save_fm DFF_P45(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2630));
DFF_save_fm DFF_P46(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2640));
DFF_save_fm DFF_P47(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2650));
DFF_save_fm DFF_P48(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2660));
DFF_save_fm DFF_P49(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2001));
DFF_save_fm DFF_P50(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2011));
DFF_save_fm DFF_P51(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2021));
DFF_save_fm DFF_P52(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2031));
DFF_save_fm DFF_P53(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2041));
DFF_save_fm DFF_P54(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2051));
DFF_save_fm DFF_P55(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2061));
DFF_save_fm DFF_P56(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2101));
DFF_save_fm DFF_P57(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2111));
DFF_save_fm DFF_P58(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2121));
DFF_save_fm DFF_P59(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2131));
DFF_save_fm DFF_P60(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2141));
DFF_save_fm DFF_P61(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2151));
DFF_save_fm DFF_P62(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2161));
DFF_save_fm DFF_P63(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2201));
DFF_save_fm DFF_P64(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2211));
DFF_save_fm DFF_P65(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2221));
DFF_save_fm DFF_P66(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2231));
DFF_save_fm DFF_P67(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2241));
DFF_save_fm DFF_P68(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2251));
DFF_save_fm DFF_P69(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2261));
DFF_save_fm DFF_P70(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2301));
DFF_save_fm DFF_P71(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2311));
DFF_save_fm DFF_P72(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2321));
DFF_save_fm DFF_P73(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2331));
DFF_save_fm DFF_P74(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2341));
DFF_save_fm DFF_P75(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2351));
DFF_save_fm DFF_P76(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2361));
DFF_save_fm DFF_P77(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2401));
DFF_save_fm DFF_P78(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2411));
DFF_save_fm DFF_P79(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2421));
DFF_save_fm DFF_P80(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2431));
DFF_save_fm DFF_P81(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2441));
DFF_save_fm DFF_P82(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2451));
DFF_save_fm DFF_P83(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2461));
DFF_save_fm DFF_P84(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2501));
DFF_save_fm DFF_P85(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2511));
DFF_save_fm DFF_P86(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2521));
DFF_save_fm DFF_P87(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2531));
DFF_save_fm DFF_P88(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2541));
DFF_save_fm DFF_P89(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2551));
DFF_save_fm DFF_P90(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2561));
DFF_save_fm DFF_P91(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2601));
DFF_save_fm DFF_P92(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2611));
DFF_save_fm DFF_P93(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2621));
DFF_save_fm DFF_P94(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2631));
DFF_save_fm DFF_P95(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2641));
DFF_save_fm DFF_P96(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2651));
DFF_save_fm DFF_P97(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2661));
DFF_save_fm DFF_P98(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2002));
DFF_save_fm DFF_P99(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2012));
DFF_save_fm DFF_P100(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2022));
DFF_save_fm DFF_P101(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2032));
DFF_save_fm DFF_P102(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2042));
DFF_save_fm DFF_P103(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2052));
DFF_save_fm DFF_P104(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2062));
DFF_save_fm DFF_P105(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2102));
DFF_save_fm DFF_P106(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2112));
DFF_save_fm DFF_P107(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2122));
DFF_save_fm DFF_P108(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2132));
DFF_save_fm DFF_P109(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2142));
DFF_save_fm DFF_P110(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2152));
DFF_save_fm DFF_P111(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2162));
DFF_save_fm DFF_P112(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2202));
DFF_save_fm DFF_P113(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2212));
DFF_save_fm DFF_P114(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2222));
DFF_save_fm DFF_P115(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2232));
DFF_save_fm DFF_P116(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2242));
DFF_save_fm DFF_P117(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2252));
DFF_save_fm DFF_P118(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2262));
DFF_save_fm DFF_P119(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2302));
DFF_save_fm DFF_P120(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2312));
DFF_save_fm DFF_P121(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2322));
DFF_save_fm DFF_P122(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2332));
DFF_save_fm DFF_P123(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2342));
DFF_save_fm DFF_P124(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2352));
DFF_save_fm DFF_P125(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2362));
DFF_save_fm DFF_P126(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2402));
DFF_save_fm DFF_P127(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2412));
DFF_save_fm DFF_P128(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2422));
DFF_save_fm DFF_P129(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2432));
DFF_save_fm DFF_P130(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2442));
DFF_save_fm DFF_P131(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2452));
DFF_save_fm DFF_P132(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2462));
DFF_save_fm DFF_P133(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2502));
DFF_save_fm DFF_P134(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2512));
DFF_save_fm DFF_P135(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2522));
DFF_save_fm DFF_P136(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2532));
DFF_save_fm DFF_P137(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2542));
DFF_save_fm DFF_P138(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2552));
DFF_save_fm DFF_P139(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2562));
DFF_save_fm DFF_P140(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2602));
DFF_save_fm DFF_P141(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2612));
DFF_save_fm DFF_P142(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2622));
DFF_save_fm DFF_P143(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2632));
DFF_save_fm DFF_P144(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2642));
DFF_save_fm DFF_P145(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2652));
DFF_save_fm DFF_P146(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2662));
DFF_save_fm DFF_P147(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2003));
DFF_save_fm DFF_P148(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2013));
DFF_save_fm DFF_P149(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2023));
DFF_save_fm DFF_P150(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2033));
DFF_save_fm DFF_P151(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2043));
DFF_save_fm DFF_P152(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2053));
DFF_save_fm DFF_P153(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2063));
DFF_save_fm DFF_P154(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2103));
DFF_save_fm DFF_P155(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2113));
DFF_save_fm DFF_P156(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2123));
DFF_save_fm DFF_P157(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2133));
DFF_save_fm DFF_P158(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2143));
DFF_save_fm DFF_P159(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2153));
DFF_save_fm DFF_P160(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2163));
DFF_save_fm DFF_P161(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2203));
DFF_save_fm DFF_P162(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2213));
DFF_save_fm DFF_P163(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2223));
DFF_save_fm DFF_P164(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2233));
DFF_save_fm DFF_P165(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2243));
DFF_save_fm DFF_P166(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2253));
DFF_save_fm DFF_P167(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2263));
DFF_save_fm DFF_P168(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2303));
DFF_save_fm DFF_P169(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2313));
DFF_save_fm DFF_P170(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2323));
DFF_save_fm DFF_P171(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2333));
DFF_save_fm DFF_P172(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2343));
DFF_save_fm DFF_P173(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2353));
DFF_save_fm DFF_P174(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2363));
DFF_save_fm DFF_P175(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2403));
DFF_save_fm DFF_P176(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2413));
DFF_save_fm DFF_P177(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2423));
DFF_save_fm DFF_P178(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2433));
DFF_save_fm DFF_P179(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2443));
DFF_save_fm DFF_P180(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2453));
DFF_save_fm DFF_P181(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2463));
DFF_save_fm DFF_P182(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2503));
DFF_save_fm DFF_P183(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2513));
DFF_save_fm DFF_P184(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2523));
DFF_save_fm DFF_P185(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2533));
DFF_save_fm DFF_P186(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2543));
DFF_save_fm DFF_P187(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2553));
DFF_save_fm DFF_P188(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2563));
DFF_save_fm DFF_P189(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2603));
DFF_save_fm DFF_P190(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2613));
DFF_save_fm DFF_P191(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2623));
DFF_save_fm DFF_P192(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2633));
DFF_save_fm DFF_P193(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2643));
DFF_save_fm DFF_P194(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2653));
DFF_save_fm DFF_P195(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2663));
DFF_save_fm DFF_P196(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2004));
DFF_save_fm DFF_P197(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2014));
DFF_save_fm DFF_P198(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2024));
DFF_save_fm DFF_P199(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2034));
DFF_save_fm DFF_P200(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2044));
DFF_save_fm DFF_P201(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2054));
DFF_save_fm DFF_P202(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2064));
DFF_save_fm DFF_P203(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2104));
DFF_save_fm DFF_P204(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2114));
DFF_save_fm DFF_P205(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2124));
DFF_save_fm DFF_P206(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2134));
DFF_save_fm DFF_P207(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2144));
DFF_save_fm DFF_P208(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2154));
DFF_save_fm DFF_P209(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2164));
DFF_save_fm DFF_P210(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2204));
DFF_save_fm DFF_P211(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2214));
DFF_save_fm DFF_P212(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2224));
DFF_save_fm DFF_P213(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2234));
DFF_save_fm DFF_P214(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2244));
DFF_save_fm DFF_P215(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2254));
DFF_save_fm DFF_P216(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2264));
DFF_save_fm DFF_P217(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2304));
DFF_save_fm DFF_P218(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2314));
DFF_save_fm DFF_P219(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2324));
DFF_save_fm DFF_P220(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2334));
DFF_save_fm DFF_P221(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2344));
DFF_save_fm DFF_P222(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2354));
DFF_save_fm DFF_P223(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2364));
DFF_save_fm DFF_P224(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2404));
DFF_save_fm DFF_P225(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2414));
DFF_save_fm DFF_P226(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2424));
DFF_save_fm DFF_P227(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2434));
DFF_save_fm DFF_P228(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2444));
DFF_save_fm DFF_P229(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2454));
DFF_save_fm DFF_P230(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2464));
DFF_save_fm DFF_P231(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2504));
DFF_save_fm DFF_P232(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2514));
DFF_save_fm DFF_P233(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2524));
DFF_save_fm DFF_P234(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2534));
DFF_save_fm DFF_P235(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2544));
DFF_save_fm DFF_P236(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2554));
DFF_save_fm DFF_P237(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2564));
DFF_save_fm DFF_P238(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2604));
DFF_save_fm DFF_P239(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2614));
DFF_save_fm DFF_P240(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2624));
DFF_save_fm DFF_P241(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2634));
DFF_save_fm DFF_P242(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2644));
DFF_save_fm DFF_P243(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2654));
DFF_save_fm DFF_P244(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2664));
DFF_save_fm DFF_P245(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2005));
DFF_save_fm DFF_P246(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2015));
DFF_save_fm DFF_P247(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2025));
DFF_save_fm DFF_P248(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2035));
DFF_save_fm DFF_P249(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2045));
DFF_save_fm DFF_P250(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2055));
DFF_save_fm DFF_P251(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2065));
DFF_save_fm DFF_P252(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2105));
DFF_save_fm DFF_P253(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2115));
DFF_save_fm DFF_P254(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2125));
DFF_save_fm DFF_P255(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2135));
DFF_save_fm DFF_P256(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2145));
DFF_save_fm DFF_P257(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2155));
DFF_save_fm DFF_P258(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2165));
DFF_save_fm DFF_P259(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2205));
DFF_save_fm DFF_P260(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2215));
DFF_save_fm DFF_P261(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2225));
DFF_save_fm DFF_P262(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2235));
DFF_save_fm DFF_P263(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2245));
DFF_save_fm DFF_P264(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2255));
DFF_save_fm DFF_P265(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2265));
DFF_save_fm DFF_P266(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2305));
DFF_save_fm DFF_P267(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2315));
DFF_save_fm DFF_P268(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2325));
DFF_save_fm DFF_P269(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2335));
DFF_save_fm DFF_P270(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2345));
DFF_save_fm DFF_P271(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2355));
DFF_save_fm DFF_P272(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2365));
DFF_save_fm DFF_P273(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2405));
DFF_save_fm DFF_P274(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2415));
DFF_save_fm DFF_P275(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2425));
DFF_save_fm DFF_P276(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2435));
DFF_save_fm DFF_P277(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2445));
DFF_save_fm DFF_P278(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2455));
DFF_save_fm DFF_P279(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2465));
DFF_save_fm DFF_P280(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2505));
DFF_save_fm DFF_P281(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2515));
DFF_save_fm DFF_P282(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2525));
DFF_save_fm DFF_P283(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2535));
DFF_save_fm DFF_P284(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2545));
DFF_save_fm DFF_P285(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2555));
DFF_save_fm DFF_P286(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2565));
DFF_save_fm DFF_P287(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2605));
DFF_save_fm DFF_P288(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2615));
DFF_save_fm DFF_P289(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2625));
DFF_save_fm DFF_P290(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2635));
DFF_save_fm DFF_P291(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2645));
DFF_save_fm DFF_P292(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2655));
DFF_save_fm DFF_P293(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2665));
DFF_save_fm DFF_P294(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2006));
DFF_save_fm DFF_P295(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2016));
DFF_save_fm DFF_P296(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2026));
DFF_save_fm DFF_P297(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2036));
DFF_save_fm DFF_P298(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2046));
DFF_save_fm DFF_P299(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2056));
DFF_save_fm DFF_P300(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2066));
DFF_save_fm DFF_P301(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2106));
DFF_save_fm DFF_P302(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2116));
DFF_save_fm DFF_P303(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2126));
DFF_save_fm DFF_P304(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2136));
DFF_save_fm DFF_P305(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2146));
DFF_save_fm DFF_P306(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2156));
DFF_save_fm DFF_P307(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2166));
DFF_save_fm DFF_P308(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2206));
DFF_save_fm DFF_P309(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2216));
DFF_save_fm DFF_P310(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2226));
DFF_save_fm DFF_P311(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2236));
DFF_save_fm DFF_P312(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2246));
DFF_save_fm DFF_P313(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2256));
DFF_save_fm DFF_P314(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2266));
DFF_save_fm DFF_P315(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2306));
DFF_save_fm DFF_P316(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2316));
DFF_save_fm DFF_P317(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2326));
DFF_save_fm DFF_P318(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2336));
DFF_save_fm DFF_P319(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2346));
DFF_save_fm DFF_P320(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2356));
DFF_save_fm DFF_P321(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2366));
DFF_save_fm DFF_P322(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2406));
DFF_save_fm DFF_P323(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2416));
DFF_save_fm DFF_P324(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2426));
DFF_save_fm DFF_P325(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2436));
DFF_save_fm DFF_P326(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2446));
DFF_save_fm DFF_P327(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2456));
DFF_save_fm DFF_P328(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2466));
DFF_save_fm DFF_P329(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2506));
DFF_save_fm DFF_P330(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2516));
DFF_save_fm DFF_P331(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2526));
DFF_save_fm DFF_P332(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2536));
DFF_save_fm DFF_P333(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2546));
DFF_save_fm DFF_P334(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2556));
DFF_save_fm DFF_P335(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2566));
DFF_save_fm DFF_P336(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2606));
DFF_save_fm DFF_P337(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2616));
DFF_save_fm DFF_P338(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2626));
DFF_save_fm DFF_P339(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2636));
DFF_save_fm DFF_P340(.clk(clk),.rstn(rstn),.reset_value(0),.q(P2646));
DFF_save_fm DFF_P341(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2656));
DFF_save_fm DFF_P342(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2666));
DFF_save_fm DFF_P343(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2007));
DFF_save_fm DFF_P344(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2017));
DFF_save_fm DFF_P345(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2027));
DFF_save_fm DFF_P346(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2037));
DFF_save_fm DFF_P347(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2047));
DFF_save_fm DFF_P348(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2057));
DFF_save_fm DFF_P349(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2067));
DFF_save_fm DFF_P350(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2107));
DFF_save_fm DFF_P351(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2117));
DFF_save_fm DFF_P352(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2127));
DFF_save_fm DFF_P353(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2137));
DFF_save_fm DFF_P354(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2147));
DFF_save_fm DFF_P355(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2157));
DFF_save_fm DFF_P356(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2167));
DFF_save_fm DFF_P357(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2207));
DFF_save_fm DFF_P358(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2217));
DFF_save_fm DFF_P359(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2227));
DFF_save_fm DFF_P360(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2237));
DFF_save_fm DFF_P361(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2247));
DFF_save_fm DFF_P362(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2257));
DFF_save_fm DFF_P363(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2267));
DFF_save_fm DFF_P364(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2307));
DFF_save_fm DFF_P365(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2317));
DFF_save_fm DFF_P366(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2327));
DFF_save_fm DFF_P367(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2337));
DFF_save_fm DFF_P368(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2347));
DFF_save_fm DFF_P369(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2357));
DFF_save_fm DFF_P370(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2367));
DFF_save_fm DFF_P371(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2407));
DFF_save_fm DFF_P372(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2417));
DFF_save_fm DFF_P373(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2427));
DFF_save_fm DFF_P374(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2437));
DFF_save_fm DFF_P375(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2447));
DFF_save_fm DFF_P376(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2457));
DFF_save_fm DFF_P377(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2467));
DFF_save_fm DFF_P378(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2507));
DFF_save_fm DFF_P379(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2517));
DFF_save_fm DFF_P380(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2527));
DFF_save_fm DFF_P381(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2537));
DFF_save_fm DFF_P382(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2547));
DFF_save_fm DFF_P383(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2557));
DFF_save_fm DFF_P384(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2567));
DFF_save_fm DFF_P385(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2607));
DFF_save_fm DFF_P386(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2617));
DFF_save_fm DFF_P387(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2627));
DFF_save_fm DFF_P388(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2637));
DFF_save_fm DFF_P389(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2647));
DFF_save_fm DFF_P390(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2657));
DFF_save_fm DFF_P391(.clk(clk),.rstn(rstn),.reset_value(1),.q(P2667));
DFF_save_fm DFF_W0(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20000));
DFF_save_fm DFF_W1(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20010));
DFF_save_fm DFF_W2(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20020));
DFF_save_fm DFF_W3(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20100));
DFF_save_fm DFF_W4(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20110));
DFF_save_fm DFF_W5(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20120));
DFF_save_fm DFF_W6(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20200));
DFF_save_fm DFF_W7(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20210));
DFF_save_fm DFF_W8(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20220));
DFF_save_fm DFF_W9(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20001));
DFF_save_fm DFF_W10(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20011));
DFF_save_fm DFF_W11(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20021));
DFF_save_fm DFF_W12(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20101));
DFF_save_fm DFF_W13(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20111));
DFF_save_fm DFF_W14(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20121));
DFF_save_fm DFF_W15(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20201));
DFF_save_fm DFF_W16(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20211));
DFF_save_fm DFF_W17(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20221));
DFF_save_fm DFF_W18(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20002));
DFF_save_fm DFF_W19(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20012));
DFF_save_fm DFF_W20(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20022));
DFF_save_fm DFF_W21(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20102));
DFF_save_fm DFF_W22(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20112));
DFF_save_fm DFF_W23(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20122));
DFF_save_fm DFF_W24(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20202));
DFF_save_fm DFF_W25(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20212));
DFF_save_fm DFF_W26(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20222));
DFF_save_fm DFF_W27(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20003));
DFF_save_fm DFF_W28(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20013));
DFF_save_fm DFF_W29(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20023));
DFF_save_fm DFF_W30(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20103));
DFF_save_fm DFF_W31(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20113));
DFF_save_fm DFF_W32(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20123));
DFF_save_fm DFF_W33(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20203));
DFF_save_fm DFF_W34(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20213));
DFF_save_fm DFF_W35(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20223));
DFF_save_fm DFF_W36(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20004));
DFF_save_fm DFF_W37(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20014));
DFF_save_fm DFF_W38(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20024));
DFF_save_fm DFF_W39(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20104));
DFF_save_fm DFF_W40(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20114));
DFF_save_fm DFF_W41(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20124));
DFF_save_fm DFF_W42(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20204));
DFF_save_fm DFF_W43(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20214));
DFF_save_fm DFF_W44(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20224));
DFF_save_fm DFF_W45(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20005));
DFF_save_fm DFF_W46(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20015));
DFF_save_fm DFF_W47(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20025));
DFF_save_fm DFF_W48(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20105));
DFF_save_fm DFF_W49(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20115));
DFF_save_fm DFF_W50(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20125));
DFF_save_fm DFF_W51(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20205));
DFF_save_fm DFF_W52(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20215));
DFF_save_fm DFF_W53(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20225));
DFF_save_fm DFF_W54(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20006));
DFF_save_fm DFF_W55(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20016));
DFF_save_fm DFF_W56(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20026));
DFF_save_fm DFF_W57(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20106));
DFF_save_fm DFF_W58(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20116));
DFF_save_fm DFF_W59(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20126));
DFF_save_fm DFF_W60(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20206));
DFF_save_fm DFF_W61(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20216));
DFF_save_fm DFF_W62(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20226));
DFF_save_fm DFF_W63(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20007));
DFF_save_fm DFF_W64(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20017));
DFF_save_fm DFF_W65(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20027));
DFF_save_fm DFF_W66(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20107));
DFF_save_fm DFF_W67(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20117));
DFF_save_fm DFF_W68(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20127));
DFF_save_fm DFF_W69(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20207));
DFF_save_fm DFF_W70(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20217));
DFF_save_fm DFF_W71(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20227));
DFF_save_fm DFF_W72(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21000));
DFF_save_fm DFF_W73(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21010));
DFF_save_fm DFF_W74(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21020));
DFF_save_fm DFF_W75(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21100));
DFF_save_fm DFF_W76(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21110));
DFF_save_fm DFF_W77(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21120));
DFF_save_fm DFF_W78(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21200));
DFF_save_fm DFF_W79(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21210));
DFF_save_fm DFF_W80(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21220));
DFF_save_fm DFF_W81(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21001));
DFF_save_fm DFF_W82(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21011));
DFF_save_fm DFF_W83(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21021));
DFF_save_fm DFF_W84(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21101));
DFF_save_fm DFF_W85(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21111));
DFF_save_fm DFF_W86(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21121));
DFF_save_fm DFF_W87(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21201));
DFF_save_fm DFF_W88(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21211));
DFF_save_fm DFF_W89(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21221));
DFF_save_fm DFF_W90(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21002));
DFF_save_fm DFF_W91(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21012));
DFF_save_fm DFF_W92(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21022));
DFF_save_fm DFF_W93(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21102));
DFF_save_fm DFF_W94(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21112));
DFF_save_fm DFF_W95(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21122));
DFF_save_fm DFF_W96(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21202));
DFF_save_fm DFF_W97(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21212));
DFF_save_fm DFF_W98(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21222));
DFF_save_fm DFF_W99(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21003));
DFF_save_fm DFF_W100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21013));
DFF_save_fm DFF_W101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21023));
DFF_save_fm DFF_W102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21103));
DFF_save_fm DFF_W103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21113));
DFF_save_fm DFF_W104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21123));
DFF_save_fm DFF_W105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21203));
DFF_save_fm DFF_W106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21213));
DFF_save_fm DFF_W107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21223));
DFF_save_fm DFF_W108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21004));
DFF_save_fm DFF_W109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21014));
DFF_save_fm DFF_W110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21024));
DFF_save_fm DFF_W111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21104));
DFF_save_fm DFF_W112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21114));
DFF_save_fm DFF_W113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21124));
DFF_save_fm DFF_W114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21204));
DFF_save_fm DFF_W115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21214));
DFF_save_fm DFF_W116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21224));
DFF_save_fm DFF_W117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21005));
DFF_save_fm DFF_W118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21015));
DFF_save_fm DFF_W119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21025));
DFF_save_fm DFF_W120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21105));
DFF_save_fm DFF_W121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21115));
DFF_save_fm DFF_W122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21125));
DFF_save_fm DFF_W123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21205));
DFF_save_fm DFF_W124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21215));
DFF_save_fm DFF_W125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21225));
DFF_save_fm DFF_W126(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21006));
DFF_save_fm DFF_W127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21016));
DFF_save_fm DFF_W128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21026));
DFF_save_fm DFF_W129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21106));
DFF_save_fm DFF_W130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21116));
DFF_save_fm DFF_W131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21126));
DFF_save_fm DFF_W132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21206));
DFF_save_fm DFF_W133(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21216));
DFF_save_fm DFF_W134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21226));
DFF_save_fm DFF_W135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21007));
DFF_save_fm DFF_W136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21017));
DFF_save_fm DFF_W137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21027));
DFF_save_fm DFF_W138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21107));
DFF_save_fm DFF_W139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21117));
DFF_save_fm DFF_W140(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21127));
DFF_save_fm DFF_W141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21207));
DFF_save_fm DFF_W142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21217));
DFF_save_fm DFF_W143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21227));
DFF_save_fm DFF_W144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22000));
DFF_save_fm DFF_W145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22010));
DFF_save_fm DFF_W146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22020));
DFF_save_fm DFF_W147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22100));
DFF_save_fm DFF_W148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22110));
DFF_save_fm DFF_W149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22120));
DFF_save_fm DFF_W150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22200));
DFF_save_fm DFF_W151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22210));
DFF_save_fm DFF_W152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22220));
DFF_save_fm DFF_W153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22001));
DFF_save_fm DFF_W154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22011));
DFF_save_fm DFF_W155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22021));
DFF_save_fm DFF_W156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22101));
DFF_save_fm DFF_W157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22111));
DFF_save_fm DFF_W158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22121));
DFF_save_fm DFF_W159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22201));
DFF_save_fm DFF_W160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22211));
DFF_save_fm DFF_W161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22221));
DFF_save_fm DFF_W162(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22002));
DFF_save_fm DFF_W163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22012));
DFF_save_fm DFF_W164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22022));
DFF_save_fm DFF_W165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22102));
DFF_save_fm DFF_W166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22112));
DFF_save_fm DFF_W167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22122));
DFF_save_fm DFF_W168(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22202));
DFF_save_fm DFF_W169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22212));
DFF_save_fm DFF_W170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22222));
DFF_save_fm DFF_W171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22003));
DFF_save_fm DFF_W172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22013));
DFF_save_fm DFF_W173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22023));
DFF_save_fm DFF_W174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22103));
DFF_save_fm DFF_W175(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22113));
DFF_save_fm DFF_W176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22123));
DFF_save_fm DFF_W177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22203));
DFF_save_fm DFF_W178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22213));
DFF_save_fm DFF_W179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22223));
DFF_save_fm DFF_W180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22004));
DFF_save_fm DFF_W181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22014));
DFF_save_fm DFF_W182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22024));
DFF_save_fm DFF_W183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22104));
DFF_save_fm DFF_W184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22114));
DFF_save_fm DFF_W185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22124));
DFF_save_fm DFF_W186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22204));
DFF_save_fm DFF_W187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22214));
DFF_save_fm DFF_W188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22224));
DFF_save_fm DFF_W189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22005));
DFF_save_fm DFF_W190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22015));
DFF_save_fm DFF_W191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22025));
DFF_save_fm DFF_W192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22105));
DFF_save_fm DFF_W193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22115));
DFF_save_fm DFF_W194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22125));
DFF_save_fm DFF_W195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22205));
DFF_save_fm DFF_W196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22215));
DFF_save_fm DFF_W197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22225));
DFF_save_fm DFF_W198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22006));
DFF_save_fm DFF_W199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22016));
DFF_save_fm DFF_W200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22026));
DFF_save_fm DFF_W201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22106));
DFF_save_fm DFF_W202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22116));
DFF_save_fm DFF_W203(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22126));
DFF_save_fm DFF_W204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22206));
DFF_save_fm DFF_W205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22216));
DFF_save_fm DFF_W206(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22226));
DFF_save_fm DFF_W207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22007));
DFF_save_fm DFF_W208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22017));
DFF_save_fm DFF_W209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22027));
DFF_save_fm DFF_W210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22107));
DFF_save_fm DFF_W211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22117));
DFF_save_fm DFF_W212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22127));
DFF_save_fm DFF_W213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22207));
DFF_save_fm DFF_W214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22217));
DFF_save_fm DFF_W215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22227));
DFF_save_fm DFF_W216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23000));
DFF_save_fm DFF_W217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23010));
DFF_save_fm DFF_W218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23020));
DFF_save_fm DFF_W219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23100));
DFF_save_fm DFF_W220(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23110));
DFF_save_fm DFF_W221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23120));
DFF_save_fm DFF_W222(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23200));
DFF_save_fm DFF_W223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23210));
DFF_save_fm DFF_W224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23220));
DFF_save_fm DFF_W225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23001));
DFF_save_fm DFF_W226(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23011));
DFF_save_fm DFF_W227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23021));
DFF_save_fm DFF_W228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23101));
DFF_save_fm DFF_W229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23111));
DFF_save_fm DFF_W230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23121));
DFF_save_fm DFF_W231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23201));
DFF_save_fm DFF_W232(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23211));
DFF_save_fm DFF_W233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23221));
DFF_save_fm DFF_W234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23002));
DFF_save_fm DFF_W235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23012));
DFF_save_fm DFF_W236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23022));
DFF_save_fm DFF_W237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23102));
DFF_save_fm DFF_W238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23112));
DFF_save_fm DFF_W239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23122));
DFF_save_fm DFF_W240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23202));
DFF_save_fm DFF_W241(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23212));
DFF_save_fm DFF_W242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23222));
DFF_save_fm DFF_W243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23003));
DFF_save_fm DFF_W244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23013));
DFF_save_fm DFF_W245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23023));
DFF_save_fm DFF_W246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23103));
DFF_save_fm DFF_W247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23113));
DFF_save_fm DFF_W248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23123));
DFF_save_fm DFF_W249(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23203));
DFF_save_fm DFF_W250(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23213));
DFF_save_fm DFF_W251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23223));
DFF_save_fm DFF_W252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23004));
DFF_save_fm DFF_W253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23014));
DFF_save_fm DFF_W254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23024));
DFF_save_fm DFF_W255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23104));
DFF_save_fm DFF_W256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23114));
DFF_save_fm DFF_W257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23124));
DFF_save_fm DFF_W258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23204));
DFF_save_fm DFF_W259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23214));
DFF_save_fm DFF_W260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23224));
DFF_save_fm DFF_W261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23005));
DFF_save_fm DFF_W262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23015));
DFF_save_fm DFF_W263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23025));
DFF_save_fm DFF_W264(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23105));
DFF_save_fm DFF_W265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23115));
DFF_save_fm DFF_W266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23125));
DFF_save_fm DFF_W267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23205));
DFF_save_fm DFF_W268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23215));
DFF_save_fm DFF_W269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23225));
DFF_save_fm DFF_W270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23006));
DFF_save_fm DFF_W271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23016));
DFF_save_fm DFF_W272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23026));
DFF_save_fm DFF_W273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23106));
DFF_save_fm DFF_W274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23116));
DFF_save_fm DFF_W275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23126));
DFF_save_fm DFF_W276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23206));
DFF_save_fm DFF_W277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23216));
DFF_save_fm DFF_W278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23226));
DFF_save_fm DFF_W279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23007));
DFF_save_fm DFF_W280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23017));
DFF_save_fm DFF_W281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23027));
DFF_save_fm DFF_W282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23107));
DFF_save_fm DFF_W283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23117));
DFF_save_fm DFF_W284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23127));
DFF_save_fm DFF_W285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23207));
DFF_save_fm DFF_W286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23217));
DFF_save_fm DFF_W287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23227));
DFF_save_fm DFF_W288(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24000));
DFF_save_fm DFF_W289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24010));
DFF_save_fm DFF_W290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24020));
DFF_save_fm DFF_W291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24100));
DFF_save_fm DFF_W292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24110));
DFF_save_fm DFF_W293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24120));
DFF_save_fm DFF_W294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24200));
DFF_save_fm DFF_W295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24210));
DFF_save_fm DFF_W296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24220));
DFF_save_fm DFF_W297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24001));
DFF_save_fm DFF_W298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24011));
DFF_save_fm DFF_W299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24021));
DFF_save_fm DFF_W300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24101));
DFF_save_fm DFF_W301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24111));
DFF_save_fm DFF_W302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24121));
DFF_save_fm DFF_W303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24201));
DFF_save_fm DFF_W304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24211));
DFF_save_fm DFF_W305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24221));
DFF_save_fm DFF_W306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24002));
DFF_save_fm DFF_W307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24012));
DFF_save_fm DFF_W308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24022));
DFF_save_fm DFF_W309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24102));
DFF_save_fm DFF_W310(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24112));
DFF_save_fm DFF_W311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24122));
DFF_save_fm DFF_W312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24202));
DFF_save_fm DFF_W313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24212));
DFF_save_fm DFF_W314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24222));
DFF_save_fm DFF_W315(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24003));
DFF_save_fm DFF_W316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24013));
DFF_save_fm DFF_W317(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24023));
DFF_save_fm DFF_W318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24103));
DFF_save_fm DFF_W319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24113));
DFF_save_fm DFF_W320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24123));
DFF_save_fm DFF_W321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24203));
DFF_save_fm DFF_W322(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24213));
DFF_save_fm DFF_W323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24223));
DFF_save_fm DFF_W324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24004));
DFF_save_fm DFF_W325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24014));
DFF_save_fm DFF_W326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24024));
DFF_save_fm DFF_W327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24104));
DFF_save_fm DFF_W328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24114));
DFF_save_fm DFF_W329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24124));
DFF_save_fm DFF_W330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24204));
DFF_save_fm DFF_W331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24214));
DFF_save_fm DFF_W332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24224));
DFF_save_fm DFF_W333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24005));
DFF_save_fm DFF_W334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24015));
DFF_save_fm DFF_W335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24025));
DFF_save_fm DFF_W336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24105));
DFF_save_fm DFF_W337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24115));
DFF_save_fm DFF_W338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24125));
DFF_save_fm DFF_W339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24205));
DFF_save_fm DFF_W340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24215));
DFF_save_fm DFF_W341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24225));
DFF_save_fm DFF_W342(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24006));
DFF_save_fm DFF_W343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24016));
DFF_save_fm DFF_W344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24026));
DFF_save_fm DFF_W345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24106));
DFF_save_fm DFF_W346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24116));
DFF_save_fm DFF_W347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24126));
DFF_save_fm DFF_W348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24206));
DFF_save_fm DFF_W349(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24216));
DFF_save_fm DFF_W350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24226));
DFF_save_fm DFF_W351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24007));
DFF_save_fm DFF_W352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24017));
DFF_save_fm DFF_W353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24027));
DFF_save_fm DFF_W354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24107));
DFF_save_fm DFF_W355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24117));
DFF_save_fm DFF_W356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24127));
DFF_save_fm DFF_W357(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24207));
DFF_save_fm DFF_W358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24217));
DFF_save_fm DFF_W359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24227));
DFF_save_fm DFF_W360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25000));
DFF_save_fm DFF_W361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25010));
DFF_save_fm DFF_W362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25020));
DFF_save_fm DFF_W363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25100));
DFF_save_fm DFF_W364(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25110));
DFF_save_fm DFF_W365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25120));
DFF_save_fm DFF_W366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25200));
DFF_save_fm DFF_W367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25210));
DFF_save_fm DFF_W368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25220));
DFF_save_fm DFF_W369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25001));
DFF_save_fm DFF_W370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25011));
DFF_save_fm DFF_W371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25021));
DFF_save_fm DFF_W372(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25101));
DFF_save_fm DFF_W373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25111));
DFF_save_fm DFF_W374(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25121));
DFF_save_fm DFF_W375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25201));
DFF_save_fm DFF_W376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25211));
DFF_save_fm DFF_W377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25221));
DFF_save_fm DFF_W378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25002));
DFF_save_fm DFF_W379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25012));
DFF_save_fm DFF_W380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25022));
DFF_save_fm DFF_W381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25102));
DFF_save_fm DFF_W382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25112));
DFF_save_fm DFF_W383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25122));
DFF_save_fm DFF_W384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25202));
DFF_save_fm DFF_W385(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25212));
DFF_save_fm DFF_W386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25222));
DFF_save_fm DFF_W387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25003));
DFF_save_fm DFF_W388(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25013));
DFF_save_fm DFF_W389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25023));
DFF_save_fm DFF_W390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25103));
DFF_save_fm DFF_W391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25113));
DFF_save_fm DFF_W392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25123));
DFF_save_fm DFF_W393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25203));
DFF_save_fm DFF_W394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25213));
DFF_save_fm DFF_W395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25223));
DFF_save_fm DFF_W396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25004));
DFF_save_fm DFF_W397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25014));
DFF_save_fm DFF_W398(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25024));
DFF_save_fm DFF_W399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25104));
DFF_save_fm DFF_W400(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25114));
DFF_save_fm DFF_W401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25124));
DFF_save_fm DFF_W402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25204));
DFF_save_fm DFF_W403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25214));
DFF_save_fm DFF_W404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25224));
DFF_save_fm DFF_W405(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25005));
DFF_save_fm DFF_W406(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25015));
DFF_save_fm DFF_W407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25025));
DFF_save_fm DFF_W408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25105));
DFF_save_fm DFF_W409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25115));
DFF_save_fm DFF_W410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25125));
DFF_save_fm DFF_W411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25205));
DFF_save_fm DFF_W412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25215));
DFF_save_fm DFF_W413(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25225));
DFF_save_fm DFF_W414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25006));
DFF_save_fm DFF_W415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25016));
DFF_save_fm DFF_W416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25026));
DFF_save_fm DFF_W417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25106));
DFF_save_fm DFF_W418(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25116));
DFF_save_fm DFF_W419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25126));
DFF_save_fm DFF_W420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25206));
DFF_save_fm DFF_W421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25216));
DFF_save_fm DFF_W422(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25226));
DFF_save_fm DFF_W423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25007));
DFF_save_fm DFF_W424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25017));
DFF_save_fm DFF_W425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25027));
DFF_save_fm DFF_W426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25107));
DFF_save_fm DFF_W427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25117));
DFF_save_fm DFF_W428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25127));
DFF_save_fm DFF_W429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25207));
DFF_save_fm DFF_W430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25217));
DFF_save_fm DFF_W431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25227));
DFF_save_fm DFF_W432(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26000));
DFF_save_fm DFF_W433(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26010));
DFF_save_fm DFF_W434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26020));
DFF_save_fm DFF_W435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26100));
DFF_save_fm DFF_W436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26110));
DFF_save_fm DFF_W437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26120));
DFF_save_fm DFF_W438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26200));
DFF_save_fm DFF_W439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26210));
DFF_save_fm DFF_W440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26220));
DFF_save_fm DFF_W441(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26001));
DFF_save_fm DFF_W442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26011));
DFF_save_fm DFF_W443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26021));
DFF_save_fm DFF_W444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26101));
DFF_save_fm DFF_W445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26111));
DFF_save_fm DFF_W446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26121));
DFF_save_fm DFF_W447(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26201));
DFF_save_fm DFF_W448(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26211));
DFF_save_fm DFF_W449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26221));
DFF_save_fm DFF_W450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26002));
DFF_save_fm DFF_W451(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26012));
DFF_save_fm DFF_W452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26022));
DFF_save_fm DFF_W453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26102));
DFF_save_fm DFF_W454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26112));
DFF_save_fm DFF_W455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26122));
DFF_save_fm DFF_W456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26202));
DFF_save_fm DFF_W457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26212));
DFF_save_fm DFF_W458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26222));
DFF_save_fm DFF_W459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26003));
DFF_save_fm DFF_W460(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26013));
DFF_save_fm DFF_W461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26023));
DFF_save_fm DFF_W462(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26103));
DFF_save_fm DFF_W463(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26113));
DFF_save_fm DFF_W464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26123));
DFF_save_fm DFF_W465(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26203));
DFF_save_fm DFF_W466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26213));
DFF_save_fm DFF_W467(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26223));
DFF_save_fm DFF_W468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26004));
DFF_save_fm DFF_W469(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26014));
DFF_save_fm DFF_W470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26024));
DFF_save_fm DFF_W471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26104));
DFF_save_fm DFF_W472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26114));
DFF_save_fm DFF_W473(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26124));
DFF_save_fm DFF_W474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26204));
DFF_save_fm DFF_W475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26214));
DFF_save_fm DFF_W476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26224));
DFF_save_fm DFF_W477(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26005));
DFF_save_fm DFF_W478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26015));
DFF_save_fm DFF_W479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26025));
DFF_save_fm DFF_W480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26105));
DFF_save_fm DFF_W481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26115));
DFF_save_fm DFF_W482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26125));
DFF_save_fm DFF_W483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26205));
DFF_save_fm DFF_W484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26215));
DFF_save_fm DFF_W485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26225));
DFF_save_fm DFF_W486(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26006));
DFF_save_fm DFF_W487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26016));
DFF_save_fm DFF_W488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26026));
DFF_save_fm DFF_W489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26106));
DFF_save_fm DFF_W490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26116));
DFF_save_fm DFF_W491(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26126));
DFF_save_fm DFF_W492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26206));
DFF_save_fm DFF_W493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26216));
DFF_save_fm DFF_W494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26226));
DFF_save_fm DFF_W495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26007));
DFF_save_fm DFF_W496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26017));
DFF_save_fm DFF_W497(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26027));
DFF_save_fm DFF_W498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26107));
DFF_save_fm DFF_W499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26117));
DFF_save_fm DFF_W500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26127));
DFF_save_fm DFF_W501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26207));
DFF_save_fm DFF_W502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26217));
DFF_save_fm DFF_W503(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26227));
DFF_save_fm DFF_W504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27000));
DFF_save_fm DFF_W505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27010));
DFF_save_fm DFF_W506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27020));
DFF_save_fm DFF_W507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27100));
DFF_save_fm DFF_W508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27110));
DFF_save_fm DFF_W509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27120));
DFF_save_fm DFF_W510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27200));
DFF_save_fm DFF_W511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27210));
DFF_save_fm DFF_W512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27220));
DFF_save_fm DFF_W513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27001));
DFF_save_fm DFF_W514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27011));
DFF_save_fm DFF_W515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27021));
DFF_save_fm DFF_W516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27101));
DFF_save_fm DFF_W517(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27111));
DFF_save_fm DFF_W518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27121));
DFF_save_fm DFF_W519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27201));
DFF_save_fm DFF_W520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27211));
DFF_save_fm DFF_W521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27221));
DFF_save_fm DFF_W522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27002));
DFF_save_fm DFF_W523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27012));
DFF_save_fm DFF_W524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27022));
DFF_save_fm DFF_W525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27102));
DFF_save_fm DFF_W526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27112));
DFF_save_fm DFF_W527(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27122));
DFF_save_fm DFF_W528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27202));
DFF_save_fm DFF_W529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27212));
DFF_save_fm DFF_W530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27222));
DFF_save_fm DFF_W531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27003));
DFF_save_fm DFF_W532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27013));
DFF_save_fm DFF_W533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27023));
DFF_save_fm DFF_W534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27103));
DFF_save_fm DFF_W535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27113));
DFF_save_fm DFF_W536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27123));
DFF_save_fm DFF_W537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27203));
DFF_save_fm DFF_W538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27213));
DFF_save_fm DFF_W539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27223));
DFF_save_fm DFF_W540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27004));
DFF_save_fm DFF_W541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27014));
DFF_save_fm DFF_W542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27024));
DFF_save_fm DFF_W543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27104));
DFF_save_fm DFF_W544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27114));
DFF_save_fm DFF_W545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27124));
DFF_save_fm DFF_W546(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27204));
DFF_save_fm DFF_W547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27214));
DFF_save_fm DFF_W548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27224));
DFF_save_fm DFF_W549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27005));
DFF_save_fm DFF_W550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27015));
DFF_save_fm DFF_W551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27025));
DFF_save_fm DFF_W552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27105));
DFF_save_fm DFF_W553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27115));
DFF_save_fm DFF_W554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27125));
DFF_save_fm DFF_W555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27205));
DFF_save_fm DFF_W556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27215));
DFF_save_fm DFF_W557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27225));
DFF_save_fm DFF_W558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27006));
DFF_save_fm DFF_W559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27016));
DFF_save_fm DFF_W560(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27026));
DFF_save_fm DFF_W561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27106));
DFF_save_fm DFF_W562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27116));
DFF_save_fm DFF_W563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27126));
DFF_save_fm DFF_W564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27206));
DFF_save_fm DFF_W565(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27216));
DFF_save_fm DFF_W566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27226));
DFF_save_fm DFF_W567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27007));
DFF_save_fm DFF_W568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27017));
DFF_save_fm DFF_W569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27027));
DFF_save_fm DFF_W570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27107));
DFF_save_fm DFF_W571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27117));
DFF_save_fm DFF_W572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27127));
DFF_save_fm DFF_W573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27207));
DFF_save_fm DFF_W574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27217));
DFF_save_fm DFF_W575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27227));
DFF_save_fm DFF_W576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28000));
DFF_save_fm DFF_W577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28010));
DFF_save_fm DFF_W578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28020));
DFF_save_fm DFF_W579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28100));
DFF_save_fm DFF_W580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28110));
DFF_save_fm DFF_W581(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28120));
DFF_save_fm DFF_W582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28200));
DFF_save_fm DFF_W583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28210));
DFF_save_fm DFF_W584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28220));
DFF_save_fm DFF_W585(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28001));
DFF_save_fm DFF_W586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28011));
DFF_save_fm DFF_W587(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28021));
DFF_save_fm DFF_W588(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28101));
DFF_save_fm DFF_W589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28111));
DFF_save_fm DFF_W590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28121));
DFF_save_fm DFF_W591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28201));
DFF_save_fm DFF_W592(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28211));
DFF_save_fm DFF_W593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28221));
DFF_save_fm DFF_W594(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28002));
DFF_save_fm DFF_W595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28012));
DFF_save_fm DFF_W596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28022));
DFF_save_fm DFF_W597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28102));
DFF_save_fm DFF_W598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28112));
DFF_save_fm DFF_W599(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28122));
DFF_save_fm DFF_W600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28202));
DFF_save_fm DFF_W601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28212));
DFF_save_fm DFF_W602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28222));
DFF_save_fm DFF_W603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28003));
DFF_save_fm DFF_W604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28013));
DFF_save_fm DFF_W605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28023));
DFF_save_fm DFF_W606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28103));
DFF_save_fm DFF_W607(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28113));
DFF_save_fm DFF_W608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28123));
DFF_save_fm DFF_W609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28203));
DFF_save_fm DFF_W610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28213));
DFF_save_fm DFF_W611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28223));
DFF_save_fm DFF_W612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28004));
DFF_save_fm DFF_W613(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28014));
DFF_save_fm DFF_W614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28024));
DFF_save_fm DFF_W615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28104));
DFF_save_fm DFF_W616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28114));
DFF_save_fm DFF_W617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28124));
DFF_save_fm DFF_W618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28204));
DFF_save_fm DFF_W619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28214));
DFF_save_fm DFF_W620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28224));
DFF_save_fm DFF_W621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28005));
DFF_save_fm DFF_W622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28015));
DFF_save_fm DFF_W623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28025));
DFF_save_fm DFF_W624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28105));
DFF_save_fm DFF_W625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28115));
DFF_save_fm DFF_W626(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28125));
DFF_save_fm DFF_W627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28205));
DFF_save_fm DFF_W628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28215));
DFF_save_fm DFF_W629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28225));
DFF_save_fm DFF_W630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28006));
DFF_save_fm DFF_W631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28016));
DFF_save_fm DFF_W632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28026));
DFF_save_fm DFF_W633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28106));
DFF_save_fm DFF_W634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28116));
DFF_save_fm DFF_W635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28126));
DFF_save_fm DFF_W636(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28206));
DFF_save_fm DFF_W637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28216));
DFF_save_fm DFF_W638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28226));
DFF_save_fm DFF_W639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28007));
DFF_save_fm DFF_W640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28017));
DFF_save_fm DFF_W641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28027));
DFF_save_fm DFF_W642(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28107));
DFF_save_fm DFF_W643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28117));
DFF_save_fm DFF_W644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28127));
DFF_save_fm DFF_W645(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28207));
DFF_save_fm DFF_W646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28217));
DFF_save_fm DFF_W647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28227));
DFF_save_fm DFF_W648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29000));
DFF_save_fm DFF_W649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29010));
DFF_save_fm DFF_W650(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29020));
DFF_save_fm DFF_W651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29100));
DFF_save_fm DFF_W652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29110));
DFF_save_fm DFF_W653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29120));
DFF_save_fm DFF_W654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29200));
DFF_save_fm DFF_W655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29210));
DFF_save_fm DFF_W656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29220));
DFF_save_fm DFF_W657(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29001));
DFF_save_fm DFF_W658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29011));
DFF_save_fm DFF_W659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29021));
DFF_save_fm DFF_W660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29101));
DFF_save_fm DFF_W661(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29111));
DFF_save_fm DFF_W662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29121));
DFF_save_fm DFF_W663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29201));
DFF_save_fm DFF_W664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29211));
DFF_save_fm DFF_W665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29221));
DFF_save_fm DFF_W666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29002));
DFF_save_fm DFF_W667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29012));
DFF_save_fm DFF_W668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29022));
DFF_save_fm DFF_W669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29102));
DFF_save_fm DFF_W670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29112));
DFF_save_fm DFF_W671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29122));
DFF_save_fm DFF_W672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29202));
DFF_save_fm DFF_W673(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29212));
DFF_save_fm DFF_W674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29222));
DFF_save_fm DFF_W675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29003));
DFF_save_fm DFF_W676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29013));
DFF_save_fm DFF_W677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29023));
DFF_save_fm DFF_W678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29103));
DFF_save_fm DFF_W679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29113));
DFF_save_fm DFF_W680(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29123));
DFF_save_fm DFF_W681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29203));
DFF_save_fm DFF_W682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29213));
DFF_save_fm DFF_W683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29223));
DFF_save_fm DFF_W684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29004));
DFF_save_fm DFF_W685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29014));
DFF_save_fm DFF_W686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29024));
DFF_save_fm DFF_W687(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29104));
DFF_save_fm DFF_W688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29114));
DFF_save_fm DFF_W689(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29124));
DFF_save_fm DFF_W690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29204));
DFF_save_fm DFF_W691(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29214));
DFF_save_fm DFF_W692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29224));
DFF_save_fm DFF_W693(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29005));
DFF_save_fm DFF_W694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29015));
DFF_save_fm DFF_W695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29025));
DFF_save_fm DFF_W696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29105));
DFF_save_fm DFF_W697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29115));
DFF_save_fm DFF_W698(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29125));
DFF_save_fm DFF_W699(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29205));
DFF_save_fm DFF_W700(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29215));
DFF_save_fm DFF_W701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29225));
DFF_save_fm DFF_W702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29006));
DFF_save_fm DFF_W703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29016));
DFF_save_fm DFF_W704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29026));
DFF_save_fm DFF_W705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29106));
DFF_save_fm DFF_W706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29116));
DFF_save_fm DFF_W707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29126));
DFF_save_fm DFF_W708(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29206));
DFF_save_fm DFF_W709(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29216));
DFF_save_fm DFF_W710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29226));
DFF_save_fm DFF_W711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29007));
DFF_save_fm DFF_W712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29017));
DFF_save_fm DFF_W713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29027));
DFF_save_fm DFF_W714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29107));
DFF_save_fm DFF_W715(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29117));
DFF_save_fm DFF_W716(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29127));
DFF_save_fm DFF_W717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29207));
DFF_save_fm DFF_W718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29217));
DFF_save_fm DFF_W719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29227));
DFF_save_fm DFF_W720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A000));
DFF_save_fm DFF_W721(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A010));
DFF_save_fm DFF_W722(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A020));
DFF_save_fm DFF_W723(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A100));
DFF_save_fm DFF_W724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A110));
DFF_save_fm DFF_W725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A120));
DFF_save_fm DFF_W726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A200));
DFF_save_fm DFF_W727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A210));
DFF_save_fm DFF_W728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A220));
DFF_save_fm DFF_W729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A001));
DFF_save_fm DFF_W730(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A011));
DFF_save_fm DFF_W731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A021));
DFF_save_fm DFF_W732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A101));
DFF_save_fm DFF_W733(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A111));
DFF_save_fm DFF_W734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A121));
DFF_save_fm DFF_W735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A201));
DFF_save_fm DFF_W736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A211));
DFF_save_fm DFF_W737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A221));
DFF_save_fm DFF_W738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A002));
DFF_save_fm DFF_W739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A012));
DFF_save_fm DFF_W740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A022));
DFF_save_fm DFF_W741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A102));
DFF_save_fm DFF_W742(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A112));
DFF_save_fm DFF_W743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A122));
DFF_save_fm DFF_W744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A202));
DFF_save_fm DFF_W745(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A212));
DFF_save_fm DFF_W746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A222));
DFF_save_fm DFF_W747(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A003));
DFF_save_fm DFF_W748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A013));
DFF_save_fm DFF_W749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A023));
DFF_save_fm DFF_W750(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A103));
DFF_save_fm DFF_W751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A113));
DFF_save_fm DFF_W752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A123));
DFF_save_fm DFF_W753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A203));
DFF_save_fm DFF_W754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A213));
DFF_save_fm DFF_W755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A223));
DFF_save_fm DFF_W756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A004));
DFF_save_fm DFF_W757(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A014));
DFF_save_fm DFF_W758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A024));
DFF_save_fm DFF_W759(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A104));
DFF_save_fm DFF_W760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A114));
DFF_save_fm DFF_W761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A124));
DFF_save_fm DFF_W762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A204));
DFF_save_fm DFF_W763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A214));
DFF_save_fm DFF_W764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A224));
DFF_save_fm DFF_W765(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A005));
DFF_save_fm DFF_W766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A015));
DFF_save_fm DFF_W767(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A025));
DFF_save_fm DFF_W768(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A105));
DFF_save_fm DFF_W769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A115));
DFF_save_fm DFF_W770(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A125));
DFF_save_fm DFF_W771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A205));
DFF_save_fm DFF_W772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A215));
DFF_save_fm DFF_W773(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A225));
DFF_save_fm DFF_W774(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A006));
DFF_save_fm DFF_W775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A016));
DFF_save_fm DFF_W776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A026));
DFF_save_fm DFF_W777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A106));
DFF_save_fm DFF_W778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A116));
DFF_save_fm DFF_W779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A126));
DFF_save_fm DFF_W780(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A206));
DFF_save_fm DFF_W781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A216));
DFF_save_fm DFF_W782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A226));
DFF_save_fm DFF_W783(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A007));
DFF_save_fm DFF_W784(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A017));
DFF_save_fm DFF_W785(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A027));
DFF_save_fm DFF_W786(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A107));
DFF_save_fm DFF_W787(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A117));
DFF_save_fm DFF_W788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A127));
DFF_save_fm DFF_W789(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A207));
DFF_save_fm DFF_W790(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A217));
DFF_save_fm DFF_W791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A227));
DFF_save_fm DFF_W792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B000));
DFF_save_fm DFF_W793(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B010));
DFF_save_fm DFF_W794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B020));
DFF_save_fm DFF_W795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B100));
DFF_save_fm DFF_W796(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B110));
DFF_save_fm DFF_W797(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B120));
DFF_save_fm DFF_W798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B200));
DFF_save_fm DFF_W799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B210));
DFF_save_fm DFF_W800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B220));
DFF_save_fm DFF_W801(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B001));
DFF_save_fm DFF_W802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B011));
DFF_save_fm DFF_W803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B021));
DFF_save_fm DFF_W804(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B101));
DFF_save_fm DFF_W805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B111));
DFF_save_fm DFF_W806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B121));
DFF_save_fm DFF_W807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B201));
DFF_save_fm DFF_W808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B211));
DFF_save_fm DFF_W809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B221));
DFF_save_fm DFF_W810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B002));
DFF_save_fm DFF_W811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B012));
DFF_save_fm DFF_W812(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B022));
DFF_save_fm DFF_W813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B102));
DFF_save_fm DFF_W814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B112));
DFF_save_fm DFF_W815(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B122));
DFF_save_fm DFF_W816(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B202));
DFF_save_fm DFF_W817(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B212));
DFF_save_fm DFF_W818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B222));
DFF_save_fm DFF_W819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B003));
DFF_save_fm DFF_W820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B013));
DFF_save_fm DFF_W821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B023));
DFF_save_fm DFF_W822(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B103));
DFF_save_fm DFF_W823(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B113));
DFF_save_fm DFF_W824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B123));
DFF_save_fm DFF_W825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B203));
DFF_save_fm DFF_W826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B213));
DFF_save_fm DFF_W827(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B223));
DFF_save_fm DFF_W828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B004));
DFF_save_fm DFF_W829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B014));
DFF_save_fm DFF_W830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B024));
DFF_save_fm DFF_W831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B104));
DFF_save_fm DFF_W832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B114));
DFF_save_fm DFF_W833(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B124));
DFF_save_fm DFF_W834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B204));
DFF_save_fm DFF_W835(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B214));
DFF_save_fm DFF_W836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B224));
DFF_save_fm DFF_W837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B005));
DFF_save_fm DFF_W838(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B015));
DFF_save_fm DFF_W839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B025));
DFF_save_fm DFF_W840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B105));
DFF_save_fm DFF_W841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B115));
DFF_save_fm DFF_W842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B125));
DFF_save_fm DFF_W843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B205));
DFF_save_fm DFF_W844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B215));
DFF_save_fm DFF_W845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B225));
DFF_save_fm DFF_W846(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B006));
DFF_save_fm DFF_W847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B016));
DFF_save_fm DFF_W848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B026));
DFF_save_fm DFF_W849(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B106));
DFF_save_fm DFF_W850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B116));
DFF_save_fm DFF_W851(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B126));
DFF_save_fm DFF_W852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B206));
DFF_save_fm DFF_W853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B216));
DFF_save_fm DFF_W854(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B226));
DFF_save_fm DFF_W855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B007));
DFF_save_fm DFF_W856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B017));
DFF_save_fm DFF_W857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B027));
DFF_save_fm DFF_W858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B107));
DFF_save_fm DFF_W859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B117));
DFF_save_fm DFF_W860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B127));
DFF_save_fm DFF_W861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B207));
DFF_save_fm DFF_W862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B217));
DFF_save_fm DFF_W863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B227));
DFF_save_fm DFF_W864(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C000));
DFF_save_fm DFF_W865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C010));
DFF_save_fm DFF_W866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C020));
DFF_save_fm DFF_W867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C100));
DFF_save_fm DFF_W868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C110));
DFF_save_fm DFF_W869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C120));
DFF_save_fm DFF_W870(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C200));
DFF_save_fm DFF_W871(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C210));
DFF_save_fm DFF_W872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C220));
DFF_save_fm DFF_W873(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C001));
DFF_save_fm DFF_W874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C011));
DFF_save_fm DFF_W875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C021));
DFF_save_fm DFF_W876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C101));
DFF_save_fm DFF_W877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C111));
DFF_save_fm DFF_W878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C121));
DFF_save_fm DFF_W879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C201));
DFF_save_fm DFF_W880(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C211));
DFF_save_fm DFF_W881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C221));
DFF_save_fm DFF_W882(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C002));
DFF_save_fm DFF_W883(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C012));
DFF_save_fm DFF_W884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C022));
DFF_save_fm DFF_W885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C102));
DFF_save_fm DFF_W886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C112));
DFF_save_fm DFF_W887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C122));
DFF_save_fm DFF_W888(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C202));
DFF_save_fm DFF_W889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C212));
DFF_save_fm DFF_W890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C222));
DFF_save_fm DFF_W891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C003));
DFF_save_fm DFF_W892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C013));
DFF_save_fm DFF_W893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C023));
DFF_save_fm DFF_W894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C103));
DFF_save_fm DFF_W895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C113));
DFF_save_fm DFF_W896(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C123));
DFF_save_fm DFF_W897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C203));
DFF_save_fm DFF_W898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C213));
DFF_save_fm DFF_W899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C223));
DFF_save_fm DFF_W900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C004));
DFF_save_fm DFF_W901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C014));
DFF_save_fm DFF_W902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C024));
DFF_save_fm DFF_W903(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C104));
DFF_save_fm DFF_W904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C114));
DFF_save_fm DFF_W905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C124));
DFF_save_fm DFF_W906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C204));
DFF_save_fm DFF_W907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C214));
DFF_save_fm DFF_W908(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C224));
DFF_save_fm DFF_W909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C005));
DFF_save_fm DFF_W910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C015));
DFF_save_fm DFF_W911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C025));
DFF_save_fm DFF_W912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C105));
DFF_save_fm DFF_W913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C115));
DFF_save_fm DFF_W914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C125));
DFF_save_fm DFF_W915(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C205));
DFF_save_fm DFF_W916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C215));
DFF_save_fm DFF_W917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C225));
DFF_save_fm DFF_W918(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C006));
DFF_save_fm DFF_W919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C016));
DFF_save_fm DFF_W920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C026));
DFF_save_fm DFF_W921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C106));
DFF_save_fm DFF_W922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C116));
DFF_save_fm DFF_W923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C126));
DFF_save_fm DFF_W924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C206));
DFF_save_fm DFF_W925(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C216));
DFF_save_fm DFF_W926(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C226));
DFF_save_fm DFF_W927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C007));
DFF_save_fm DFF_W928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C017));
DFF_save_fm DFF_W929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C027));
DFF_save_fm DFF_W930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C107));
DFF_save_fm DFF_W931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C117));
DFF_save_fm DFF_W932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C127));
DFF_save_fm DFF_W933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C207));
DFF_save_fm DFF_W934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C217));
DFF_save_fm DFF_W935(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C227));
DFF_save_fm DFF_W936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D000));
DFF_save_fm DFF_W937(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D010));
DFF_save_fm DFF_W938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D020));
DFF_save_fm DFF_W939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D100));
DFF_save_fm DFF_W940(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D110));
DFF_save_fm DFF_W941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D120));
DFF_save_fm DFF_W942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D200));
DFF_save_fm DFF_W943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D210));
DFF_save_fm DFF_W944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D220));
DFF_save_fm DFF_W945(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D001));
DFF_save_fm DFF_W946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D011));
DFF_save_fm DFF_W947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D021));
DFF_save_fm DFF_W948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D101));
DFF_save_fm DFF_W949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D111));
DFF_save_fm DFF_W950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D121));
DFF_save_fm DFF_W951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D201));
DFF_save_fm DFF_W952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D211));
DFF_save_fm DFF_W953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D221));
DFF_save_fm DFF_W954(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D002));
DFF_save_fm DFF_W955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D012));
DFF_save_fm DFF_W956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D022));
DFF_save_fm DFF_W957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D102));
DFF_save_fm DFF_W958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D112));
DFF_save_fm DFF_W959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D122));
DFF_save_fm DFF_W960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D202));
DFF_save_fm DFF_W961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D212));
DFF_save_fm DFF_W962(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D222));
DFF_save_fm DFF_W963(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D003));
DFF_save_fm DFF_W964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D013));
DFF_save_fm DFF_W965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D023));
DFF_save_fm DFF_W966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D103));
DFF_save_fm DFF_W967(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D113));
DFF_save_fm DFF_W968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D123));
DFF_save_fm DFF_W969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D203));
DFF_save_fm DFF_W970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D213));
DFF_save_fm DFF_W971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D223));
DFF_save_fm DFF_W972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D004));
DFF_save_fm DFF_W973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D014));
DFF_save_fm DFF_W974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D024));
DFF_save_fm DFF_W975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D104));
DFF_save_fm DFF_W976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D114));
DFF_save_fm DFF_W977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D124));
DFF_save_fm DFF_W978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D204));
DFF_save_fm DFF_W979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D214));
DFF_save_fm DFF_W980(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D224));
DFF_save_fm DFF_W981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D005));
DFF_save_fm DFF_W982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D015));
DFF_save_fm DFF_W983(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D025));
DFF_save_fm DFF_W984(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D105));
DFF_save_fm DFF_W985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D115));
DFF_save_fm DFF_W986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D125));
DFF_save_fm DFF_W987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D205));
DFF_save_fm DFF_W988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D215));
DFF_save_fm DFF_W989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D225));
DFF_save_fm DFF_W990(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D006));
DFF_save_fm DFF_W991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D016));
DFF_save_fm DFF_W992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D026));
DFF_save_fm DFF_W993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D106));
DFF_save_fm DFF_W994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D116));
DFF_save_fm DFF_W995(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D126));
DFF_save_fm DFF_W996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D206));
DFF_save_fm DFF_W997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D216));
DFF_save_fm DFF_W998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D226));
DFF_save_fm DFF_W999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D007));
DFF_save_fm DFF_W1000(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D017));
DFF_save_fm DFF_W1001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D027));
DFF_save_fm DFF_W1002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D107));
DFF_save_fm DFF_W1003(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D117));
DFF_save_fm DFF_W1004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D127));
DFF_save_fm DFF_W1005(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D207));
DFF_save_fm DFF_W1006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D217));
DFF_save_fm DFF_W1007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D227));
DFF_save_fm DFF_W1008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E000));
DFF_save_fm DFF_W1009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E010));
DFF_save_fm DFF_W1010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E020));
DFF_save_fm DFF_W1011(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E100));
DFF_save_fm DFF_W1012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E110));
DFF_save_fm DFF_W1013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E120));
DFF_save_fm DFF_W1014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E200));
DFF_save_fm DFF_W1015(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E210));
DFF_save_fm DFF_W1016(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E220));
DFF_save_fm DFF_W1017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E001));
DFF_save_fm DFF_W1018(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E011));
DFF_save_fm DFF_W1019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E021));
DFF_save_fm DFF_W1020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E101));
DFF_save_fm DFF_W1021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E111));
DFF_save_fm DFF_W1022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E121));
DFF_save_fm DFF_W1023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E201));
DFF_save_fm DFF_W1024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E211));
DFF_save_fm DFF_W1025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E221));
DFF_save_fm DFF_W1026(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E002));
DFF_save_fm DFF_W1027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E012));
DFF_save_fm DFF_W1028(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E022));
DFF_save_fm DFF_W1029(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E102));
DFF_save_fm DFF_W1030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E112));
DFF_save_fm DFF_W1031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E122));
DFF_save_fm DFF_W1032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E202));
DFF_save_fm DFF_W1033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E212));
DFF_save_fm DFF_W1034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E222));
DFF_save_fm DFF_W1035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E003));
DFF_save_fm DFF_W1036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E013));
DFF_save_fm DFF_W1037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E023));
DFF_save_fm DFF_W1038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E103));
DFF_save_fm DFF_W1039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E113));
DFF_save_fm DFF_W1040(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E123));
DFF_save_fm DFF_W1041(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E203));
DFF_save_fm DFF_W1042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E213));
DFF_save_fm DFF_W1043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E223));
DFF_save_fm DFF_W1044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E004));
DFF_save_fm DFF_W1045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E014));
DFF_save_fm DFF_W1046(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E024));
DFF_save_fm DFF_W1047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E104));
DFF_save_fm DFF_W1048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E114));
DFF_save_fm DFF_W1049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E124));
DFF_save_fm DFF_W1050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E204));
DFF_save_fm DFF_W1051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E214));
DFF_save_fm DFF_W1052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E224));
DFF_save_fm DFF_W1053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E005));
DFF_save_fm DFF_W1054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E015));
DFF_save_fm DFF_W1055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E025));
DFF_save_fm DFF_W1056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E105));
DFF_save_fm DFF_W1057(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E115));
DFF_save_fm DFF_W1058(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E125));
DFF_save_fm DFF_W1059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E205));
DFF_save_fm DFF_W1060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E215));
DFF_save_fm DFF_W1061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E225));
DFF_save_fm DFF_W1062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E006));
DFF_save_fm DFF_W1063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E016));
DFF_save_fm DFF_W1064(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E026));
DFF_save_fm DFF_W1065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E106));
DFF_save_fm DFF_W1066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E116));
DFF_save_fm DFF_W1067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E126));
DFF_save_fm DFF_W1068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E206));
DFF_save_fm DFF_W1069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E216));
DFF_save_fm DFF_W1070(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E226));
DFF_save_fm DFF_W1071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E007));
DFF_save_fm DFF_W1072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E017));
DFF_save_fm DFF_W1073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E027));
DFF_save_fm DFF_W1074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E107));
DFF_save_fm DFF_W1075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E117));
DFF_save_fm DFF_W1076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E127));
DFF_save_fm DFF_W1077(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E207));
DFF_save_fm DFF_W1078(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E217));
DFF_save_fm DFF_W1079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E227));
DFF_save_fm DFF_W1080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F000));
DFF_save_fm DFF_W1081(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F010));
DFF_save_fm DFF_W1082(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F020));
DFF_save_fm DFF_W1083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F100));
DFF_save_fm DFF_W1084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F110));
DFF_save_fm DFF_W1085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F120));
DFF_save_fm DFF_W1086(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F200));
DFF_save_fm DFF_W1087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F210));
DFF_save_fm DFF_W1088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F220));
DFF_save_fm DFF_W1089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F001));
DFF_save_fm DFF_W1090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F011));
DFF_save_fm DFF_W1091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F021));
DFF_save_fm DFF_W1092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F101));
DFF_save_fm DFF_W1093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F111));
DFF_save_fm DFF_W1094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F121));
DFF_save_fm DFF_W1095(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F201));
DFF_save_fm DFF_W1096(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F211));
DFF_save_fm DFF_W1097(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F221));
DFF_save_fm DFF_W1098(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F002));
DFF_save_fm DFF_W1099(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F012));
DFF_save_fm DFF_W1100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F022));
DFF_save_fm DFF_W1101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F102));
DFF_save_fm DFF_W1102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F112));
DFF_save_fm DFF_W1103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F122));
DFF_save_fm DFF_W1104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F202));
DFF_save_fm DFF_W1105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F212));
DFF_save_fm DFF_W1106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F222));
DFF_save_fm DFF_W1107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F003));
DFF_save_fm DFF_W1108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F013));
DFF_save_fm DFF_W1109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F023));
DFF_save_fm DFF_W1110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F103));
DFF_save_fm DFF_W1111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F113));
DFF_save_fm DFF_W1112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F123));
DFF_save_fm DFF_W1113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F203));
DFF_save_fm DFF_W1114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F213));
DFF_save_fm DFF_W1115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F223));
DFF_save_fm DFF_W1116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F004));
DFF_save_fm DFF_W1117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F014));
DFF_save_fm DFF_W1118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F024));
DFF_save_fm DFF_W1119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F104));
DFF_save_fm DFF_W1120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F114));
DFF_save_fm DFF_W1121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F124));
DFF_save_fm DFF_W1122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F204));
DFF_save_fm DFF_W1123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F214));
DFF_save_fm DFF_W1124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F224));
DFF_save_fm DFF_W1125(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F005));
DFF_save_fm DFF_W1126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F015));
DFF_save_fm DFF_W1127(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F025));
DFF_save_fm DFF_W1128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F105));
DFF_save_fm DFF_W1129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F115));
DFF_save_fm DFF_W1130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F125));
DFF_save_fm DFF_W1131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F205));
DFF_save_fm DFF_W1132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F215));
DFF_save_fm DFF_W1133(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F225));
DFF_save_fm DFF_W1134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F006));
DFF_save_fm DFF_W1135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F016));
DFF_save_fm DFF_W1136(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F026));
DFF_save_fm DFF_W1137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F106));
DFF_save_fm DFF_W1138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F116));
DFF_save_fm DFF_W1139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F126));
DFF_save_fm DFF_W1140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F206));
DFF_save_fm DFF_W1141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F216));
DFF_save_fm DFF_W1142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F226));
DFF_save_fm DFF_W1143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F007));
DFF_save_fm DFF_W1144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F017));
DFF_save_fm DFF_W1145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F027));
DFF_save_fm DFF_W1146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F107));
DFF_save_fm DFF_W1147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F117));
DFF_save_fm DFF_W1148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F127));
DFF_save_fm DFF_W1149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F207));
DFF_save_fm DFF_W1150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F217));
DFF_save_fm DFF_W1151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F227));
ninexnine_unit ninexnine_unit_0(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20000)
);

ninexnine_unit ninexnine_unit_1(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21000)
);

ninexnine_unit ninexnine_unit_2(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22000)
);

ninexnine_unit ninexnine_unit_3(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23000)
);

ninexnine_unit ninexnine_unit_4(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24000)
);

ninexnine_unit ninexnine_unit_5(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25000)
);

ninexnine_unit ninexnine_unit_6(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26000)
);

ninexnine_unit ninexnine_unit_7(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27000)
);

assign C2000=c20000+c21000+c22000+c23000+c24000+c25000+c26000+c27000;
assign A2000=(C2000>=0)?1:0;

assign P3000=A2000;

ninexnine_unit ninexnine_unit_8(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20010)
);

ninexnine_unit ninexnine_unit_9(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21010)
);

ninexnine_unit ninexnine_unit_10(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22010)
);

ninexnine_unit ninexnine_unit_11(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23010)
);

ninexnine_unit ninexnine_unit_12(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24010)
);

ninexnine_unit ninexnine_unit_13(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25010)
);

ninexnine_unit ninexnine_unit_14(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26010)
);

ninexnine_unit ninexnine_unit_15(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27010)
);

assign C2010=c20010+c21010+c22010+c23010+c24010+c25010+c26010+c27010;
assign A2010=(C2010>=0)?1:0;

assign P3010=A2010;

ninexnine_unit ninexnine_unit_16(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20020)
);

ninexnine_unit ninexnine_unit_17(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21020)
);

ninexnine_unit ninexnine_unit_18(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22020)
);

ninexnine_unit ninexnine_unit_19(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23020)
);

ninexnine_unit ninexnine_unit_20(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24020)
);

ninexnine_unit ninexnine_unit_21(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25020)
);

ninexnine_unit ninexnine_unit_22(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26020)
);

ninexnine_unit ninexnine_unit_23(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27020)
);

assign C2020=c20020+c21020+c22020+c23020+c24020+c25020+c26020+c27020;
assign A2020=(C2020>=0)?1:0;

assign P3020=A2020;

ninexnine_unit ninexnine_unit_24(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20030)
);

ninexnine_unit ninexnine_unit_25(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21030)
);

ninexnine_unit ninexnine_unit_26(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22030)
);

ninexnine_unit ninexnine_unit_27(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23030)
);

ninexnine_unit ninexnine_unit_28(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24030)
);

ninexnine_unit ninexnine_unit_29(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25030)
);

ninexnine_unit ninexnine_unit_30(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26030)
);

ninexnine_unit ninexnine_unit_31(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27030)
);

assign C2030=c20030+c21030+c22030+c23030+c24030+c25030+c26030+c27030;
assign A2030=(C2030>=0)?1:0;

assign P3030=A2030;

ninexnine_unit ninexnine_unit_32(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20040)
);

ninexnine_unit ninexnine_unit_33(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21040)
);

ninexnine_unit ninexnine_unit_34(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22040)
);

ninexnine_unit ninexnine_unit_35(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23040)
);

ninexnine_unit ninexnine_unit_36(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24040)
);

ninexnine_unit ninexnine_unit_37(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25040)
);

ninexnine_unit ninexnine_unit_38(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26040)
);

ninexnine_unit ninexnine_unit_39(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27040)
);

assign C2040=c20040+c21040+c22040+c23040+c24040+c25040+c26040+c27040;
assign A2040=(C2040>=0)?1:0;

assign P3040=A2040;

ninexnine_unit ninexnine_unit_40(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20100)
);

ninexnine_unit ninexnine_unit_41(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21100)
);

ninexnine_unit ninexnine_unit_42(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22100)
);

ninexnine_unit ninexnine_unit_43(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23100)
);

ninexnine_unit ninexnine_unit_44(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24100)
);

ninexnine_unit ninexnine_unit_45(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25100)
);

ninexnine_unit ninexnine_unit_46(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26100)
);

ninexnine_unit ninexnine_unit_47(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27100)
);

assign C2100=c20100+c21100+c22100+c23100+c24100+c25100+c26100+c27100;
assign A2100=(C2100>=0)?1:0;

assign P3100=A2100;

ninexnine_unit ninexnine_unit_48(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20110)
);

ninexnine_unit ninexnine_unit_49(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21110)
);

ninexnine_unit ninexnine_unit_50(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22110)
);

ninexnine_unit ninexnine_unit_51(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23110)
);

ninexnine_unit ninexnine_unit_52(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24110)
);

ninexnine_unit ninexnine_unit_53(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25110)
);

ninexnine_unit ninexnine_unit_54(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26110)
);

ninexnine_unit ninexnine_unit_55(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27110)
);

assign C2110=c20110+c21110+c22110+c23110+c24110+c25110+c26110+c27110;
assign A2110=(C2110>=0)?1:0;

assign P3110=A2110;

ninexnine_unit ninexnine_unit_56(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20120)
);

ninexnine_unit ninexnine_unit_57(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21120)
);

ninexnine_unit ninexnine_unit_58(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22120)
);

ninexnine_unit ninexnine_unit_59(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23120)
);

ninexnine_unit ninexnine_unit_60(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24120)
);

ninexnine_unit ninexnine_unit_61(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25120)
);

ninexnine_unit ninexnine_unit_62(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26120)
);

ninexnine_unit ninexnine_unit_63(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27120)
);

assign C2120=c20120+c21120+c22120+c23120+c24120+c25120+c26120+c27120;
assign A2120=(C2120>=0)?1:0;

assign P3120=A2120;

ninexnine_unit ninexnine_unit_64(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20130)
);

ninexnine_unit ninexnine_unit_65(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21130)
);

ninexnine_unit ninexnine_unit_66(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22130)
);

ninexnine_unit ninexnine_unit_67(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23130)
);

ninexnine_unit ninexnine_unit_68(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24130)
);

ninexnine_unit ninexnine_unit_69(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25130)
);

ninexnine_unit ninexnine_unit_70(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26130)
);

ninexnine_unit ninexnine_unit_71(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27130)
);

assign C2130=c20130+c21130+c22130+c23130+c24130+c25130+c26130+c27130;
assign A2130=(C2130>=0)?1:0;

assign P3130=A2130;

ninexnine_unit ninexnine_unit_72(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20140)
);

ninexnine_unit ninexnine_unit_73(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21140)
);

ninexnine_unit ninexnine_unit_74(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22140)
);

ninexnine_unit ninexnine_unit_75(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23140)
);

ninexnine_unit ninexnine_unit_76(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24140)
);

ninexnine_unit ninexnine_unit_77(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25140)
);

ninexnine_unit ninexnine_unit_78(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26140)
);

ninexnine_unit ninexnine_unit_79(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27140)
);

assign C2140=c20140+c21140+c22140+c23140+c24140+c25140+c26140+c27140;
assign A2140=(C2140>=0)?1:0;

assign P3140=A2140;

ninexnine_unit ninexnine_unit_80(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20200)
);

ninexnine_unit ninexnine_unit_81(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21200)
);

ninexnine_unit ninexnine_unit_82(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22200)
);

ninexnine_unit ninexnine_unit_83(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23200)
);

ninexnine_unit ninexnine_unit_84(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24200)
);

ninexnine_unit ninexnine_unit_85(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25200)
);

ninexnine_unit ninexnine_unit_86(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26200)
);

ninexnine_unit ninexnine_unit_87(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27200)
);

assign C2200=c20200+c21200+c22200+c23200+c24200+c25200+c26200+c27200;
assign A2200=(C2200>=0)?1:0;

assign P3200=A2200;

ninexnine_unit ninexnine_unit_88(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20210)
);

ninexnine_unit ninexnine_unit_89(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21210)
);

ninexnine_unit ninexnine_unit_90(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22210)
);

ninexnine_unit ninexnine_unit_91(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23210)
);

ninexnine_unit ninexnine_unit_92(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24210)
);

ninexnine_unit ninexnine_unit_93(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25210)
);

ninexnine_unit ninexnine_unit_94(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26210)
);

ninexnine_unit ninexnine_unit_95(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27210)
);

assign C2210=c20210+c21210+c22210+c23210+c24210+c25210+c26210+c27210;
assign A2210=(C2210>=0)?1:0;

assign P3210=A2210;

ninexnine_unit ninexnine_unit_96(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20220)
);

ninexnine_unit ninexnine_unit_97(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21220)
);

ninexnine_unit ninexnine_unit_98(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22220)
);

ninexnine_unit ninexnine_unit_99(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23220)
);

ninexnine_unit ninexnine_unit_100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24220)
);

ninexnine_unit ninexnine_unit_101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25220)
);

ninexnine_unit ninexnine_unit_102(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26220)
);

ninexnine_unit ninexnine_unit_103(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27220)
);

assign C2220=c20220+c21220+c22220+c23220+c24220+c25220+c26220+c27220;
assign A2220=(C2220>=0)?1:0;

assign P3220=A2220;

ninexnine_unit ninexnine_unit_104(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20230)
);

ninexnine_unit ninexnine_unit_105(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21230)
);

ninexnine_unit ninexnine_unit_106(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22230)
);

ninexnine_unit ninexnine_unit_107(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23230)
);

ninexnine_unit ninexnine_unit_108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24230)
);

ninexnine_unit ninexnine_unit_109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25230)
);

ninexnine_unit ninexnine_unit_110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26230)
);

ninexnine_unit ninexnine_unit_111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27230)
);

assign C2230=c20230+c21230+c22230+c23230+c24230+c25230+c26230+c27230;
assign A2230=(C2230>=0)?1:0;

assign P3230=A2230;

ninexnine_unit ninexnine_unit_112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20240)
);

ninexnine_unit ninexnine_unit_113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21240)
);

ninexnine_unit ninexnine_unit_114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22240)
);

ninexnine_unit ninexnine_unit_115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23240)
);

ninexnine_unit ninexnine_unit_116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24240)
);

ninexnine_unit ninexnine_unit_117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25240)
);

ninexnine_unit ninexnine_unit_118(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26240)
);

ninexnine_unit ninexnine_unit_119(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27240)
);

assign C2240=c20240+c21240+c22240+c23240+c24240+c25240+c26240+c27240;
assign A2240=(C2240>=0)?1:0;

assign P3240=A2240;

ninexnine_unit ninexnine_unit_120(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20300)
);

ninexnine_unit ninexnine_unit_121(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21300)
);

ninexnine_unit ninexnine_unit_122(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22300)
);

ninexnine_unit ninexnine_unit_123(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23300)
);

ninexnine_unit ninexnine_unit_124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24300)
);

ninexnine_unit ninexnine_unit_125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25300)
);

ninexnine_unit ninexnine_unit_126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26300)
);

ninexnine_unit ninexnine_unit_127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27300)
);

assign C2300=c20300+c21300+c22300+c23300+c24300+c25300+c26300+c27300;
assign A2300=(C2300>=0)?1:0;

assign P3300=A2300;

ninexnine_unit ninexnine_unit_128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20310)
);

ninexnine_unit ninexnine_unit_129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21310)
);

ninexnine_unit ninexnine_unit_130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22310)
);

ninexnine_unit ninexnine_unit_131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23310)
);

ninexnine_unit ninexnine_unit_132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24310)
);

ninexnine_unit ninexnine_unit_133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25310)
);

ninexnine_unit ninexnine_unit_134(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26310)
);

ninexnine_unit ninexnine_unit_135(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27310)
);

assign C2310=c20310+c21310+c22310+c23310+c24310+c25310+c26310+c27310;
assign A2310=(C2310>=0)?1:0;

assign P3310=A2310;

ninexnine_unit ninexnine_unit_136(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20320)
);

ninexnine_unit ninexnine_unit_137(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21320)
);

ninexnine_unit ninexnine_unit_138(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22320)
);

ninexnine_unit ninexnine_unit_139(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23320)
);

ninexnine_unit ninexnine_unit_140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24320)
);

ninexnine_unit ninexnine_unit_141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25320)
);

ninexnine_unit ninexnine_unit_142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26320)
);

ninexnine_unit ninexnine_unit_143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27320)
);

assign C2320=c20320+c21320+c22320+c23320+c24320+c25320+c26320+c27320;
assign A2320=(C2320>=0)?1:0;

assign P3320=A2320;

ninexnine_unit ninexnine_unit_144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20330)
);

ninexnine_unit ninexnine_unit_145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21330)
);

ninexnine_unit ninexnine_unit_146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22330)
);

ninexnine_unit ninexnine_unit_147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23330)
);

ninexnine_unit ninexnine_unit_148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24330)
);

ninexnine_unit ninexnine_unit_149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25330)
);

ninexnine_unit ninexnine_unit_150(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26330)
);

ninexnine_unit ninexnine_unit_151(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27330)
);

assign C2330=c20330+c21330+c22330+c23330+c24330+c25330+c26330+c27330;
assign A2330=(C2330>=0)?1:0;

assign P3330=A2330;

ninexnine_unit ninexnine_unit_152(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20340)
);

ninexnine_unit ninexnine_unit_153(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21340)
);

ninexnine_unit ninexnine_unit_154(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22340)
);

ninexnine_unit ninexnine_unit_155(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23340)
);

ninexnine_unit ninexnine_unit_156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24340)
);

ninexnine_unit ninexnine_unit_157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25340)
);

ninexnine_unit ninexnine_unit_158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26340)
);

ninexnine_unit ninexnine_unit_159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27340)
);

assign C2340=c20340+c21340+c22340+c23340+c24340+c25340+c26340+c27340;
assign A2340=(C2340>=0)?1:0;

assign P3340=A2340;

ninexnine_unit ninexnine_unit_160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20400)
);

ninexnine_unit ninexnine_unit_161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21400)
);

ninexnine_unit ninexnine_unit_162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22400)
);

ninexnine_unit ninexnine_unit_163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23400)
);

ninexnine_unit ninexnine_unit_164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24400)
);

ninexnine_unit ninexnine_unit_165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25400)
);

ninexnine_unit ninexnine_unit_166(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26400)
);

ninexnine_unit ninexnine_unit_167(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27400)
);

assign C2400=c20400+c21400+c22400+c23400+c24400+c25400+c26400+c27400;
assign A2400=(C2400>=0)?1:0;

assign P3400=A2400;

ninexnine_unit ninexnine_unit_168(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20410)
);

ninexnine_unit ninexnine_unit_169(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21410)
);

ninexnine_unit ninexnine_unit_170(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22410)
);

ninexnine_unit ninexnine_unit_171(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23410)
);

ninexnine_unit ninexnine_unit_172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24410)
);

ninexnine_unit ninexnine_unit_173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25410)
);

ninexnine_unit ninexnine_unit_174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26410)
);

ninexnine_unit ninexnine_unit_175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27410)
);

assign C2410=c20410+c21410+c22410+c23410+c24410+c25410+c26410+c27410;
assign A2410=(C2410>=0)?1:0;

assign P3410=A2410;

ninexnine_unit ninexnine_unit_176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20420)
);

ninexnine_unit ninexnine_unit_177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21420)
);

ninexnine_unit ninexnine_unit_178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22420)
);

ninexnine_unit ninexnine_unit_179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23420)
);

ninexnine_unit ninexnine_unit_180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24420)
);

ninexnine_unit ninexnine_unit_181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25420)
);

ninexnine_unit ninexnine_unit_182(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26420)
);

ninexnine_unit ninexnine_unit_183(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27420)
);

assign C2420=c20420+c21420+c22420+c23420+c24420+c25420+c26420+c27420;
assign A2420=(C2420>=0)?1:0;

assign P3420=A2420;

ninexnine_unit ninexnine_unit_184(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20430)
);

ninexnine_unit ninexnine_unit_185(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21430)
);

ninexnine_unit ninexnine_unit_186(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22430)
);

ninexnine_unit ninexnine_unit_187(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23430)
);

ninexnine_unit ninexnine_unit_188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24430)
);

ninexnine_unit ninexnine_unit_189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25430)
);

ninexnine_unit ninexnine_unit_190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26430)
);

ninexnine_unit ninexnine_unit_191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27430)
);

assign C2430=c20430+c21430+c22430+c23430+c24430+c25430+c26430+c27430;
assign A2430=(C2430>=0)?1:0;

assign P3430=A2430;

ninexnine_unit ninexnine_unit_192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20440)
);

ninexnine_unit ninexnine_unit_193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21440)
);

ninexnine_unit ninexnine_unit_194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22440)
);

ninexnine_unit ninexnine_unit_195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23440)
);

ninexnine_unit ninexnine_unit_196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24440)
);

ninexnine_unit ninexnine_unit_197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25440)
);

ninexnine_unit ninexnine_unit_198(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26440)
);

ninexnine_unit ninexnine_unit_199(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27440)
);

assign C2440=c20440+c21440+c22440+c23440+c24440+c25440+c26440+c27440;
assign A2440=(C2440>=0)?1:0;

assign P3440=A2440;

ninexnine_unit ninexnine_unit_200(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20001)
);

ninexnine_unit ninexnine_unit_201(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21001)
);

ninexnine_unit ninexnine_unit_202(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22001)
);

ninexnine_unit ninexnine_unit_203(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23001)
);

ninexnine_unit ninexnine_unit_204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24001)
);

ninexnine_unit ninexnine_unit_205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25001)
);

ninexnine_unit ninexnine_unit_206(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26001)
);

ninexnine_unit ninexnine_unit_207(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27001)
);

assign C2001=c20001+c21001+c22001+c23001+c24001+c25001+c26001+c27001;
assign A2001=(C2001>=0)?1:0;

assign P3001=A2001;

ninexnine_unit ninexnine_unit_208(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20011)
);

ninexnine_unit ninexnine_unit_209(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21011)
);

ninexnine_unit ninexnine_unit_210(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22011)
);

ninexnine_unit ninexnine_unit_211(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23011)
);

ninexnine_unit ninexnine_unit_212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24011)
);

ninexnine_unit ninexnine_unit_213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25011)
);

ninexnine_unit ninexnine_unit_214(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26011)
);

ninexnine_unit ninexnine_unit_215(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27011)
);

assign C2011=c20011+c21011+c22011+c23011+c24011+c25011+c26011+c27011;
assign A2011=(C2011>=0)?1:0;

assign P3011=A2011;

ninexnine_unit ninexnine_unit_216(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20021)
);

ninexnine_unit ninexnine_unit_217(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21021)
);

ninexnine_unit ninexnine_unit_218(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22021)
);

ninexnine_unit ninexnine_unit_219(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23021)
);

ninexnine_unit ninexnine_unit_220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24021)
);

ninexnine_unit ninexnine_unit_221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25021)
);

ninexnine_unit ninexnine_unit_222(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26021)
);

ninexnine_unit ninexnine_unit_223(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27021)
);

assign C2021=c20021+c21021+c22021+c23021+c24021+c25021+c26021+c27021;
assign A2021=(C2021>=0)?1:0;

assign P3021=A2021;

ninexnine_unit ninexnine_unit_224(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20031)
);

ninexnine_unit ninexnine_unit_225(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21031)
);

ninexnine_unit ninexnine_unit_226(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22031)
);

ninexnine_unit ninexnine_unit_227(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23031)
);

ninexnine_unit ninexnine_unit_228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24031)
);

ninexnine_unit ninexnine_unit_229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25031)
);

ninexnine_unit ninexnine_unit_230(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26031)
);

ninexnine_unit ninexnine_unit_231(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27031)
);

assign C2031=c20031+c21031+c22031+c23031+c24031+c25031+c26031+c27031;
assign A2031=(C2031>=0)?1:0;

assign P3031=A2031;

ninexnine_unit ninexnine_unit_232(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20041)
);

ninexnine_unit ninexnine_unit_233(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21041)
);

ninexnine_unit ninexnine_unit_234(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22041)
);

ninexnine_unit ninexnine_unit_235(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23041)
);

ninexnine_unit ninexnine_unit_236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24041)
);

ninexnine_unit ninexnine_unit_237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25041)
);

ninexnine_unit ninexnine_unit_238(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26041)
);

ninexnine_unit ninexnine_unit_239(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27041)
);

assign C2041=c20041+c21041+c22041+c23041+c24041+c25041+c26041+c27041;
assign A2041=(C2041>=0)?1:0;

assign P3041=A2041;

ninexnine_unit ninexnine_unit_240(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20101)
);

ninexnine_unit ninexnine_unit_241(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21101)
);

ninexnine_unit ninexnine_unit_242(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22101)
);

ninexnine_unit ninexnine_unit_243(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23101)
);

ninexnine_unit ninexnine_unit_244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24101)
);

ninexnine_unit ninexnine_unit_245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25101)
);

ninexnine_unit ninexnine_unit_246(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26101)
);

ninexnine_unit ninexnine_unit_247(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27101)
);

assign C2101=c20101+c21101+c22101+c23101+c24101+c25101+c26101+c27101;
assign A2101=(C2101>=0)?1:0;

assign P3101=A2101;

ninexnine_unit ninexnine_unit_248(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20111)
);

ninexnine_unit ninexnine_unit_249(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21111)
);

ninexnine_unit ninexnine_unit_250(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22111)
);

ninexnine_unit ninexnine_unit_251(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23111)
);

ninexnine_unit ninexnine_unit_252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24111)
);

ninexnine_unit ninexnine_unit_253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25111)
);

ninexnine_unit ninexnine_unit_254(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26111)
);

ninexnine_unit ninexnine_unit_255(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27111)
);

assign C2111=c20111+c21111+c22111+c23111+c24111+c25111+c26111+c27111;
assign A2111=(C2111>=0)?1:0;

assign P3111=A2111;

ninexnine_unit ninexnine_unit_256(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20121)
);

ninexnine_unit ninexnine_unit_257(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21121)
);

ninexnine_unit ninexnine_unit_258(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22121)
);

ninexnine_unit ninexnine_unit_259(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23121)
);

ninexnine_unit ninexnine_unit_260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24121)
);

ninexnine_unit ninexnine_unit_261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25121)
);

ninexnine_unit ninexnine_unit_262(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26121)
);

ninexnine_unit ninexnine_unit_263(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27121)
);

assign C2121=c20121+c21121+c22121+c23121+c24121+c25121+c26121+c27121;
assign A2121=(C2121>=0)?1:0;

assign P3121=A2121;

ninexnine_unit ninexnine_unit_264(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20131)
);

ninexnine_unit ninexnine_unit_265(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21131)
);

ninexnine_unit ninexnine_unit_266(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22131)
);

ninexnine_unit ninexnine_unit_267(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23131)
);

ninexnine_unit ninexnine_unit_268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24131)
);

ninexnine_unit ninexnine_unit_269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25131)
);

ninexnine_unit ninexnine_unit_270(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26131)
);

ninexnine_unit ninexnine_unit_271(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27131)
);

assign C2131=c20131+c21131+c22131+c23131+c24131+c25131+c26131+c27131;
assign A2131=(C2131>=0)?1:0;

assign P3131=A2131;

ninexnine_unit ninexnine_unit_272(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20141)
);

ninexnine_unit ninexnine_unit_273(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21141)
);

ninexnine_unit ninexnine_unit_274(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22141)
);

ninexnine_unit ninexnine_unit_275(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23141)
);

ninexnine_unit ninexnine_unit_276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24141)
);

ninexnine_unit ninexnine_unit_277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25141)
);

ninexnine_unit ninexnine_unit_278(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26141)
);

ninexnine_unit ninexnine_unit_279(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27141)
);

assign C2141=c20141+c21141+c22141+c23141+c24141+c25141+c26141+c27141;
assign A2141=(C2141>=0)?1:0;

assign P3141=A2141;

ninexnine_unit ninexnine_unit_280(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20201)
);

ninexnine_unit ninexnine_unit_281(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21201)
);

ninexnine_unit ninexnine_unit_282(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22201)
);

ninexnine_unit ninexnine_unit_283(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23201)
);

ninexnine_unit ninexnine_unit_284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24201)
);

ninexnine_unit ninexnine_unit_285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25201)
);

ninexnine_unit ninexnine_unit_286(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26201)
);

ninexnine_unit ninexnine_unit_287(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27201)
);

assign C2201=c20201+c21201+c22201+c23201+c24201+c25201+c26201+c27201;
assign A2201=(C2201>=0)?1:0;

assign P3201=A2201;

ninexnine_unit ninexnine_unit_288(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20211)
);

ninexnine_unit ninexnine_unit_289(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21211)
);

ninexnine_unit ninexnine_unit_290(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22211)
);

ninexnine_unit ninexnine_unit_291(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23211)
);

ninexnine_unit ninexnine_unit_292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24211)
);

ninexnine_unit ninexnine_unit_293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25211)
);

ninexnine_unit ninexnine_unit_294(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26211)
);

ninexnine_unit ninexnine_unit_295(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27211)
);

assign C2211=c20211+c21211+c22211+c23211+c24211+c25211+c26211+c27211;
assign A2211=(C2211>=0)?1:0;

assign P3211=A2211;

ninexnine_unit ninexnine_unit_296(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20221)
);

ninexnine_unit ninexnine_unit_297(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21221)
);

ninexnine_unit ninexnine_unit_298(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22221)
);

ninexnine_unit ninexnine_unit_299(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23221)
);

ninexnine_unit ninexnine_unit_300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24221)
);

ninexnine_unit ninexnine_unit_301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25221)
);

ninexnine_unit ninexnine_unit_302(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26221)
);

ninexnine_unit ninexnine_unit_303(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27221)
);

assign C2221=c20221+c21221+c22221+c23221+c24221+c25221+c26221+c27221;
assign A2221=(C2221>=0)?1:0;

assign P3221=A2221;

ninexnine_unit ninexnine_unit_304(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20231)
);

ninexnine_unit ninexnine_unit_305(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21231)
);

ninexnine_unit ninexnine_unit_306(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22231)
);

ninexnine_unit ninexnine_unit_307(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23231)
);

ninexnine_unit ninexnine_unit_308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24231)
);

ninexnine_unit ninexnine_unit_309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25231)
);

ninexnine_unit ninexnine_unit_310(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26231)
);

ninexnine_unit ninexnine_unit_311(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27231)
);

assign C2231=c20231+c21231+c22231+c23231+c24231+c25231+c26231+c27231;
assign A2231=(C2231>=0)?1:0;

assign P3231=A2231;

ninexnine_unit ninexnine_unit_312(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20241)
);

ninexnine_unit ninexnine_unit_313(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21241)
);

ninexnine_unit ninexnine_unit_314(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22241)
);

ninexnine_unit ninexnine_unit_315(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23241)
);

ninexnine_unit ninexnine_unit_316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24241)
);

ninexnine_unit ninexnine_unit_317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25241)
);

ninexnine_unit ninexnine_unit_318(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26241)
);

ninexnine_unit ninexnine_unit_319(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27241)
);

assign C2241=c20241+c21241+c22241+c23241+c24241+c25241+c26241+c27241;
assign A2241=(C2241>=0)?1:0;

assign P3241=A2241;

ninexnine_unit ninexnine_unit_320(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20301)
);

ninexnine_unit ninexnine_unit_321(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21301)
);

ninexnine_unit ninexnine_unit_322(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22301)
);

ninexnine_unit ninexnine_unit_323(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23301)
);

ninexnine_unit ninexnine_unit_324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24301)
);

ninexnine_unit ninexnine_unit_325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25301)
);

ninexnine_unit ninexnine_unit_326(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26301)
);

ninexnine_unit ninexnine_unit_327(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27301)
);

assign C2301=c20301+c21301+c22301+c23301+c24301+c25301+c26301+c27301;
assign A2301=(C2301>=0)?1:0;

assign P3301=A2301;

ninexnine_unit ninexnine_unit_328(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20311)
);

ninexnine_unit ninexnine_unit_329(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21311)
);

ninexnine_unit ninexnine_unit_330(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22311)
);

ninexnine_unit ninexnine_unit_331(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23311)
);

ninexnine_unit ninexnine_unit_332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24311)
);

ninexnine_unit ninexnine_unit_333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25311)
);

ninexnine_unit ninexnine_unit_334(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26311)
);

ninexnine_unit ninexnine_unit_335(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27311)
);

assign C2311=c20311+c21311+c22311+c23311+c24311+c25311+c26311+c27311;
assign A2311=(C2311>=0)?1:0;

assign P3311=A2311;

ninexnine_unit ninexnine_unit_336(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20321)
);

ninexnine_unit ninexnine_unit_337(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21321)
);

ninexnine_unit ninexnine_unit_338(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22321)
);

ninexnine_unit ninexnine_unit_339(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23321)
);

ninexnine_unit ninexnine_unit_340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24321)
);

ninexnine_unit ninexnine_unit_341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25321)
);

ninexnine_unit ninexnine_unit_342(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26321)
);

ninexnine_unit ninexnine_unit_343(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27321)
);

assign C2321=c20321+c21321+c22321+c23321+c24321+c25321+c26321+c27321;
assign A2321=(C2321>=0)?1:0;

assign P3321=A2321;

ninexnine_unit ninexnine_unit_344(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20331)
);

ninexnine_unit ninexnine_unit_345(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21331)
);

ninexnine_unit ninexnine_unit_346(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22331)
);

ninexnine_unit ninexnine_unit_347(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23331)
);

ninexnine_unit ninexnine_unit_348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24331)
);

ninexnine_unit ninexnine_unit_349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25331)
);

ninexnine_unit ninexnine_unit_350(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26331)
);

ninexnine_unit ninexnine_unit_351(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27331)
);

assign C2331=c20331+c21331+c22331+c23331+c24331+c25331+c26331+c27331;
assign A2331=(C2331>=0)?1:0;

assign P3331=A2331;

ninexnine_unit ninexnine_unit_352(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20341)
);

ninexnine_unit ninexnine_unit_353(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21341)
);

ninexnine_unit ninexnine_unit_354(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22341)
);

ninexnine_unit ninexnine_unit_355(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23341)
);

ninexnine_unit ninexnine_unit_356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24341)
);

ninexnine_unit ninexnine_unit_357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25341)
);

ninexnine_unit ninexnine_unit_358(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26341)
);

ninexnine_unit ninexnine_unit_359(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27341)
);

assign C2341=c20341+c21341+c22341+c23341+c24341+c25341+c26341+c27341;
assign A2341=(C2341>=0)?1:0;

assign P3341=A2341;

ninexnine_unit ninexnine_unit_360(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20401)
);

ninexnine_unit ninexnine_unit_361(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21401)
);

ninexnine_unit ninexnine_unit_362(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22401)
);

ninexnine_unit ninexnine_unit_363(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23401)
);

ninexnine_unit ninexnine_unit_364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24401)
);

ninexnine_unit ninexnine_unit_365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25401)
);

ninexnine_unit ninexnine_unit_366(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26401)
);

ninexnine_unit ninexnine_unit_367(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27401)
);

assign C2401=c20401+c21401+c22401+c23401+c24401+c25401+c26401+c27401;
assign A2401=(C2401>=0)?1:0;

assign P3401=A2401;

ninexnine_unit ninexnine_unit_368(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20411)
);

ninexnine_unit ninexnine_unit_369(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21411)
);

ninexnine_unit ninexnine_unit_370(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22411)
);

ninexnine_unit ninexnine_unit_371(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23411)
);

ninexnine_unit ninexnine_unit_372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24411)
);

ninexnine_unit ninexnine_unit_373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25411)
);

ninexnine_unit ninexnine_unit_374(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26411)
);

ninexnine_unit ninexnine_unit_375(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27411)
);

assign C2411=c20411+c21411+c22411+c23411+c24411+c25411+c26411+c27411;
assign A2411=(C2411>=0)?1:0;

assign P3411=A2411;

ninexnine_unit ninexnine_unit_376(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20421)
);

ninexnine_unit ninexnine_unit_377(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21421)
);

ninexnine_unit ninexnine_unit_378(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22421)
);

ninexnine_unit ninexnine_unit_379(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23421)
);

ninexnine_unit ninexnine_unit_380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24421)
);

ninexnine_unit ninexnine_unit_381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25421)
);

ninexnine_unit ninexnine_unit_382(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26421)
);

ninexnine_unit ninexnine_unit_383(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27421)
);

assign C2421=c20421+c21421+c22421+c23421+c24421+c25421+c26421+c27421;
assign A2421=(C2421>=0)?1:0;

assign P3421=A2421;

ninexnine_unit ninexnine_unit_384(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20431)
);

ninexnine_unit ninexnine_unit_385(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21431)
);

ninexnine_unit ninexnine_unit_386(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22431)
);

ninexnine_unit ninexnine_unit_387(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23431)
);

ninexnine_unit ninexnine_unit_388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24431)
);

ninexnine_unit ninexnine_unit_389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25431)
);

ninexnine_unit ninexnine_unit_390(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26431)
);

ninexnine_unit ninexnine_unit_391(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27431)
);

assign C2431=c20431+c21431+c22431+c23431+c24431+c25431+c26431+c27431;
assign A2431=(C2431>=0)?1:0;

assign P3431=A2431;

ninexnine_unit ninexnine_unit_392(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20441)
);

ninexnine_unit ninexnine_unit_393(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21441)
);

ninexnine_unit ninexnine_unit_394(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22441)
);

ninexnine_unit ninexnine_unit_395(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23441)
);

ninexnine_unit ninexnine_unit_396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24441)
);

ninexnine_unit ninexnine_unit_397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25441)
);

ninexnine_unit ninexnine_unit_398(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26441)
);

ninexnine_unit ninexnine_unit_399(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27441)
);

assign C2441=c20441+c21441+c22441+c23441+c24441+c25441+c26441+c27441;
assign A2441=(C2441>=0)?1:0;

assign P3441=A2441;

ninexnine_unit ninexnine_unit_400(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20002)
);

ninexnine_unit ninexnine_unit_401(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21002)
);

ninexnine_unit ninexnine_unit_402(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22002)
);

ninexnine_unit ninexnine_unit_403(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23002)
);

ninexnine_unit ninexnine_unit_404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24002)
);

ninexnine_unit ninexnine_unit_405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25002)
);

ninexnine_unit ninexnine_unit_406(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26002)
);

ninexnine_unit ninexnine_unit_407(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27002)
);

assign C2002=c20002+c21002+c22002+c23002+c24002+c25002+c26002+c27002;
assign A2002=(C2002>=0)?1:0;

assign P3002=A2002;

ninexnine_unit ninexnine_unit_408(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20012)
);

ninexnine_unit ninexnine_unit_409(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21012)
);

ninexnine_unit ninexnine_unit_410(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22012)
);

ninexnine_unit ninexnine_unit_411(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23012)
);

ninexnine_unit ninexnine_unit_412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24012)
);

ninexnine_unit ninexnine_unit_413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25012)
);

ninexnine_unit ninexnine_unit_414(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26012)
);

ninexnine_unit ninexnine_unit_415(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27012)
);

assign C2012=c20012+c21012+c22012+c23012+c24012+c25012+c26012+c27012;
assign A2012=(C2012>=0)?1:0;

assign P3012=A2012;

ninexnine_unit ninexnine_unit_416(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20022)
);

ninexnine_unit ninexnine_unit_417(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21022)
);

ninexnine_unit ninexnine_unit_418(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22022)
);

ninexnine_unit ninexnine_unit_419(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23022)
);

ninexnine_unit ninexnine_unit_420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24022)
);

ninexnine_unit ninexnine_unit_421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25022)
);

ninexnine_unit ninexnine_unit_422(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26022)
);

ninexnine_unit ninexnine_unit_423(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27022)
);

assign C2022=c20022+c21022+c22022+c23022+c24022+c25022+c26022+c27022;
assign A2022=(C2022>=0)?1:0;

assign P3022=A2022;

ninexnine_unit ninexnine_unit_424(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20032)
);

ninexnine_unit ninexnine_unit_425(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21032)
);

ninexnine_unit ninexnine_unit_426(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22032)
);

ninexnine_unit ninexnine_unit_427(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23032)
);

ninexnine_unit ninexnine_unit_428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24032)
);

ninexnine_unit ninexnine_unit_429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25032)
);

ninexnine_unit ninexnine_unit_430(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26032)
);

ninexnine_unit ninexnine_unit_431(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27032)
);

assign C2032=c20032+c21032+c22032+c23032+c24032+c25032+c26032+c27032;
assign A2032=(C2032>=0)?1:0;

assign P3032=A2032;

ninexnine_unit ninexnine_unit_432(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20042)
);

ninexnine_unit ninexnine_unit_433(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21042)
);

ninexnine_unit ninexnine_unit_434(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22042)
);

ninexnine_unit ninexnine_unit_435(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23042)
);

ninexnine_unit ninexnine_unit_436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24042)
);

ninexnine_unit ninexnine_unit_437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25042)
);

ninexnine_unit ninexnine_unit_438(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26042)
);

ninexnine_unit ninexnine_unit_439(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27042)
);

assign C2042=c20042+c21042+c22042+c23042+c24042+c25042+c26042+c27042;
assign A2042=(C2042>=0)?1:0;

assign P3042=A2042;

ninexnine_unit ninexnine_unit_440(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20102)
);

ninexnine_unit ninexnine_unit_441(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21102)
);

ninexnine_unit ninexnine_unit_442(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22102)
);

ninexnine_unit ninexnine_unit_443(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23102)
);

ninexnine_unit ninexnine_unit_444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24102)
);

ninexnine_unit ninexnine_unit_445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25102)
);

ninexnine_unit ninexnine_unit_446(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26102)
);

ninexnine_unit ninexnine_unit_447(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27102)
);

assign C2102=c20102+c21102+c22102+c23102+c24102+c25102+c26102+c27102;
assign A2102=(C2102>=0)?1:0;

assign P3102=A2102;

ninexnine_unit ninexnine_unit_448(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20112)
);

ninexnine_unit ninexnine_unit_449(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21112)
);

ninexnine_unit ninexnine_unit_450(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22112)
);

ninexnine_unit ninexnine_unit_451(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23112)
);

ninexnine_unit ninexnine_unit_452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24112)
);

ninexnine_unit ninexnine_unit_453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25112)
);

ninexnine_unit ninexnine_unit_454(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26112)
);

ninexnine_unit ninexnine_unit_455(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27112)
);

assign C2112=c20112+c21112+c22112+c23112+c24112+c25112+c26112+c27112;
assign A2112=(C2112>=0)?1:0;

assign P3112=A2112;

ninexnine_unit ninexnine_unit_456(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20122)
);

ninexnine_unit ninexnine_unit_457(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21122)
);

ninexnine_unit ninexnine_unit_458(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22122)
);

ninexnine_unit ninexnine_unit_459(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23122)
);

ninexnine_unit ninexnine_unit_460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24122)
);

ninexnine_unit ninexnine_unit_461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25122)
);

ninexnine_unit ninexnine_unit_462(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26122)
);

ninexnine_unit ninexnine_unit_463(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27122)
);

assign C2122=c20122+c21122+c22122+c23122+c24122+c25122+c26122+c27122;
assign A2122=(C2122>=0)?1:0;

assign P3122=A2122;

ninexnine_unit ninexnine_unit_464(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20132)
);

ninexnine_unit ninexnine_unit_465(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21132)
);

ninexnine_unit ninexnine_unit_466(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22132)
);

ninexnine_unit ninexnine_unit_467(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23132)
);

ninexnine_unit ninexnine_unit_468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24132)
);

ninexnine_unit ninexnine_unit_469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25132)
);

ninexnine_unit ninexnine_unit_470(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26132)
);

ninexnine_unit ninexnine_unit_471(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27132)
);

assign C2132=c20132+c21132+c22132+c23132+c24132+c25132+c26132+c27132;
assign A2132=(C2132>=0)?1:0;

assign P3132=A2132;

ninexnine_unit ninexnine_unit_472(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20142)
);

ninexnine_unit ninexnine_unit_473(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21142)
);

ninexnine_unit ninexnine_unit_474(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22142)
);

ninexnine_unit ninexnine_unit_475(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23142)
);

ninexnine_unit ninexnine_unit_476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24142)
);

ninexnine_unit ninexnine_unit_477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25142)
);

ninexnine_unit ninexnine_unit_478(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26142)
);

ninexnine_unit ninexnine_unit_479(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27142)
);

assign C2142=c20142+c21142+c22142+c23142+c24142+c25142+c26142+c27142;
assign A2142=(C2142>=0)?1:0;

assign P3142=A2142;

ninexnine_unit ninexnine_unit_480(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20202)
);

ninexnine_unit ninexnine_unit_481(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21202)
);

ninexnine_unit ninexnine_unit_482(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22202)
);

ninexnine_unit ninexnine_unit_483(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23202)
);

ninexnine_unit ninexnine_unit_484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24202)
);

ninexnine_unit ninexnine_unit_485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25202)
);

ninexnine_unit ninexnine_unit_486(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26202)
);

ninexnine_unit ninexnine_unit_487(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27202)
);

assign C2202=c20202+c21202+c22202+c23202+c24202+c25202+c26202+c27202;
assign A2202=(C2202>=0)?1:0;

assign P3202=A2202;

ninexnine_unit ninexnine_unit_488(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20212)
);

ninexnine_unit ninexnine_unit_489(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21212)
);

ninexnine_unit ninexnine_unit_490(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22212)
);

ninexnine_unit ninexnine_unit_491(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23212)
);

ninexnine_unit ninexnine_unit_492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24212)
);

ninexnine_unit ninexnine_unit_493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25212)
);

ninexnine_unit ninexnine_unit_494(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26212)
);

ninexnine_unit ninexnine_unit_495(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27212)
);

assign C2212=c20212+c21212+c22212+c23212+c24212+c25212+c26212+c27212;
assign A2212=(C2212>=0)?1:0;

assign P3212=A2212;

ninexnine_unit ninexnine_unit_496(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20222)
);

ninexnine_unit ninexnine_unit_497(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21222)
);

ninexnine_unit ninexnine_unit_498(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22222)
);

ninexnine_unit ninexnine_unit_499(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23222)
);

ninexnine_unit ninexnine_unit_500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24222)
);

ninexnine_unit ninexnine_unit_501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25222)
);

ninexnine_unit ninexnine_unit_502(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26222)
);

ninexnine_unit ninexnine_unit_503(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27222)
);

assign C2222=c20222+c21222+c22222+c23222+c24222+c25222+c26222+c27222;
assign A2222=(C2222>=0)?1:0;

assign P3222=A2222;

ninexnine_unit ninexnine_unit_504(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20232)
);

ninexnine_unit ninexnine_unit_505(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21232)
);

ninexnine_unit ninexnine_unit_506(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22232)
);

ninexnine_unit ninexnine_unit_507(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23232)
);

ninexnine_unit ninexnine_unit_508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24232)
);

ninexnine_unit ninexnine_unit_509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25232)
);

ninexnine_unit ninexnine_unit_510(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26232)
);

ninexnine_unit ninexnine_unit_511(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27232)
);

assign C2232=c20232+c21232+c22232+c23232+c24232+c25232+c26232+c27232;
assign A2232=(C2232>=0)?1:0;

assign P3232=A2232;

ninexnine_unit ninexnine_unit_512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20242)
);

ninexnine_unit ninexnine_unit_513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21242)
);

ninexnine_unit ninexnine_unit_514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22242)
);

ninexnine_unit ninexnine_unit_515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23242)
);

ninexnine_unit ninexnine_unit_516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24242)
);

ninexnine_unit ninexnine_unit_517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25242)
);

ninexnine_unit ninexnine_unit_518(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26242)
);

ninexnine_unit ninexnine_unit_519(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27242)
);

assign C2242=c20242+c21242+c22242+c23242+c24242+c25242+c26242+c27242;
assign A2242=(C2242>=0)?1:0;

assign P3242=A2242;

ninexnine_unit ninexnine_unit_520(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20302)
);

ninexnine_unit ninexnine_unit_521(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21302)
);

ninexnine_unit ninexnine_unit_522(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22302)
);

ninexnine_unit ninexnine_unit_523(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23302)
);

ninexnine_unit ninexnine_unit_524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24302)
);

ninexnine_unit ninexnine_unit_525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25302)
);

ninexnine_unit ninexnine_unit_526(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26302)
);

ninexnine_unit ninexnine_unit_527(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27302)
);

assign C2302=c20302+c21302+c22302+c23302+c24302+c25302+c26302+c27302;
assign A2302=(C2302>=0)?1:0;

assign P3302=A2302;

ninexnine_unit ninexnine_unit_528(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20312)
);

ninexnine_unit ninexnine_unit_529(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21312)
);

ninexnine_unit ninexnine_unit_530(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22312)
);

ninexnine_unit ninexnine_unit_531(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23312)
);

ninexnine_unit ninexnine_unit_532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24312)
);

ninexnine_unit ninexnine_unit_533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25312)
);

ninexnine_unit ninexnine_unit_534(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26312)
);

ninexnine_unit ninexnine_unit_535(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27312)
);

assign C2312=c20312+c21312+c22312+c23312+c24312+c25312+c26312+c27312;
assign A2312=(C2312>=0)?1:0;

assign P3312=A2312;

ninexnine_unit ninexnine_unit_536(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20322)
);

ninexnine_unit ninexnine_unit_537(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21322)
);

ninexnine_unit ninexnine_unit_538(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22322)
);

ninexnine_unit ninexnine_unit_539(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23322)
);

ninexnine_unit ninexnine_unit_540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24322)
);

ninexnine_unit ninexnine_unit_541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25322)
);

ninexnine_unit ninexnine_unit_542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26322)
);

ninexnine_unit ninexnine_unit_543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27322)
);

assign C2322=c20322+c21322+c22322+c23322+c24322+c25322+c26322+c27322;
assign A2322=(C2322>=0)?1:0;

assign P3322=A2322;

ninexnine_unit ninexnine_unit_544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20332)
);

ninexnine_unit ninexnine_unit_545(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21332)
);

ninexnine_unit ninexnine_unit_546(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22332)
);

ninexnine_unit ninexnine_unit_547(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23332)
);

ninexnine_unit ninexnine_unit_548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24332)
);

ninexnine_unit ninexnine_unit_549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25332)
);

ninexnine_unit ninexnine_unit_550(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26332)
);

ninexnine_unit ninexnine_unit_551(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27332)
);

assign C2332=c20332+c21332+c22332+c23332+c24332+c25332+c26332+c27332;
assign A2332=(C2332>=0)?1:0;

assign P3332=A2332;

ninexnine_unit ninexnine_unit_552(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20342)
);

ninexnine_unit ninexnine_unit_553(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21342)
);

ninexnine_unit ninexnine_unit_554(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22342)
);

ninexnine_unit ninexnine_unit_555(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23342)
);

ninexnine_unit ninexnine_unit_556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24342)
);

ninexnine_unit ninexnine_unit_557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25342)
);

ninexnine_unit ninexnine_unit_558(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26342)
);

ninexnine_unit ninexnine_unit_559(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27342)
);

assign C2342=c20342+c21342+c22342+c23342+c24342+c25342+c26342+c27342;
assign A2342=(C2342>=0)?1:0;

assign P3342=A2342;

ninexnine_unit ninexnine_unit_560(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20402)
);

ninexnine_unit ninexnine_unit_561(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21402)
);

ninexnine_unit ninexnine_unit_562(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22402)
);

ninexnine_unit ninexnine_unit_563(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23402)
);

ninexnine_unit ninexnine_unit_564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24402)
);

ninexnine_unit ninexnine_unit_565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25402)
);

ninexnine_unit ninexnine_unit_566(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26402)
);

ninexnine_unit ninexnine_unit_567(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27402)
);

assign C2402=c20402+c21402+c22402+c23402+c24402+c25402+c26402+c27402;
assign A2402=(C2402>=0)?1:0;

assign P3402=A2402;

ninexnine_unit ninexnine_unit_568(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20412)
);

ninexnine_unit ninexnine_unit_569(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21412)
);

ninexnine_unit ninexnine_unit_570(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22412)
);

ninexnine_unit ninexnine_unit_571(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23412)
);

ninexnine_unit ninexnine_unit_572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24412)
);

ninexnine_unit ninexnine_unit_573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25412)
);

ninexnine_unit ninexnine_unit_574(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26412)
);

ninexnine_unit ninexnine_unit_575(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27412)
);

assign C2412=c20412+c21412+c22412+c23412+c24412+c25412+c26412+c27412;
assign A2412=(C2412>=0)?1:0;

assign P3412=A2412;

ninexnine_unit ninexnine_unit_576(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20422)
);

ninexnine_unit ninexnine_unit_577(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21422)
);

ninexnine_unit ninexnine_unit_578(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22422)
);

ninexnine_unit ninexnine_unit_579(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23422)
);

ninexnine_unit ninexnine_unit_580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24422)
);

ninexnine_unit ninexnine_unit_581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25422)
);

ninexnine_unit ninexnine_unit_582(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26422)
);

ninexnine_unit ninexnine_unit_583(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27422)
);

assign C2422=c20422+c21422+c22422+c23422+c24422+c25422+c26422+c27422;
assign A2422=(C2422>=0)?1:0;

assign P3422=A2422;

ninexnine_unit ninexnine_unit_584(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20432)
);

ninexnine_unit ninexnine_unit_585(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21432)
);

ninexnine_unit ninexnine_unit_586(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22432)
);

ninexnine_unit ninexnine_unit_587(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23432)
);

ninexnine_unit ninexnine_unit_588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24432)
);

ninexnine_unit ninexnine_unit_589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25432)
);

ninexnine_unit ninexnine_unit_590(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26432)
);

ninexnine_unit ninexnine_unit_591(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27432)
);

assign C2432=c20432+c21432+c22432+c23432+c24432+c25432+c26432+c27432;
assign A2432=(C2432>=0)?1:0;

assign P3432=A2432;

ninexnine_unit ninexnine_unit_592(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20442)
);

ninexnine_unit ninexnine_unit_593(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21442)
);

ninexnine_unit ninexnine_unit_594(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22442)
);

ninexnine_unit ninexnine_unit_595(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23442)
);

ninexnine_unit ninexnine_unit_596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24442)
);

ninexnine_unit ninexnine_unit_597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25442)
);

ninexnine_unit ninexnine_unit_598(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26442)
);

ninexnine_unit ninexnine_unit_599(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27442)
);

assign C2442=c20442+c21442+c22442+c23442+c24442+c25442+c26442+c27442;
assign A2442=(C2442>=0)?1:0;

assign P3442=A2442;

ninexnine_unit ninexnine_unit_600(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20003)
);

ninexnine_unit ninexnine_unit_601(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21003)
);

ninexnine_unit ninexnine_unit_602(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22003)
);

ninexnine_unit ninexnine_unit_603(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23003)
);

ninexnine_unit ninexnine_unit_604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24003)
);

ninexnine_unit ninexnine_unit_605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25003)
);

ninexnine_unit ninexnine_unit_606(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26003)
);

ninexnine_unit ninexnine_unit_607(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27003)
);

assign C2003=c20003+c21003+c22003+c23003+c24003+c25003+c26003+c27003;
assign A2003=(C2003>=0)?1:0;

assign P3003=A2003;

ninexnine_unit ninexnine_unit_608(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20013)
);

ninexnine_unit ninexnine_unit_609(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21013)
);

ninexnine_unit ninexnine_unit_610(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22013)
);

ninexnine_unit ninexnine_unit_611(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23013)
);

ninexnine_unit ninexnine_unit_612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24013)
);

ninexnine_unit ninexnine_unit_613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25013)
);

ninexnine_unit ninexnine_unit_614(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26013)
);

ninexnine_unit ninexnine_unit_615(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27013)
);

assign C2013=c20013+c21013+c22013+c23013+c24013+c25013+c26013+c27013;
assign A2013=(C2013>=0)?1:0;

assign P3013=A2013;

ninexnine_unit ninexnine_unit_616(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20023)
);

ninexnine_unit ninexnine_unit_617(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21023)
);

ninexnine_unit ninexnine_unit_618(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22023)
);

ninexnine_unit ninexnine_unit_619(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23023)
);

ninexnine_unit ninexnine_unit_620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24023)
);

ninexnine_unit ninexnine_unit_621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25023)
);

ninexnine_unit ninexnine_unit_622(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26023)
);

ninexnine_unit ninexnine_unit_623(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27023)
);

assign C2023=c20023+c21023+c22023+c23023+c24023+c25023+c26023+c27023;
assign A2023=(C2023>=0)?1:0;

assign P3023=A2023;

ninexnine_unit ninexnine_unit_624(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20033)
);

ninexnine_unit ninexnine_unit_625(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21033)
);

ninexnine_unit ninexnine_unit_626(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22033)
);

ninexnine_unit ninexnine_unit_627(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23033)
);

ninexnine_unit ninexnine_unit_628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24033)
);

ninexnine_unit ninexnine_unit_629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25033)
);

ninexnine_unit ninexnine_unit_630(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26033)
);

ninexnine_unit ninexnine_unit_631(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27033)
);

assign C2033=c20033+c21033+c22033+c23033+c24033+c25033+c26033+c27033;
assign A2033=(C2033>=0)?1:0;

assign P3033=A2033;

ninexnine_unit ninexnine_unit_632(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20043)
);

ninexnine_unit ninexnine_unit_633(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21043)
);

ninexnine_unit ninexnine_unit_634(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22043)
);

ninexnine_unit ninexnine_unit_635(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23043)
);

ninexnine_unit ninexnine_unit_636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24043)
);

ninexnine_unit ninexnine_unit_637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25043)
);

ninexnine_unit ninexnine_unit_638(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26043)
);

ninexnine_unit ninexnine_unit_639(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27043)
);

assign C2043=c20043+c21043+c22043+c23043+c24043+c25043+c26043+c27043;
assign A2043=(C2043>=0)?1:0;

assign P3043=A2043;

ninexnine_unit ninexnine_unit_640(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20103)
);

ninexnine_unit ninexnine_unit_641(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21103)
);

ninexnine_unit ninexnine_unit_642(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22103)
);

ninexnine_unit ninexnine_unit_643(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23103)
);

ninexnine_unit ninexnine_unit_644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24103)
);

ninexnine_unit ninexnine_unit_645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25103)
);

ninexnine_unit ninexnine_unit_646(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26103)
);

ninexnine_unit ninexnine_unit_647(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27103)
);

assign C2103=c20103+c21103+c22103+c23103+c24103+c25103+c26103+c27103;
assign A2103=(C2103>=0)?1:0;

assign P3103=A2103;

ninexnine_unit ninexnine_unit_648(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20113)
);

ninexnine_unit ninexnine_unit_649(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21113)
);

ninexnine_unit ninexnine_unit_650(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22113)
);

ninexnine_unit ninexnine_unit_651(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23113)
);

ninexnine_unit ninexnine_unit_652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24113)
);

ninexnine_unit ninexnine_unit_653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25113)
);

ninexnine_unit ninexnine_unit_654(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26113)
);

ninexnine_unit ninexnine_unit_655(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27113)
);

assign C2113=c20113+c21113+c22113+c23113+c24113+c25113+c26113+c27113;
assign A2113=(C2113>=0)?1:0;

assign P3113=A2113;

ninexnine_unit ninexnine_unit_656(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20123)
);

ninexnine_unit ninexnine_unit_657(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21123)
);

ninexnine_unit ninexnine_unit_658(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22123)
);

ninexnine_unit ninexnine_unit_659(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23123)
);

ninexnine_unit ninexnine_unit_660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24123)
);

ninexnine_unit ninexnine_unit_661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25123)
);

ninexnine_unit ninexnine_unit_662(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26123)
);

ninexnine_unit ninexnine_unit_663(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27123)
);

assign C2123=c20123+c21123+c22123+c23123+c24123+c25123+c26123+c27123;
assign A2123=(C2123>=0)?1:0;

assign P3123=A2123;

ninexnine_unit ninexnine_unit_664(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20133)
);

ninexnine_unit ninexnine_unit_665(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21133)
);

ninexnine_unit ninexnine_unit_666(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22133)
);

ninexnine_unit ninexnine_unit_667(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23133)
);

ninexnine_unit ninexnine_unit_668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24133)
);

ninexnine_unit ninexnine_unit_669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25133)
);

ninexnine_unit ninexnine_unit_670(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26133)
);

ninexnine_unit ninexnine_unit_671(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27133)
);

assign C2133=c20133+c21133+c22133+c23133+c24133+c25133+c26133+c27133;
assign A2133=(C2133>=0)?1:0;

assign P3133=A2133;

ninexnine_unit ninexnine_unit_672(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20143)
);

ninexnine_unit ninexnine_unit_673(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21143)
);

ninexnine_unit ninexnine_unit_674(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22143)
);

ninexnine_unit ninexnine_unit_675(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23143)
);

ninexnine_unit ninexnine_unit_676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24143)
);

ninexnine_unit ninexnine_unit_677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25143)
);

ninexnine_unit ninexnine_unit_678(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26143)
);

ninexnine_unit ninexnine_unit_679(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27143)
);

assign C2143=c20143+c21143+c22143+c23143+c24143+c25143+c26143+c27143;
assign A2143=(C2143>=0)?1:0;

assign P3143=A2143;

ninexnine_unit ninexnine_unit_680(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20203)
);

ninexnine_unit ninexnine_unit_681(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21203)
);

ninexnine_unit ninexnine_unit_682(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22203)
);

ninexnine_unit ninexnine_unit_683(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23203)
);

ninexnine_unit ninexnine_unit_684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24203)
);

ninexnine_unit ninexnine_unit_685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25203)
);

ninexnine_unit ninexnine_unit_686(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26203)
);

ninexnine_unit ninexnine_unit_687(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27203)
);

assign C2203=c20203+c21203+c22203+c23203+c24203+c25203+c26203+c27203;
assign A2203=(C2203>=0)?1:0;

assign P3203=A2203;

ninexnine_unit ninexnine_unit_688(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20213)
);

ninexnine_unit ninexnine_unit_689(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21213)
);

ninexnine_unit ninexnine_unit_690(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22213)
);

ninexnine_unit ninexnine_unit_691(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23213)
);

ninexnine_unit ninexnine_unit_692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24213)
);

ninexnine_unit ninexnine_unit_693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25213)
);

ninexnine_unit ninexnine_unit_694(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26213)
);

ninexnine_unit ninexnine_unit_695(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27213)
);

assign C2213=c20213+c21213+c22213+c23213+c24213+c25213+c26213+c27213;
assign A2213=(C2213>=0)?1:0;

assign P3213=A2213;

ninexnine_unit ninexnine_unit_696(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20223)
);

ninexnine_unit ninexnine_unit_697(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21223)
);

ninexnine_unit ninexnine_unit_698(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22223)
);

ninexnine_unit ninexnine_unit_699(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23223)
);

ninexnine_unit ninexnine_unit_700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24223)
);

ninexnine_unit ninexnine_unit_701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25223)
);

ninexnine_unit ninexnine_unit_702(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26223)
);

ninexnine_unit ninexnine_unit_703(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27223)
);

assign C2223=c20223+c21223+c22223+c23223+c24223+c25223+c26223+c27223;
assign A2223=(C2223>=0)?1:0;

assign P3223=A2223;

ninexnine_unit ninexnine_unit_704(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20233)
);

ninexnine_unit ninexnine_unit_705(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21233)
);

ninexnine_unit ninexnine_unit_706(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22233)
);

ninexnine_unit ninexnine_unit_707(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23233)
);

ninexnine_unit ninexnine_unit_708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24233)
);

ninexnine_unit ninexnine_unit_709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25233)
);

ninexnine_unit ninexnine_unit_710(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26233)
);

ninexnine_unit ninexnine_unit_711(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27233)
);

assign C2233=c20233+c21233+c22233+c23233+c24233+c25233+c26233+c27233;
assign A2233=(C2233>=0)?1:0;

assign P3233=A2233;

ninexnine_unit ninexnine_unit_712(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20243)
);

ninexnine_unit ninexnine_unit_713(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21243)
);

ninexnine_unit ninexnine_unit_714(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22243)
);

ninexnine_unit ninexnine_unit_715(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23243)
);

ninexnine_unit ninexnine_unit_716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24243)
);

ninexnine_unit ninexnine_unit_717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25243)
);

ninexnine_unit ninexnine_unit_718(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26243)
);

ninexnine_unit ninexnine_unit_719(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27243)
);

assign C2243=c20243+c21243+c22243+c23243+c24243+c25243+c26243+c27243;
assign A2243=(C2243>=0)?1:0;

assign P3243=A2243;

ninexnine_unit ninexnine_unit_720(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20303)
);

ninexnine_unit ninexnine_unit_721(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21303)
);

ninexnine_unit ninexnine_unit_722(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22303)
);

ninexnine_unit ninexnine_unit_723(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23303)
);

ninexnine_unit ninexnine_unit_724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24303)
);

ninexnine_unit ninexnine_unit_725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25303)
);

ninexnine_unit ninexnine_unit_726(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26303)
);

ninexnine_unit ninexnine_unit_727(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27303)
);

assign C2303=c20303+c21303+c22303+c23303+c24303+c25303+c26303+c27303;
assign A2303=(C2303>=0)?1:0;

assign P3303=A2303;

ninexnine_unit ninexnine_unit_728(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20313)
);

ninexnine_unit ninexnine_unit_729(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21313)
);

ninexnine_unit ninexnine_unit_730(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22313)
);

ninexnine_unit ninexnine_unit_731(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23313)
);

ninexnine_unit ninexnine_unit_732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24313)
);

ninexnine_unit ninexnine_unit_733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25313)
);

ninexnine_unit ninexnine_unit_734(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26313)
);

ninexnine_unit ninexnine_unit_735(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27313)
);

assign C2313=c20313+c21313+c22313+c23313+c24313+c25313+c26313+c27313;
assign A2313=(C2313>=0)?1:0;

assign P3313=A2313;

ninexnine_unit ninexnine_unit_736(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20323)
);

ninexnine_unit ninexnine_unit_737(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21323)
);

ninexnine_unit ninexnine_unit_738(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22323)
);

ninexnine_unit ninexnine_unit_739(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23323)
);

ninexnine_unit ninexnine_unit_740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24323)
);

ninexnine_unit ninexnine_unit_741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25323)
);

ninexnine_unit ninexnine_unit_742(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26323)
);

ninexnine_unit ninexnine_unit_743(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27323)
);

assign C2323=c20323+c21323+c22323+c23323+c24323+c25323+c26323+c27323;
assign A2323=(C2323>=0)?1:0;

assign P3323=A2323;

ninexnine_unit ninexnine_unit_744(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20333)
);

ninexnine_unit ninexnine_unit_745(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21333)
);

ninexnine_unit ninexnine_unit_746(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22333)
);

ninexnine_unit ninexnine_unit_747(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23333)
);

ninexnine_unit ninexnine_unit_748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24333)
);

ninexnine_unit ninexnine_unit_749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25333)
);

ninexnine_unit ninexnine_unit_750(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26333)
);

ninexnine_unit ninexnine_unit_751(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27333)
);

assign C2333=c20333+c21333+c22333+c23333+c24333+c25333+c26333+c27333;
assign A2333=(C2333>=0)?1:0;

assign P3333=A2333;

ninexnine_unit ninexnine_unit_752(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20343)
);

ninexnine_unit ninexnine_unit_753(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21343)
);

ninexnine_unit ninexnine_unit_754(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22343)
);

ninexnine_unit ninexnine_unit_755(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23343)
);

ninexnine_unit ninexnine_unit_756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24343)
);

ninexnine_unit ninexnine_unit_757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25343)
);

ninexnine_unit ninexnine_unit_758(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26343)
);

ninexnine_unit ninexnine_unit_759(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27343)
);

assign C2343=c20343+c21343+c22343+c23343+c24343+c25343+c26343+c27343;
assign A2343=(C2343>=0)?1:0;

assign P3343=A2343;

ninexnine_unit ninexnine_unit_760(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20403)
);

ninexnine_unit ninexnine_unit_761(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21403)
);

ninexnine_unit ninexnine_unit_762(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22403)
);

ninexnine_unit ninexnine_unit_763(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23403)
);

ninexnine_unit ninexnine_unit_764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24403)
);

ninexnine_unit ninexnine_unit_765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25403)
);

ninexnine_unit ninexnine_unit_766(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26403)
);

ninexnine_unit ninexnine_unit_767(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27403)
);

assign C2403=c20403+c21403+c22403+c23403+c24403+c25403+c26403+c27403;
assign A2403=(C2403>=0)?1:0;

assign P3403=A2403;

ninexnine_unit ninexnine_unit_768(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20413)
);

ninexnine_unit ninexnine_unit_769(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21413)
);

ninexnine_unit ninexnine_unit_770(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22413)
);

ninexnine_unit ninexnine_unit_771(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23413)
);

ninexnine_unit ninexnine_unit_772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24413)
);

ninexnine_unit ninexnine_unit_773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25413)
);

ninexnine_unit ninexnine_unit_774(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26413)
);

ninexnine_unit ninexnine_unit_775(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27413)
);

assign C2413=c20413+c21413+c22413+c23413+c24413+c25413+c26413+c27413;
assign A2413=(C2413>=0)?1:0;

assign P3413=A2413;

ninexnine_unit ninexnine_unit_776(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20423)
);

ninexnine_unit ninexnine_unit_777(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21423)
);

ninexnine_unit ninexnine_unit_778(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22423)
);

ninexnine_unit ninexnine_unit_779(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23423)
);

ninexnine_unit ninexnine_unit_780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24423)
);

ninexnine_unit ninexnine_unit_781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25423)
);

ninexnine_unit ninexnine_unit_782(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26423)
);

ninexnine_unit ninexnine_unit_783(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27423)
);

assign C2423=c20423+c21423+c22423+c23423+c24423+c25423+c26423+c27423;
assign A2423=(C2423>=0)?1:0;

assign P3423=A2423;

ninexnine_unit ninexnine_unit_784(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20433)
);

ninexnine_unit ninexnine_unit_785(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21433)
);

ninexnine_unit ninexnine_unit_786(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22433)
);

ninexnine_unit ninexnine_unit_787(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23433)
);

ninexnine_unit ninexnine_unit_788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24433)
);

ninexnine_unit ninexnine_unit_789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25433)
);

ninexnine_unit ninexnine_unit_790(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26433)
);

ninexnine_unit ninexnine_unit_791(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27433)
);

assign C2433=c20433+c21433+c22433+c23433+c24433+c25433+c26433+c27433;
assign A2433=(C2433>=0)?1:0;

assign P3433=A2433;

ninexnine_unit ninexnine_unit_792(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20443)
);

ninexnine_unit ninexnine_unit_793(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21443)
);

ninexnine_unit ninexnine_unit_794(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22443)
);

ninexnine_unit ninexnine_unit_795(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23443)
);

ninexnine_unit ninexnine_unit_796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24443)
);

ninexnine_unit ninexnine_unit_797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25443)
);

ninexnine_unit ninexnine_unit_798(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26443)
);

ninexnine_unit ninexnine_unit_799(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27443)
);

assign C2443=c20443+c21443+c22443+c23443+c24443+c25443+c26443+c27443;
assign A2443=(C2443>=0)?1:0;

assign P3443=A2443;

ninexnine_unit ninexnine_unit_800(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20004)
);

ninexnine_unit ninexnine_unit_801(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21004)
);

ninexnine_unit ninexnine_unit_802(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22004)
);

ninexnine_unit ninexnine_unit_803(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23004)
);

ninexnine_unit ninexnine_unit_804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24004)
);

ninexnine_unit ninexnine_unit_805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25004)
);

ninexnine_unit ninexnine_unit_806(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26004)
);

ninexnine_unit ninexnine_unit_807(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27004)
);

assign C2004=c20004+c21004+c22004+c23004+c24004+c25004+c26004+c27004;
assign A2004=(C2004>=0)?1:0;

assign P3004=A2004;

ninexnine_unit ninexnine_unit_808(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20014)
);

ninexnine_unit ninexnine_unit_809(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21014)
);

ninexnine_unit ninexnine_unit_810(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22014)
);

ninexnine_unit ninexnine_unit_811(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23014)
);

ninexnine_unit ninexnine_unit_812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24014)
);

ninexnine_unit ninexnine_unit_813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25014)
);

ninexnine_unit ninexnine_unit_814(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26014)
);

ninexnine_unit ninexnine_unit_815(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27014)
);

assign C2014=c20014+c21014+c22014+c23014+c24014+c25014+c26014+c27014;
assign A2014=(C2014>=0)?1:0;

assign P3014=A2014;

ninexnine_unit ninexnine_unit_816(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20024)
);

ninexnine_unit ninexnine_unit_817(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21024)
);

ninexnine_unit ninexnine_unit_818(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22024)
);

ninexnine_unit ninexnine_unit_819(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23024)
);

ninexnine_unit ninexnine_unit_820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24024)
);

ninexnine_unit ninexnine_unit_821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25024)
);

ninexnine_unit ninexnine_unit_822(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26024)
);

ninexnine_unit ninexnine_unit_823(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27024)
);

assign C2024=c20024+c21024+c22024+c23024+c24024+c25024+c26024+c27024;
assign A2024=(C2024>=0)?1:0;

assign P3024=A2024;

ninexnine_unit ninexnine_unit_824(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20034)
);

ninexnine_unit ninexnine_unit_825(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21034)
);

ninexnine_unit ninexnine_unit_826(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22034)
);

ninexnine_unit ninexnine_unit_827(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23034)
);

ninexnine_unit ninexnine_unit_828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24034)
);

ninexnine_unit ninexnine_unit_829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25034)
);

ninexnine_unit ninexnine_unit_830(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26034)
);

ninexnine_unit ninexnine_unit_831(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27034)
);

assign C2034=c20034+c21034+c22034+c23034+c24034+c25034+c26034+c27034;
assign A2034=(C2034>=0)?1:0;

assign P3034=A2034;

ninexnine_unit ninexnine_unit_832(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20044)
);

ninexnine_unit ninexnine_unit_833(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21044)
);

ninexnine_unit ninexnine_unit_834(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22044)
);

ninexnine_unit ninexnine_unit_835(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23044)
);

ninexnine_unit ninexnine_unit_836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24044)
);

ninexnine_unit ninexnine_unit_837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25044)
);

ninexnine_unit ninexnine_unit_838(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26044)
);

ninexnine_unit ninexnine_unit_839(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27044)
);

assign C2044=c20044+c21044+c22044+c23044+c24044+c25044+c26044+c27044;
assign A2044=(C2044>=0)?1:0;

assign P3044=A2044;

ninexnine_unit ninexnine_unit_840(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20104)
);

ninexnine_unit ninexnine_unit_841(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21104)
);

ninexnine_unit ninexnine_unit_842(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22104)
);

ninexnine_unit ninexnine_unit_843(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23104)
);

ninexnine_unit ninexnine_unit_844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24104)
);

ninexnine_unit ninexnine_unit_845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25104)
);

ninexnine_unit ninexnine_unit_846(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26104)
);

ninexnine_unit ninexnine_unit_847(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27104)
);

assign C2104=c20104+c21104+c22104+c23104+c24104+c25104+c26104+c27104;
assign A2104=(C2104>=0)?1:0;

assign P3104=A2104;

ninexnine_unit ninexnine_unit_848(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20114)
);

ninexnine_unit ninexnine_unit_849(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21114)
);

ninexnine_unit ninexnine_unit_850(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22114)
);

ninexnine_unit ninexnine_unit_851(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23114)
);

ninexnine_unit ninexnine_unit_852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24114)
);

ninexnine_unit ninexnine_unit_853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25114)
);

ninexnine_unit ninexnine_unit_854(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26114)
);

ninexnine_unit ninexnine_unit_855(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27114)
);

assign C2114=c20114+c21114+c22114+c23114+c24114+c25114+c26114+c27114;
assign A2114=(C2114>=0)?1:0;

assign P3114=A2114;

ninexnine_unit ninexnine_unit_856(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20124)
);

ninexnine_unit ninexnine_unit_857(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21124)
);

ninexnine_unit ninexnine_unit_858(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22124)
);

ninexnine_unit ninexnine_unit_859(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23124)
);

ninexnine_unit ninexnine_unit_860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24124)
);

ninexnine_unit ninexnine_unit_861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25124)
);

ninexnine_unit ninexnine_unit_862(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26124)
);

ninexnine_unit ninexnine_unit_863(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27124)
);

assign C2124=c20124+c21124+c22124+c23124+c24124+c25124+c26124+c27124;
assign A2124=(C2124>=0)?1:0;

assign P3124=A2124;

ninexnine_unit ninexnine_unit_864(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20134)
);

ninexnine_unit ninexnine_unit_865(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21134)
);

ninexnine_unit ninexnine_unit_866(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22134)
);

ninexnine_unit ninexnine_unit_867(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23134)
);

ninexnine_unit ninexnine_unit_868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24134)
);

ninexnine_unit ninexnine_unit_869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25134)
);

ninexnine_unit ninexnine_unit_870(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26134)
);

ninexnine_unit ninexnine_unit_871(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27134)
);

assign C2134=c20134+c21134+c22134+c23134+c24134+c25134+c26134+c27134;
assign A2134=(C2134>=0)?1:0;

assign P3134=A2134;

ninexnine_unit ninexnine_unit_872(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20144)
);

ninexnine_unit ninexnine_unit_873(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21144)
);

ninexnine_unit ninexnine_unit_874(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22144)
);

ninexnine_unit ninexnine_unit_875(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23144)
);

ninexnine_unit ninexnine_unit_876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24144)
);

ninexnine_unit ninexnine_unit_877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25144)
);

ninexnine_unit ninexnine_unit_878(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26144)
);

ninexnine_unit ninexnine_unit_879(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27144)
);

assign C2144=c20144+c21144+c22144+c23144+c24144+c25144+c26144+c27144;
assign A2144=(C2144>=0)?1:0;

assign P3144=A2144;

ninexnine_unit ninexnine_unit_880(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20204)
);

ninexnine_unit ninexnine_unit_881(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21204)
);

ninexnine_unit ninexnine_unit_882(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22204)
);

ninexnine_unit ninexnine_unit_883(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23204)
);

ninexnine_unit ninexnine_unit_884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24204)
);

ninexnine_unit ninexnine_unit_885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25204)
);

ninexnine_unit ninexnine_unit_886(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26204)
);

ninexnine_unit ninexnine_unit_887(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27204)
);

assign C2204=c20204+c21204+c22204+c23204+c24204+c25204+c26204+c27204;
assign A2204=(C2204>=0)?1:0;

assign P3204=A2204;

ninexnine_unit ninexnine_unit_888(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20214)
);

ninexnine_unit ninexnine_unit_889(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21214)
);

ninexnine_unit ninexnine_unit_890(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22214)
);

ninexnine_unit ninexnine_unit_891(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23214)
);

ninexnine_unit ninexnine_unit_892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24214)
);

ninexnine_unit ninexnine_unit_893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25214)
);

ninexnine_unit ninexnine_unit_894(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26214)
);

ninexnine_unit ninexnine_unit_895(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27214)
);

assign C2214=c20214+c21214+c22214+c23214+c24214+c25214+c26214+c27214;
assign A2214=(C2214>=0)?1:0;

assign P3214=A2214;

ninexnine_unit ninexnine_unit_896(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20224)
);

ninexnine_unit ninexnine_unit_897(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21224)
);

ninexnine_unit ninexnine_unit_898(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22224)
);

ninexnine_unit ninexnine_unit_899(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23224)
);

ninexnine_unit ninexnine_unit_900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24224)
);

ninexnine_unit ninexnine_unit_901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25224)
);

ninexnine_unit ninexnine_unit_902(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26224)
);

ninexnine_unit ninexnine_unit_903(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27224)
);

assign C2224=c20224+c21224+c22224+c23224+c24224+c25224+c26224+c27224;
assign A2224=(C2224>=0)?1:0;

assign P3224=A2224;

ninexnine_unit ninexnine_unit_904(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20234)
);

ninexnine_unit ninexnine_unit_905(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21234)
);

ninexnine_unit ninexnine_unit_906(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22234)
);

ninexnine_unit ninexnine_unit_907(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23234)
);

ninexnine_unit ninexnine_unit_908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24234)
);

ninexnine_unit ninexnine_unit_909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25234)
);

ninexnine_unit ninexnine_unit_910(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26234)
);

ninexnine_unit ninexnine_unit_911(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27234)
);

assign C2234=c20234+c21234+c22234+c23234+c24234+c25234+c26234+c27234;
assign A2234=(C2234>=0)?1:0;

assign P3234=A2234;

ninexnine_unit ninexnine_unit_912(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20244)
);

ninexnine_unit ninexnine_unit_913(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21244)
);

ninexnine_unit ninexnine_unit_914(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22244)
);

ninexnine_unit ninexnine_unit_915(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23244)
);

ninexnine_unit ninexnine_unit_916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24244)
);

ninexnine_unit ninexnine_unit_917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25244)
);

ninexnine_unit ninexnine_unit_918(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26244)
);

ninexnine_unit ninexnine_unit_919(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27244)
);

assign C2244=c20244+c21244+c22244+c23244+c24244+c25244+c26244+c27244;
assign A2244=(C2244>=0)?1:0;

assign P3244=A2244;

ninexnine_unit ninexnine_unit_920(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20304)
);

ninexnine_unit ninexnine_unit_921(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21304)
);

ninexnine_unit ninexnine_unit_922(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22304)
);

ninexnine_unit ninexnine_unit_923(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23304)
);

ninexnine_unit ninexnine_unit_924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24304)
);

ninexnine_unit ninexnine_unit_925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25304)
);

ninexnine_unit ninexnine_unit_926(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26304)
);

ninexnine_unit ninexnine_unit_927(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27304)
);

assign C2304=c20304+c21304+c22304+c23304+c24304+c25304+c26304+c27304;
assign A2304=(C2304>=0)?1:0;

assign P3304=A2304;

ninexnine_unit ninexnine_unit_928(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20314)
);

ninexnine_unit ninexnine_unit_929(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21314)
);

ninexnine_unit ninexnine_unit_930(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22314)
);

ninexnine_unit ninexnine_unit_931(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23314)
);

ninexnine_unit ninexnine_unit_932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24314)
);

ninexnine_unit ninexnine_unit_933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25314)
);

ninexnine_unit ninexnine_unit_934(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26314)
);

ninexnine_unit ninexnine_unit_935(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27314)
);

assign C2314=c20314+c21314+c22314+c23314+c24314+c25314+c26314+c27314;
assign A2314=(C2314>=0)?1:0;

assign P3314=A2314;

ninexnine_unit ninexnine_unit_936(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20324)
);

ninexnine_unit ninexnine_unit_937(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21324)
);

ninexnine_unit ninexnine_unit_938(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22324)
);

ninexnine_unit ninexnine_unit_939(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23324)
);

ninexnine_unit ninexnine_unit_940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24324)
);

ninexnine_unit ninexnine_unit_941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25324)
);

ninexnine_unit ninexnine_unit_942(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26324)
);

ninexnine_unit ninexnine_unit_943(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27324)
);

assign C2324=c20324+c21324+c22324+c23324+c24324+c25324+c26324+c27324;
assign A2324=(C2324>=0)?1:0;

assign P3324=A2324;

ninexnine_unit ninexnine_unit_944(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20334)
);

ninexnine_unit ninexnine_unit_945(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21334)
);

ninexnine_unit ninexnine_unit_946(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22334)
);

ninexnine_unit ninexnine_unit_947(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23334)
);

ninexnine_unit ninexnine_unit_948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24334)
);

ninexnine_unit ninexnine_unit_949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25334)
);

ninexnine_unit ninexnine_unit_950(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26334)
);

ninexnine_unit ninexnine_unit_951(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27334)
);

assign C2334=c20334+c21334+c22334+c23334+c24334+c25334+c26334+c27334;
assign A2334=(C2334>=0)?1:0;

assign P3334=A2334;

ninexnine_unit ninexnine_unit_952(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20344)
);

ninexnine_unit ninexnine_unit_953(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21344)
);

ninexnine_unit ninexnine_unit_954(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22344)
);

ninexnine_unit ninexnine_unit_955(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23344)
);

ninexnine_unit ninexnine_unit_956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24344)
);

ninexnine_unit ninexnine_unit_957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25344)
);

ninexnine_unit ninexnine_unit_958(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26344)
);

ninexnine_unit ninexnine_unit_959(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27344)
);

assign C2344=c20344+c21344+c22344+c23344+c24344+c25344+c26344+c27344;
assign A2344=(C2344>=0)?1:0;

assign P3344=A2344;

ninexnine_unit ninexnine_unit_960(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20404)
);

ninexnine_unit ninexnine_unit_961(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21404)
);

ninexnine_unit ninexnine_unit_962(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22404)
);

ninexnine_unit ninexnine_unit_963(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23404)
);

ninexnine_unit ninexnine_unit_964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24404)
);

ninexnine_unit ninexnine_unit_965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25404)
);

ninexnine_unit ninexnine_unit_966(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26404)
);

ninexnine_unit ninexnine_unit_967(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27404)
);

assign C2404=c20404+c21404+c22404+c23404+c24404+c25404+c26404+c27404;
assign A2404=(C2404>=0)?1:0;

assign P3404=A2404;

ninexnine_unit ninexnine_unit_968(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20414)
);

ninexnine_unit ninexnine_unit_969(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21414)
);

ninexnine_unit ninexnine_unit_970(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22414)
);

ninexnine_unit ninexnine_unit_971(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23414)
);

ninexnine_unit ninexnine_unit_972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24414)
);

ninexnine_unit ninexnine_unit_973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25414)
);

ninexnine_unit ninexnine_unit_974(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26414)
);

ninexnine_unit ninexnine_unit_975(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27414)
);

assign C2414=c20414+c21414+c22414+c23414+c24414+c25414+c26414+c27414;
assign A2414=(C2414>=0)?1:0;

assign P3414=A2414;

ninexnine_unit ninexnine_unit_976(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20424)
);

ninexnine_unit ninexnine_unit_977(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21424)
);

ninexnine_unit ninexnine_unit_978(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22424)
);

ninexnine_unit ninexnine_unit_979(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23424)
);

ninexnine_unit ninexnine_unit_980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24424)
);

ninexnine_unit ninexnine_unit_981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25424)
);

ninexnine_unit ninexnine_unit_982(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26424)
);

ninexnine_unit ninexnine_unit_983(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27424)
);

assign C2424=c20424+c21424+c22424+c23424+c24424+c25424+c26424+c27424;
assign A2424=(C2424>=0)?1:0;

assign P3424=A2424;

ninexnine_unit ninexnine_unit_984(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20434)
);

ninexnine_unit ninexnine_unit_985(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21434)
);

ninexnine_unit ninexnine_unit_986(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22434)
);

ninexnine_unit ninexnine_unit_987(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23434)
);

ninexnine_unit ninexnine_unit_988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24434)
);

ninexnine_unit ninexnine_unit_989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25434)
);

ninexnine_unit ninexnine_unit_990(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26434)
);

ninexnine_unit ninexnine_unit_991(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27434)
);

assign C2434=c20434+c21434+c22434+c23434+c24434+c25434+c26434+c27434;
assign A2434=(C2434>=0)?1:0;

assign P3434=A2434;

ninexnine_unit ninexnine_unit_992(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20444)
);

ninexnine_unit ninexnine_unit_993(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21444)
);

ninexnine_unit ninexnine_unit_994(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22444)
);

ninexnine_unit ninexnine_unit_995(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23444)
);

ninexnine_unit ninexnine_unit_996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24444)
);

ninexnine_unit ninexnine_unit_997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25444)
);

ninexnine_unit ninexnine_unit_998(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26444)
);

ninexnine_unit ninexnine_unit_999(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27444)
);

assign C2444=c20444+c21444+c22444+c23444+c24444+c25444+c26444+c27444;
assign A2444=(C2444>=0)?1:0;

assign P3444=A2444;

ninexnine_unit ninexnine_unit_1000(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20005)
);

ninexnine_unit ninexnine_unit_1001(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21005)
);

ninexnine_unit ninexnine_unit_1002(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22005)
);

ninexnine_unit ninexnine_unit_1003(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23005)
);

ninexnine_unit ninexnine_unit_1004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24005)
);

ninexnine_unit ninexnine_unit_1005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25005)
);

ninexnine_unit ninexnine_unit_1006(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26005)
);

ninexnine_unit ninexnine_unit_1007(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27005)
);

assign C2005=c20005+c21005+c22005+c23005+c24005+c25005+c26005+c27005;
assign A2005=(C2005>=0)?1:0;

assign P3005=A2005;

ninexnine_unit ninexnine_unit_1008(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20015)
);

ninexnine_unit ninexnine_unit_1009(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21015)
);

ninexnine_unit ninexnine_unit_1010(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22015)
);

ninexnine_unit ninexnine_unit_1011(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23015)
);

ninexnine_unit ninexnine_unit_1012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24015)
);

ninexnine_unit ninexnine_unit_1013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25015)
);

ninexnine_unit ninexnine_unit_1014(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26015)
);

ninexnine_unit ninexnine_unit_1015(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27015)
);

assign C2015=c20015+c21015+c22015+c23015+c24015+c25015+c26015+c27015;
assign A2015=(C2015>=0)?1:0;

assign P3015=A2015;

ninexnine_unit ninexnine_unit_1016(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20025)
);

ninexnine_unit ninexnine_unit_1017(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21025)
);

ninexnine_unit ninexnine_unit_1018(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22025)
);

ninexnine_unit ninexnine_unit_1019(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23025)
);

ninexnine_unit ninexnine_unit_1020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24025)
);

ninexnine_unit ninexnine_unit_1021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25025)
);

ninexnine_unit ninexnine_unit_1022(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26025)
);

ninexnine_unit ninexnine_unit_1023(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27025)
);

assign C2025=c20025+c21025+c22025+c23025+c24025+c25025+c26025+c27025;
assign A2025=(C2025>=0)?1:0;

assign P3025=A2025;

ninexnine_unit ninexnine_unit_1024(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20035)
);

ninexnine_unit ninexnine_unit_1025(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21035)
);

ninexnine_unit ninexnine_unit_1026(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22035)
);

ninexnine_unit ninexnine_unit_1027(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23035)
);

ninexnine_unit ninexnine_unit_1028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24035)
);

ninexnine_unit ninexnine_unit_1029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25035)
);

ninexnine_unit ninexnine_unit_1030(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26035)
);

ninexnine_unit ninexnine_unit_1031(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27035)
);

assign C2035=c20035+c21035+c22035+c23035+c24035+c25035+c26035+c27035;
assign A2035=(C2035>=0)?1:0;

assign P3035=A2035;

ninexnine_unit ninexnine_unit_1032(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20045)
);

ninexnine_unit ninexnine_unit_1033(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21045)
);

ninexnine_unit ninexnine_unit_1034(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22045)
);

ninexnine_unit ninexnine_unit_1035(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23045)
);

ninexnine_unit ninexnine_unit_1036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24045)
);

ninexnine_unit ninexnine_unit_1037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25045)
);

ninexnine_unit ninexnine_unit_1038(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26045)
);

ninexnine_unit ninexnine_unit_1039(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27045)
);

assign C2045=c20045+c21045+c22045+c23045+c24045+c25045+c26045+c27045;
assign A2045=(C2045>=0)?1:0;

assign P3045=A2045;

ninexnine_unit ninexnine_unit_1040(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20105)
);

ninexnine_unit ninexnine_unit_1041(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21105)
);

ninexnine_unit ninexnine_unit_1042(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22105)
);

ninexnine_unit ninexnine_unit_1043(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23105)
);

ninexnine_unit ninexnine_unit_1044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24105)
);

ninexnine_unit ninexnine_unit_1045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25105)
);

ninexnine_unit ninexnine_unit_1046(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26105)
);

ninexnine_unit ninexnine_unit_1047(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27105)
);

assign C2105=c20105+c21105+c22105+c23105+c24105+c25105+c26105+c27105;
assign A2105=(C2105>=0)?1:0;

assign P3105=A2105;

ninexnine_unit ninexnine_unit_1048(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20115)
);

ninexnine_unit ninexnine_unit_1049(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21115)
);

ninexnine_unit ninexnine_unit_1050(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22115)
);

ninexnine_unit ninexnine_unit_1051(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23115)
);

ninexnine_unit ninexnine_unit_1052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24115)
);

ninexnine_unit ninexnine_unit_1053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25115)
);

ninexnine_unit ninexnine_unit_1054(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26115)
);

ninexnine_unit ninexnine_unit_1055(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27115)
);

assign C2115=c20115+c21115+c22115+c23115+c24115+c25115+c26115+c27115;
assign A2115=(C2115>=0)?1:0;

assign P3115=A2115;

ninexnine_unit ninexnine_unit_1056(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20125)
);

ninexnine_unit ninexnine_unit_1057(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21125)
);

ninexnine_unit ninexnine_unit_1058(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22125)
);

ninexnine_unit ninexnine_unit_1059(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23125)
);

ninexnine_unit ninexnine_unit_1060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24125)
);

ninexnine_unit ninexnine_unit_1061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25125)
);

ninexnine_unit ninexnine_unit_1062(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26125)
);

ninexnine_unit ninexnine_unit_1063(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27125)
);

assign C2125=c20125+c21125+c22125+c23125+c24125+c25125+c26125+c27125;
assign A2125=(C2125>=0)?1:0;

assign P3125=A2125;

ninexnine_unit ninexnine_unit_1064(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20135)
);

ninexnine_unit ninexnine_unit_1065(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21135)
);

ninexnine_unit ninexnine_unit_1066(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22135)
);

ninexnine_unit ninexnine_unit_1067(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23135)
);

ninexnine_unit ninexnine_unit_1068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24135)
);

ninexnine_unit ninexnine_unit_1069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25135)
);

ninexnine_unit ninexnine_unit_1070(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26135)
);

ninexnine_unit ninexnine_unit_1071(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27135)
);

assign C2135=c20135+c21135+c22135+c23135+c24135+c25135+c26135+c27135;
assign A2135=(C2135>=0)?1:0;

assign P3135=A2135;

ninexnine_unit ninexnine_unit_1072(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20145)
);

ninexnine_unit ninexnine_unit_1073(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21145)
);

ninexnine_unit ninexnine_unit_1074(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22145)
);

ninexnine_unit ninexnine_unit_1075(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23145)
);

ninexnine_unit ninexnine_unit_1076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24145)
);

ninexnine_unit ninexnine_unit_1077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25145)
);

ninexnine_unit ninexnine_unit_1078(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26145)
);

ninexnine_unit ninexnine_unit_1079(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27145)
);

assign C2145=c20145+c21145+c22145+c23145+c24145+c25145+c26145+c27145;
assign A2145=(C2145>=0)?1:0;

assign P3145=A2145;

ninexnine_unit ninexnine_unit_1080(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20205)
);

ninexnine_unit ninexnine_unit_1081(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21205)
);

ninexnine_unit ninexnine_unit_1082(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22205)
);

ninexnine_unit ninexnine_unit_1083(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23205)
);

ninexnine_unit ninexnine_unit_1084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24205)
);

ninexnine_unit ninexnine_unit_1085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25205)
);

ninexnine_unit ninexnine_unit_1086(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26205)
);

ninexnine_unit ninexnine_unit_1087(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27205)
);

assign C2205=c20205+c21205+c22205+c23205+c24205+c25205+c26205+c27205;
assign A2205=(C2205>=0)?1:0;

assign P3205=A2205;

ninexnine_unit ninexnine_unit_1088(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20215)
);

ninexnine_unit ninexnine_unit_1089(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21215)
);

ninexnine_unit ninexnine_unit_1090(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22215)
);

ninexnine_unit ninexnine_unit_1091(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23215)
);

ninexnine_unit ninexnine_unit_1092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24215)
);

ninexnine_unit ninexnine_unit_1093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25215)
);

ninexnine_unit ninexnine_unit_1094(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26215)
);

ninexnine_unit ninexnine_unit_1095(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27215)
);

assign C2215=c20215+c21215+c22215+c23215+c24215+c25215+c26215+c27215;
assign A2215=(C2215>=0)?1:0;

assign P3215=A2215;

ninexnine_unit ninexnine_unit_1096(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20225)
);

ninexnine_unit ninexnine_unit_1097(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21225)
);

ninexnine_unit ninexnine_unit_1098(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22225)
);

ninexnine_unit ninexnine_unit_1099(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23225)
);

ninexnine_unit ninexnine_unit_1100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24225)
);

ninexnine_unit ninexnine_unit_1101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25225)
);

ninexnine_unit ninexnine_unit_1102(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26225)
);

ninexnine_unit ninexnine_unit_1103(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27225)
);

assign C2225=c20225+c21225+c22225+c23225+c24225+c25225+c26225+c27225;
assign A2225=(C2225>=0)?1:0;

assign P3225=A2225;

ninexnine_unit ninexnine_unit_1104(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20235)
);

ninexnine_unit ninexnine_unit_1105(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21235)
);

ninexnine_unit ninexnine_unit_1106(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22235)
);

ninexnine_unit ninexnine_unit_1107(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23235)
);

ninexnine_unit ninexnine_unit_1108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24235)
);

ninexnine_unit ninexnine_unit_1109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25235)
);

ninexnine_unit ninexnine_unit_1110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26235)
);

ninexnine_unit ninexnine_unit_1111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27235)
);

assign C2235=c20235+c21235+c22235+c23235+c24235+c25235+c26235+c27235;
assign A2235=(C2235>=0)?1:0;

assign P3235=A2235;

ninexnine_unit ninexnine_unit_1112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20245)
);

ninexnine_unit ninexnine_unit_1113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21245)
);

ninexnine_unit ninexnine_unit_1114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22245)
);

ninexnine_unit ninexnine_unit_1115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23245)
);

ninexnine_unit ninexnine_unit_1116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24245)
);

ninexnine_unit ninexnine_unit_1117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25245)
);

ninexnine_unit ninexnine_unit_1118(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26245)
);

ninexnine_unit ninexnine_unit_1119(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27245)
);

assign C2245=c20245+c21245+c22245+c23245+c24245+c25245+c26245+c27245;
assign A2245=(C2245>=0)?1:0;

assign P3245=A2245;

ninexnine_unit ninexnine_unit_1120(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20305)
);

ninexnine_unit ninexnine_unit_1121(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21305)
);

ninexnine_unit ninexnine_unit_1122(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22305)
);

ninexnine_unit ninexnine_unit_1123(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23305)
);

ninexnine_unit ninexnine_unit_1124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24305)
);

ninexnine_unit ninexnine_unit_1125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25305)
);

ninexnine_unit ninexnine_unit_1126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26305)
);

ninexnine_unit ninexnine_unit_1127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27305)
);

assign C2305=c20305+c21305+c22305+c23305+c24305+c25305+c26305+c27305;
assign A2305=(C2305>=0)?1:0;

assign P3305=A2305;

ninexnine_unit ninexnine_unit_1128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20315)
);

ninexnine_unit ninexnine_unit_1129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21315)
);

ninexnine_unit ninexnine_unit_1130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22315)
);

ninexnine_unit ninexnine_unit_1131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23315)
);

ninexnine_unit ninexnine_unit_1132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24315)
);

ninexnine_unit ninexnine_unit_1133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25315)
);

ninexnine_unit ninexnine_unit_1134(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26315)
);

ninexnine_unit ninexnine_unit_1135(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27315)
);

assign C2315=c20315+c21315+c22315+c23315+c24315+c25315+c26315+c27315;
assign A2315=(C2315>=0)?1:0;

assign P3315=A2315;

ninexnine_unit ninexnine_unit_1136(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20325)
);

ninexnine_unit ninexnine_unit_1137(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21325)
);

ninexnine_unit ninexnine_unit_1138(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22325)
);

ninexnine_unit ninexnine_unit_1139(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23325)
);

ninexnine_unit ninexnine_unit_1140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24325)
);

ninexnine_unit ninexnine_unit_1141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25325)
);

ninexnine_unit ninexnine_unit_1142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26325)
);

ninexnine_unit ninexnine_unit_1143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27325)
);

assign C2325=c20325+c21325+c22325+c23325+c24325+c25325+c26325+c27325;
assign A2325=(C2325>=0)?1:0;

assign P3325=A2325;

ninexnine_unit ninexnine_unit_1144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20335)
);

ninexnine_unit ninexnine_unit_1145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21335)
);

ninexnine_unit ninexnine_unit_1146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22335)
);

ninexnine_unit ninexnine_unit_1147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23335)
);

ninexnine_unit ninexnine_unit_1148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24335)
);

ninexnine_unit ninexnine_unit_1149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25335)
);

ninexnine_unit ninexnine_unit_1150(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26335)
);

ninexnine_unit ninexnine_unit_1151(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27335)
);

assign C2335=c20335+c21335+c22335+c23335+c24335+c25335+c26335+c27335;
assign A2335=(C2335>=0)?1:0;

assign P3335=A2335;

ninexnine_unit ninexnine_unit_1152(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20345)
);

ninexnine_unit ninexnine_unit_1153(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21345)
);

ninexnine_unit ninexnine_unit_1154(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22345)
);

ninexnine_unit ninexnine_unit_1155(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23345)
);

ninexnine_unit ninexnine_unit_1156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24345)
);

ninexnine_unit ninexnine_unit_1157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25345)
);

ninexnine_unit ninexnine_unit_1158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26345)
);

ninexnine_unit ninexnine_unit_1159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27345)
);

assign C2345=c20345+c21345+c22345+c23345+c24345+c25345+c26345+c27345;
assign A2345=(C2345>=0)?1:0;

assign P3345=A2345;

ninexnine_unit ninexnine_unit_1160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20405)
);

ninexnine_unit ninexnine_unit_1161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21405)
);

ninexnine_unit ninexnine_unit_1162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22405)
);

ninexnine_unit ninexnine_unit_1163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23405)
);

ninexnine_unit ninexnine_unit_1164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24405)
);

ninexnine_unit ninexnine_unit_1165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25405)
);

ninexnine_unit ninexnine_unit_1166(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26405)
);

ninexnine_unit ninexnine_unit_1167(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27405)
);

assign C2405=c20405+c21405+c22405+c23405+c24405+c25405+c26405+c27405;
assign A2405=(C2405>=0)?1:0;

assign P3405=A2405;

ninexnine_unit ninexnine_unit_1168(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20415)
);

ninexnine_unit ninexnine_unit_1169(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21415)
);

ninexnine_unit ninexnine_unit_1170(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22415)
);

ninexnine_unit ninexnine_unit_1171(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23415)
);

ninexnine_unit ninexnine_unit_1172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24415)
);

ninexnine_unit ninexnine_unit_1173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25415)
);

ninexnine_unit ninexnine_unit_1174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26415)
);

ninexnine_unit ninexnine_unit_1175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27415)
);

assign C2415=c20415+c21415+c22415+c23415+c24415+c25415+c26415+c27415;
assign A2415=(C2415>=0)?1:0;

assign P3415=A2415;

ninexnine_unit ninexnine_unit_1176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20425)
);

ninexnine_unit ninexnine_unit_1177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21425)
);

ninexnine_unit ninexnine_unit_1178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22425)
);

ninexnine_unit ninexnine_unit_1179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23425)
);

ninexnine_unit ninexnine_unit_1180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24425)
);

ninexnine_unit ninexnine_unit_1181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25425)
);

ninexnine_unit ninexnine_unit_1182(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26425)
);

ninexnine_unit ninexnine_unit_1183(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27425)
);

assign C2425=c20425+c21425+c22425+c23425+c24425+c25425+c26425+c27425;
assign A2425=(C2425>=0)?1:0;

assign P3425=A2425;

ninexnine_unit ninexnine_unit_1184(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20435)
);

ninexnine_unit ninexnine_unit_1185(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21435)
);

ninexnine_unit ninexnine_unit_1186(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22435)
);

ninexnine_unit ninexnine_unit_1187(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23435)
);

ninexnine_unit ninexnine_unit_1188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24435)
);

ninexnine_unit ninexnine_unit_1189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25435)
);

ninexnine_unit ninexnine_unit_1190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26435)
);

ninexnine_unit ninexnine_unit_1191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27435)
);

assign C2435=c20435+c21435+c22435+c23435+c24435+c25435+c26435+c27435;
assign A2435=(C2435>=0)?1:0;

assign P3435=A2435;

ninexnine_unit ninexnine_unit_1192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20445)
);

ninexnine_unit ninexnine_unit_1193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21445)
);

ninexnine_unit ninexnine_unit_1194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22445)
);

ninexnine_unit ninexnine_unit_1195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23445)
);

ninexnine_unit ninexnine_unit_1196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24445)
);

ninexnine_unit ninexnine_unit_1197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25445)
);

ninexnine_unit ninexnine_unit_1198(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26445)
);

ninexnine_unit ninexnine_unit_1199(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27445)
);

assign C2445=c20445+c21445+c22445+c23445+c24445+c25445+c26445+c27445;
assign A2445=(C2445>=0)?1:0;

assign P3445=A2445;

ninexnine_unit ninexnine_unit_1200(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20006)
);

ninexnine_unit ninexnine_unit_1201(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21006)
);

ninexnine_unit ninexnine_unit_1202(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22006)
);

ninexnine_unit ninexnine_unit_1203(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23006)
);

ninexnine_unit ninexnine_unit_1204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24006)
);

ninexnine_unit ninexnine_unit_1205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25006)
);

ninexnine_unit ninexnine_unit_1206(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26006)
);

ninexnine_unit ninexnine_unit_1207(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27006)
);

assign C2006=c20006+c21006+c22006+c23006+c24006+c25006+c26006+c27006;
assign A2006=(C2006>=0)?1:0;

assign P3006=A2006;

ninexnine_unit ninexnine_unit_1208(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20016)
);

ninexnine_unit ninexnine_unit_1209(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21016)
);

ninexnine_unit ninexnine_unit_1210(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22016)
);

ninexnine_unit ninexnine_unit_1211(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23016)
);

ninexnine_unit ninexnine_unit_1212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24016)
);

ninexnine_unit ninexnine_unit_1213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25016)
);

ninexnine_unit ninexnine_unit_1214(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26016)
);

ninexnine_unit ninexnine_unit_1215(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27016)
);

assign C2016=c20016+c21016+c22016+c23016+c24016+c25016+c26016+c27016;
assign A2016=(C2016>=0)?1:0;

assign P3016=A2016;

ninexnine_unit ninexnine_unit_1216(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20026)
);

ninexnine_unit ninexnine_unit_1217(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21026)
);

ninexnine_unit ninexnine_unit_1218(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22026)
);

ninexnine_unit ninexnine_unit_1219(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23026)
);

ninexnine_unit ninexnine_unit_1220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24026)
);

ninexnine_unit ninexnine_unit_1221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25026)
);

ninexnine_unit ninexnine_unit_1222(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26026)
);

ninexnine_unit ninexnine_unit_1223(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27026)
);

assign C2026=c20026+c21026+c22026+c23026+c24026+c25026+c26026+c27026;
assign A2026=(C2026>=0)?1:0;

assign P3026=A2026;

ninexnine_unit ninexnine_unit_1224(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20036)
);

ninexnine_unit ninexnine_unit_1225(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21036)
);

ninexnine_unit ninexnine_unit_1226(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22036)
);

ninexnine_unit ninexnine_unit_1227(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23036)
);

ninexnine_unit ninexnine_unit_1228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24036)
);

ninexnine_unit ninexnine_unit_1229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25036)
);

ninexnine_unit ninexnine_unit_1230(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26036)
);

ninexnine_unit ninexnine_unit_1231(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27036)
);

assign C2036=c20036+c21036+c22036+c23036+c24036+c25036+c26036+c27036;
assign A2036=(C2036>=0)?1:0;

assign P3036=A2036;

ninexnine_unit ninexnine_unit_1232(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20046)
);

ninexnine_unit ninexnine_unit_1233(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21046)
);

ninexnine_unit ninexnine_unit_1234(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22046)
);

ninexnine_unit ninexnine_unit_1235(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23046)
);

ninexnine_unit ninexnine_unit_1236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24046)
);

ninexnine_unit ninexnine_unit_1237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25046)
);

ninexnine_unit ninexnine_unit_1238(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26046)
);

ninexnine_unit ninexnine_unit_1239(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27046)
);

assign C2046=c20046+c21046+c22046+c23046+c24046+c25046+c26046+c27046;
assign A2046=(C2046>=0)?1:0;

assign P3046=A2046;

ninexnine_unit ninexnine_unit_1240(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20106)
);

ninexnine_unit ninexnine_unit_1241(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21106)
);

ninexnine_unit ninexnine_unit_1242(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22106)
);

ninexnine_unit ninexnine_unit_1243(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23106)
);

ninexnine_unit ninexnine_unit_1244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24106)
);

ninexnine_unit ninexnine_unit_1245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25106)
);

ninexnine_unit ninexnine_unit_1246(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26106)
);

ninexnine_unit ninexnine_unit_1247(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27106)
);

assign C2106=c20106+c21106+c22106+c23106+c24106+c25106+c26106+c27106;
assign A2106=(C2106>=0)?1:0;

assign P3106=A2106;

ninexnine_unit ninexnine_unit_1248(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20116)
);

ninexnine_unit ninexnine_unit_1249(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21116)
);

ninexnine_unit ninexnine_unit_1250(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22116)
);

ninexnine_unit ninexnine_unit_1251(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23116)
);

ninexnine_unit ninexnine_unit_1252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24116)
);

ninexnine_unit ninexnine_unit_1253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25116)
);

ninexnine_unit ninexnine_unit_1254(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26116)
);

ninexnine_unit ninexnine_unit_1255(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27116)
);

assign C2116=c20116+c21116+c22116+c23116+c24116+c25116+c26116+c27116;
assign A2116=(C2116>=0)?1:0;

assign P3116=A2116;

ninexnine_unit ninexnine_unit_1256(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20126)
);

ninexnine_unit ninexnine_unit_1257(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21126)
);

ninexnine_unit ninexnine_unit_1258(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22126)
);

ninexnine_unit ninexnine_unit_1259(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23126)
);

ninexnine_unit ninexnine_unit_1260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24126)
);

ninexnine_unit ninexnine_unit_1261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25126)
);

ninexnine_unit ninexnine_unit_1262(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26126)
);

ninexnine_unit ninexnine_unit_1263(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27126)
);

assign C2126=c20126+c21126+c22126+c23126+c24126+c25126+c26126+c27126;
assign A2126=(C2126>=0)?1:0;

assign P3126=A2126;

ninexnine_unit ninexnine_unit_1264(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20136)
);

ninexnine_unit ninexnine_unit_1265(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21136)
);

ninexnine_unit ninexnine_unit_1266(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22136)
);

ninexnine_unit ninexnine_unit_1267(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23136)
);

ninexnine_unit ninexnine_unit_1268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24136)
);

ninexnine_unit ninexnine_unit_1269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25136)
);

ninexnine_unit ninexnine_unit_1270(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26136)
);

ninexnine_unit ninexnine_unit_1271(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27136)
);

assign C2136=c20136+c21136+c22136+c23136+c24136+c25136+c26136+c27136;
assign A2136=(C2136>=0)?1:0;

assign P3136=A2136;

ninexnine_unit ninexnine_unit_1272(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20146)
);

ninexnine_unit ninexnine_unit_1273(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21146)
);

ninexnine_unit ninexnine_unit_1274(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22146)
);

ninexnine_unit ninexnine_unit_1275(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23146)
);

ninexnine_unit ninexnine_unit_1276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24146)
);

ninexnine_unit ninexnine_unit_1277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25146)
);

ninexnine_unit ninexnine_unit_1278(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26146)
);

ninexnine_unit ninexnine_unit_1279(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27146)
);

assign C2146=c20146+c21146+c22146+c23146+c24146+c25146+c26146+c27146;
assign A2146=(C2146>=0)?1:0;

assign P3146=A2146;

ninexnine_unit ninexnine_unit_1280(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20206)
);

ninexnine_unit ninexnine_unit_1281(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21206)
);

ninexnine_unit ninexnine_unit_1282(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22206)
);

ninexnine_unit ninexnine_unit_1283(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23206)
);

ninexnine_unit ninexnine_unit_1284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24206)
);

ninexnine_unit ninexnine_unit_1285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25206)
);

ninexnine_unit ninexnine_unit_1286(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26206)
);

ninexnine_unit ninexnine_unit_1287(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27206)
);

assign C2206=c20206+c21206+c22206+c23206+c24206+c25206+c26206+c27206;
assign A2206=(C2206>=0)?1:0;

assign P3206=A2206;

ninexnine_unit ninexnine_unit_1288(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20216)
);

ninexnine_unit ninexnine_unit_1289(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21216)
);

ninexnine_unit ninexnine_unit_1290(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22216)
);

ninexnine_unit ninexnine_unit_1291(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23216)
);

ninexnine_unit ninexnine_unit_1292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24216)
);

ninexnine_unit ninexnine_unit_1293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25216)
);

ninexnine_unit ninexnine_unit_1294(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26216)
);

ninexnine_unit ninexnine_unit_1295(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27216)
);

assign C2216=c20216+c21216+c22216+c23216+c24216+c25216+c26216+c27216;
assign A2216=(C2216>=0)?1:0;

assign P3216=A2216;

ninexnine_unit ninexnine_unit_1296(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20226)
);

ninexnine_unit ninexnine_unit_1297(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21226)
);

ninexnine_unit ninexnine_unit_1298(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22226)
);

ninexnine_unit ninexnine_unit_1299(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23226)
);

ninexnine_unit ninexnine_unit_1300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24226)
);

ninexnine_unit ninexnine_unit_1301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25226)
);

ninexnine_unit ninexnine_unit_1302(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26226)
);

ninexnine_unit ninexnine_unit_1303(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27226)
);

assign C2226=c20226+c21226+c22226+c23226+c24226+c25226+c26226+c27226;
assign A2226=(C2226>=0)?1:0;

assign P3226=A2226;

ninexnine_unit ninexnine_unit_1304(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20236)
);

ninexnine_unit ninexnine_unit_1305(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21236)
);

ninexnine_unit ninexnine_unit_1306(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22236)
);

ninexnine_unit ninexnine_unit_1307(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23236)
);

ninexnine_unit ninexnine_unit_1308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24236)
);

ninexnine_unit ninexnine_unit_1309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25236)
);

ninexnine_unit ninexnine_unit_1310(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26236)
);

ninexnine_unit ninexnine_unit_1311(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27236)
);

assign C2236=c20236+c21236+c22236+c23236+c24236+c25236+c26236+c27236;
assign A2236=(C2236>=0)?1:0;

assign P3236=A2236;

ninexnine_unit ninexnine_unit_1312(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20246)
);

ninexnine_unit ninexnine_unit_1313(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21246)
);

ninexnine_unit ninexnine_unit_1314(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22246)
);

ninexnine_unit ninexnine_unit_1315(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23246)
);

ninexnine_unit ninexnine_unit_1316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24246)
);

ninexnine_unit ninexnine_unit_1317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25246)
);

ninexnine_unit ninexnine_unit_1318(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26246)
);

ninexnine_unit ninexnine_unit_1319(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27246)
);

assign C2246=c20246+c21246+c22246+c23246+c24246+c25246+c26246+c27246;
assign A2246=(C2246>=0)?1:0;

assign P3246=A2246;

ninexnine_unit ninexnine_unit_1320(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20306)
);

ninexnine_unit ninexnine_unit_1321(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21306)
);

ninexnine_unit ninexnine_unit_1322(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22306)
);

ninexnine_unit ninexnine_unit_1323(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23306)
);

ninexnine_unit ninexnine_unit_1324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24306)
);

ninexnine_unit ninexnine_unit_1325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25306)
);

ninexnine_unit ninexnine_unit_1326(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26306)
);

ninexnine_unit ninexnine_unit_1327(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27306)
);

assign C2306=c20306+c21306+c22306+c23306+c24306+c25306+c26306+c27306;
assign A2306=(C2306>=0)?1:0;

assign P3306=A2306;

ninexnine_unit ninexnine_unit_1328(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20316)
);

ninexnine_unit ninexnine_unit_1329(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21316)
);

ninexnine_unit ninexnine_unit_1330(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22316)
);

ninexnine_unit ninexnine_unit_1331(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23316)
);

ninexnine_unit ninexnine_unit_1332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24316)
);

ninexnine_unit ninexnine_unit_1333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25316)
);

ninexnine_unit ninexnine_unit_1334(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26316)
);

ninexnine_unit ninexnine_unit_1335(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27316)
);

assign C2316=c20316+c21316+c22316+c23316+c24316+c25316+c26316+c27316;
assign A2316=(C2316>=0)?1:0;

assign P3316=A2316;

ninexnine_unit ninexnine_unit_1336(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20326)
);

ninexnine_unit ninexnine_unit_1337(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21326)
);

ninexnine_unit ninexnine_unit_1338(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22326)
);

ninexnine_unit ninexnine_unit_1339(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23326)
);

ninexnine_unit ninexnine_unit_1340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24326)
);

ninexnine_unit ninexnine_unit_1341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25326)
);

ninexnine_unit ninexnine_unit_1342(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26326)
);

ninexnine_unit ninexnine_unit_1343(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27326)
);

assign C2326=c20326+c21326+c22326+c23326+c24326+c25326+c26326+c27326;
assign A2326=(C2326>=0)?1:0;

assign P3326=A2326;

ninexnine_unit ninexnine_unit_1344(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20336)
);

ninexnine_unit ninexnine_unit_1345(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21336)
);

ninexnine_unit ninexnine_unit_1346(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22336)
);

ninexnine_unit ninexnine_unit_1347(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23336)
);

ninexnine_unit ninexnine_unit_1348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24336)
);

ninexnine_unit ninexnine_unit_1349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25336)
);

ninexnine_unit ninexnine_unit_1350(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26336)
);

ninexnine_unit ninexnine_unit_1351(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27336)
);

assign C2336=c20336+c21336+c22336+c23336+c24336+c25336+c26336+c27336;
assign A2336=(C2336>=0)?1:0;

assign P3336=A2336;

ninexnine_unit ninexnine_unit_1352(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20346)
);

ninexnine_unit ninexnine_unit_1353(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21346)
);

ninexnine_unit ninexnine_unit_1354(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22346)
);

ninexnine_unit ninexnine_unit_1355(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23346)
);

ninexnine_unit ninexnine_unit_1356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24346)
);

ninexnine_unit ninexnine_unit_1357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25346)
);

ninexnine_unit ninexnine_unit_1358(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26346)
);

ninexnine_unit ninexnine_unit_1359(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27346)
);

assign C2346=c20346+c21346+c22346+c23346+c24346+c25346+c26346+c27346;
assign A2346=(C2346>=0)?1:0;

assign P3346=A2346;

ninexnine_unit ninexnine_unit_1360(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20406)
);

ninexnine_unit ninexnine_unit_1361(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21406)
);

ninexnine_unit ninexnine_unit_1362(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22406)
);

ninexnine_unit ninexnine_unit_1363(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23406)
);

ninexnine_unit ninexnine_unit_1364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24406)
);

ninexnine_unit ninexnine_unit_1365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25406)
);

ninexnine_unit ninexnine_unit_1366(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26406)
);

ninexnine_unit ninexnine_unit_1367(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27406)
);

assign C2406=c20406+c21406+c22406+c23406+c24406+c25406+c26406+c27406;
assign A2406=(C2406>=0)?1:0;

assign P3406=A2406;

ninexnine_unit ninexnine_unit_1368(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20416)
);

ninexnine_unit ninexnine_unit_1369(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21416)
);

ninexnine_unit ninexnine_unit_1370(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22416)
);

ninexnine_unit ninexnine_unit_1371(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23416)
);

ninexnine_unit ninexnine_unit_1372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24416)
);

ninexnine_unit ninexnine_unit_1373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25416)
);

ninexnine_unit ninexnine_unit_1374(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26416)
);

ninexnine_unit ninexnine_unit_1375(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27416)
);

assign C2416=c20416+c21416+c22416+c23416+c24416+c25416+c26416+c27416;
assign A2416=(C2416>=0)?1:0;

assign P3416=A2416;

ninexnine_unit ninexnine_unit_1376(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20426)
);

ninexnine_unit ninexnine_unit_1377(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21426)
);

ninexnine_unit ninexnine_unit_1378(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22426)
);

ninexnine_unit ninexnine_unit_1379(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23426)
);

ninexnine_unit ninexnine_unit_1380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24426)
);

ninexnine_unit ninexnine_unit_1381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25426)
);

ninexnine_unit ninexnine_unit_1382(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26426)
);

ninexnine_unit ninexnine_unit_1383(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27426)
);

assign C2426=c20426+c21426+c22426+c23426+c24426+c25426+c26426+c27426;
assign A2426=(C2426>=0)?1:0;

assign P3426=A2426;

ninexnine_unit ninexnine_unit_1384(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20436)
);

ninexnine_unit ninexnine_unit_1385(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21436)
);

ninexnine_unit ninexnine_unit_1386(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22436)
);

ninexnine_unit ninexnine_unit_1387(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23436)
);

ninexnine_unit ninexnine_unit_1388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24436)
);

ninexnine_unit ninexnine_unit_1389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25436)
);

ninexnine_unit ninexnine_unit_1390(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26436)
);

ninexnine_unit ninexnine_unit_1391(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27436)
);

assign C2436=c20436+c21436+c22436+c23436+c24436+c25436+c26436+c27436;
assign A2436=(C2436>=0)?1:0;

assign P3436=A2436;

ninexnine_unit ninexnine_unit_1392(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20446)
);

ninexnine_unit ninexnine_unit_1393(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21446)
);

ninexnine_unit ninexnine_unit_1394(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22446)
);

ninexnine_unit ninexnine_unit_1395(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23446)
);

ninexnine_unit ninexnine_unit_1396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24446)
);

ninexnine_unit ninexnine_unit_1397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25446)
);

ninexnine_unit ninexnine_unit_1398(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26446)
);

ninexnine_unit ninexnine_unit_1399(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27446)
);

assign C2446=c20446+c21446+c22446+c23446+c24446+c25446+c26446+c27446;
assign A2446=(C2446>=0)?1:0;

assign P3446=A2446;

ninexnine_unit ninexnine_unit_1400(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20007)
);

ninexnine_unit ninexnine_unit_1401(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21007)
);

ninexnine_unit ninexnine_unit_1402(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22007)
);

ninexnine_unit ninexnine_unit_1403(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23007)
);

ninexnine_unit ninexnine_unit_1404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24007)
);

ninexnine_unit ninexnine_unit_1405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25007)
);

ninexnine_unit ninexnine_unit_1406(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26007)
);

ninexnine_unit ninexnine_unit_1407(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27007)
);

assign C2007=c20007+c21007+c22007+c23007+c24007+c25007+c26007+c27007;
assign A2007=(C2007>=0)?1:0;

assign P3007=A2007;

ninexnine_unit ninexnine_unit_1408(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20017)
);

ninexnine_unit ninexnine_unit_1409(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21017)
);

ninexnine_unit ninexnine_unit_1410(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22017)
);

ninexnine_unit ninexnine_unit_1411(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23017)
);

ninexnine_unit ninexnine_unit_1412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24017)
);

ninexnine_unit ninexnine_unit_1413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25017)
);

ninexnine_unit ninexnine_unit_1414(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26017)
);

ninexnine_unit ninexnine_unit_1415(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27017)
);

assign C2017=c20017+c21017+c22017+c23017+c24017+c25017+c26017+c27017;
assign A2017=(C2017>=0)?1:0;

assign P3017=A2017;

ninexnine_unit ninexnine_unit_1416(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20027)
);

ninexnine_unit ninexnine_unit_1417(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21027)
);

ninexnine_unit ninexnine_unit_1418(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22027)
);

ninexnine_unit ninexnine_unit_1419(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23027)
);

ninexnine_unit ninexnine_unit_1420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24027)
);

ninexnine_unit ninexnine_unit_1421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25027)
);

ninexnine_unit ninexnine_unit_1422(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26027)
);

ninexnine_unit ninexnine_unit_1423(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27027)
);

assign C2027=c20027+c21027+c22027+c23027+c24027+c25027+c26027+c27027;
assign A2027=(C2027>=0)?1:0;

assign P3027=A2027;

ninexnine_unit ninexnine_unit_1424(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20037)
);

ninexnine_unit ninexnine_unit_1425(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21037)
);

ninexnine_unit ninexnine_unit_1426(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22037)
);

ninexnine_unit ninexnine_unit_1427(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23037)
);

ninexnine_unit ninexnine_unit_1428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24037)
);

ninexnine_unit ninexnine_unit_1429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25037)
);

ninexnine_unit ninexnine_unit_1430(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26037)
);

ninexnine_unit ninexnine_unit_1431(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27037)
);

assign C2037=c20037+c21037+c22037+c23037+c24037+c25037+c26037+c27037;
assign A2037=(C2037>=0)?1:0;

assign P3037=A2037;

ninexnine_unit ninexnine_unit_1432(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20047)
);

ninexnine_unit ninexnine_unit_1433(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21047)
);

ninexnine_unit ninexnine_unit_1434(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22047)
);

ninexnine_unit ninexnine_unit_1435(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23047)
);

ninexnine_unit ninexnine_unit_1436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24047)
);

ninexnine_unit ninexnine_unit_1437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25047)
);

ninexnine_unit ninexnine_unit_1438(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26047)
);

ninexnine_unit ninexnine_unit_1439(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27047)
);

assign C2047=c20047+c21047+c22047+c23047+c24047+c25047+c26047+c27047;
assign A2047=(C2047>=0)?1:0;

assign P3047=A2047;

ninexnine_unit ninexnine_unit_1440(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20107)
);

ninexnine_unit ninexnine_unit_1441(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21107)
);

ninexnine_unit ninexnine_unit_1442(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22107)
);

ninexnine_unit ninexnine_unit_1443(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23107)
);

ninexnine_unit ninexnine_unit_1444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24107)
);

ninexnine_unit ninexnine_unit_1445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25107)
);

ninexnine_unit ninexnine_unit_1446(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26107)
);

ninexnine_unit ninexnine_unit_1447(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27107)
);

assign C2107=c20107+c21107+c22107+c23107+c24107+c25107+c26107+c27107;
assign A2107=(C2107>=0)?1:0;

assign P3107=A2107;

ninexnine_unit ninexnine_unit_1448(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20117)
);

ninexnine_unit ninexnine_unit_1449(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21117)
);

ninexnine_unit ninexnine_unit_1450(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22117)
);

ninexnine_unit ninexnine_unit_1451(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23117)
);

ninexnine_unit ninexnine_unit_1452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24117)
);

ninexnine_unit ninexnine_unit_1453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25117)
);

ninexnine_unit ninexnine_unit_1454(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26117)
);

ninexnine_unit ninexnine_unit_1455(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27117)
);

assign C2117=c20117+c21117+c22117+c23117+c24117+c25117+c26117+c27117;
assign A2117=(C2117>=0)?1:0;

assign P3117=A2117;

ninexnine_unit ninexnine_unit_1456(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20127)
);

ninexnine_unit ninexnine_unit_1457(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21127)
);

ninexnine_unit ninexnine_unit_1458(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22127)
);

ninexnine_unit ninexnine_unit_1459(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23127)
);

ninexnine_unit ninexnine_unit_1460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24127)
);

ninexnine_unit ninexnine_unit_1461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25127)
);

ninexnine_unit ninexnine_unit_1462(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26127)
);

ninexnine_unit ninexnine_unit_1463(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27127)
);

assign C2127=c20127+c21127+c22127+c23127+c24127+c25127+c26127+c27127;
assign A2127=(C2127>=0)?1:0;

assign P3127=A2127;

ninexnine_unit ninexnine_unit_1464(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20137)
);

ninexnine_unit ninexnine_unit_1465(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21137)
);

ninexnine_unit ninexnine_unit_1466(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22137)
);

ninexnine_unit ninexnine_unit_1467(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23137)
);

ninexnine_unit ninexnine_unit_1468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24137)
);

ninexnine_unit ninexnine_unit_1469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25137)
);

ninexnine_unit ninexnine_unit_1470(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26137)
);

ninexnine_unit ninexnine_unit_1471(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27137)
);

assign C2137=c20137+c21137+c22137+c23137+c24137+c25137+c26137+c27137;
assign A2137=(C2137>=0)?1:0;

assign P3137=A2137;

ninexnine_unit ninexnine_unit_1472(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20147)
);

ninexnine_unit ninexnine_unit_1473(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21147)
);

ninexnine_unit ninexnine_unit_1474(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22147)
);

ninexnine_unit ninexnine_unit_1475(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23147)
);

ninexnine_unit ninexnine_unit_1476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24147)
);

ninexnine_unit ninexnine_unit_1477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25147)
);

ninexnine_unit ninexnine_unit_1478(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26147)
);

ninexnine_unit ninexnine_unit_1479(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27147)
);

assign C2147=c20147+c21147+c22147+c23147+c24147+c25147+c26147+c27147;
assign A2147=(C2147>=0)?1:0;

assign P3147=A2147;

ninexnine_unit ninexnine_unit_1480(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20207)
);

ninexnine_unit ninexnine_unit_1481(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21207)
);

ninexnine_unit ninexnine_unit_1482(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22207)
);

ninexnine_unit ninexnine_unit_1483(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23207)
);

ninexnine_unit ninexnine_unit_1484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24207)
);

ninexnine_unit ninexnine_unit_1485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25207)
);

ninexnine_unit ninexnine_unit_1486(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26207)
);

ninexnine_unit ninexnine_unit_1487(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27207)
);

assign C2207=c20207+c21207+c22207+c23207+c24207+c25207+c26207+c27207;
assign A2207=(C2207>=0)?1:0;

assign P3207=A2207;

ninexnine_unit ninexnine_unit_1488(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20217)
);

ninexnine_unit ninexnine_unit_1489(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21217)
);

ninexnine_unit ninexnine_unit_1490(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22217)
);

ninexnine_unit ninexnine_unit_1491(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23217)
);

ninexnine_unit ninexnine_unit_1492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24217)
);

ninexnine_unit ninexnine_unit_1493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25217)
);

ninexnine_unit ninexnine_unit_1494(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26217)
);

ninexnine_unit ninexnine_unit_1495(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27217)
);

assign C2217=c20217+c21217+c22217+c23217+c24217+c25217+c26217+c27217;
assign A2217=(C2217>=0)?1:0;

assign P3217=A2217;

ninexnine_unit ninexnine_unit_1496(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20227)
);

ninexnine_unit ninexnine_unit_1497(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21227)
);

ninexnine_unit ninexnine_unit_1498(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22227)
);

ninexnine_unit ninexnine_unit_1499(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23227)
);

ninexnine_unit ninexnine_unit_1500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24227)
);

ninexnine_unit ninexnine_unit_1501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25227)
);

ninexnine_unit ninexnine_unit_1502(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26227)
);

ninexnine_unit ninexnine_unit_1503(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27227)
);

assign C2227=c20227+c21227+c22227+c23227+c24227+c25227+c26227+c27227;
assign A2227=(C2227>=0)?1:0;

assign P3227=A2227;

ninexnine_unit ninexnine_unit_1504(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20237)
);

ninexnine_unit ninexnine_unit_1505(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21237)
);

ninexnine_unit ninexnine_unit_1506(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22237)
);

ninexnine_unit ninexnine_unit_1507(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23237)
);

ninexnine_unit ninexnine_unit_1508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24237)
);

ninexnine_unit ninexnine_unit_1509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25237)
);

ninexnine_unit ninexnine_unit_1510(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26237)
);

ninexnine_unit ninexnine_unit_1511(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27237)
);

assign C2237=c20237+c21237+c22237+c23237+c24237+c25237+c26237+c27237;
assign A2237=(C2237>=0)?1:0;

assign P3237=A2237;

ninexnine_unit ninexnine_unit_1512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20247)
);

ninexnine_unit ninexnine_unit_1513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21247)
);

ninexnine_unit ninexnine_unit_1514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22247)
);

ninexnine_unit ninexnine_unit_1515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23247)
);

ninexnine_unit ninexnine_unit_1516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24247)
);

ninexnine_unit ninexnine_unit_1517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25247)
);

ninexnine_unit ninexnine_unit_1518(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26247)
);

ninexnine_unit ninexnine_unit_1519(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27247)
);

assign C2247=c20247+c21247+c22247+c23247+c24247+c25247+c26247+c27247;
assign A2247=(C2247>=0)?1:0;

assign P3247=A2247;

ninexnine_unit ninexnine_unit_1520(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20307)
);

ninexnine_unit ninexnine_unit_1521(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21307)
);

ninexnine_unit ninexnine_unit_1522(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22307)
);

ninexnine_unit ninexnine_unit_1523(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23307)
);

ninexnine_unit ninexnine_unit_1524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24307)
);

ninexnine_unit ninexnine_unit_1525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25307)
);

ninexnine_unit ninexnine_unit_1526(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26307)
);

ninexnine_unit ninexnine_unit_1527(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27307)
);

assign C2307=c20307+c21307+c22307+c23307+c24307+c25307+c26307+c27307;
assign A2307=(C2307>=0)?1:0;

assign P3307=A2307;

ninexnine_unit ninexnine_unit_1528(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20317)
);

ninexnine_unit ninexnine_unit_1529(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21317)
);

ninexnine_unit ninexnine_unit_1530(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22317)
);

ninexnine_unit ninexnine_unit_1531(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23317)
);

ninexnine_unit ninexnine_unit_1532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24317)
);

ninexnine_unit ninexnine_unit_1533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25317)
);

ninexnine_unit ninexnine_unit_1534(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26317)
);

ninexnine_unit ninexnine_unit_1535(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27317)
);

assign C2317=c20317+c21317+c22317+c23317+c24317+c25317+c26317+c27317;
assign A2317=(C2317>=0)?1:0;

assign P3317=A2317;

ninexnine_unit ninexnine_unit_1536(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20327)
);

ninexnine_unit ninexnine_unit_1537(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21327)
);

ninexnine_unit ninexnine_unit_1538(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22327)
);

ninexnine_unit ninexnine_unit_1539(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23327)
);

ninexnine_unit ninexnine_unit_1540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24327)
);

ninexnine_unit ninexnine_unit_1541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25327)
);

ninexnine_unit ninexnine_unit_1542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26327)
);

ninexnine_unit ninexnine_unit_1543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27327)
);

assign C2327=c20327+c21327+c22327+c23327+c24327+c25327+c26327+c27327;
assign A2327=(C2327>=0)?1:0;

assign P3327=A2327;

ninexnine_unit ninexnine_unit_1544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20337)
);

ninexnine_unit ninexnine_unit_1545(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21337)
);

ninexnine_unit ninexnine_unit_1546(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22337)
);

ninexnine_unit ninexnine_unit_1547(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23337)
);

ninexnine_unit ninexnine_unit_1548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24337)
);

ninexnine_unit ninexnine_unit_1549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25337)
);

ninexnine_unit ninexnine_unit_1550(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26337)
);

ninexnine_unit ninexnine_unit_1551(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27337)
);

assign C2337=c20337+c21337+c22337+c23337+c24337+c25337+c26337+c27337;
assign A2337=(C2337>=0)?1:0;

assign P3337=A2337;

ninexnine_unit ninexnine_unit_1552(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20347)
);

ninexnine_unit ninexnine_unit_1553(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21347)
);

ninexnine_unit ninexnine_unit_1554(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22347)
);

ninexnine_unit ninexnine_unit_1555(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23347)
);

ninexnine_unit ninexnine_unit_1556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24347)
);

ninexnine_unit ninexnine_unit_1557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25347)
);

ninexnine_unit ninexnine_unit_1558(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26347)
);

ninexnine_unit ninexnine_unit_1559(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27347)
);

assign C2347=c20347+c21347+c22347+c23347+c24347+c25347+c26347+c27347;
assign A2347=(C2347>=0)?1:0;

assign P3347=A2347;

ninexnine_unit ninexnine_unit_1560(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20407)
);

ninexnine_unit ninexnine_unit_1561(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21407)
);

ninexnine_unit ninexnine_unit_1562(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22407)
);

ninexnine_unit ninexnine_unit_1563(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23407)
);

ninexnine_unit ninexnine_unit_1564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24407)
);

ninexnine_unit ninexnine_unit_1565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25407)
);

ninexnine_unit ninexnine_unit_1566(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26407)
);

ninexnine_unit ninexnine_unit_1567(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27407)
);

assign C2407=c20407+c21407+c22407+c23407+c24407+c25407+c26407+c27407;
assign A2407=(C2407>=0)?1:0;

assign P3407=A2407;

ninexnine_unit ninexnine_unit_1568(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20417)
);

ninexnine_unit ninexnine_unit_1569(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21417)
);

ninexnine_unit ninexnine_unit_1570(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22417)
);

ninexnine_unit ninexnine_unit_1571(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23417)
);

ninexnine_unit ninexnine_unit_1572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24417)
);

ninexnine_unit ninexnine_unit_1573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25417)
);

ninexnine_unit ninexnine_unit_1574(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26417)
);

ninexnine_unit ninexnine_unit_1575(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27417)
);

assign C2417=c20417+c21417+c22417+c23417+c24417+c25417+c26417+c27417;
assign A2417=(C2417>=0)?1:0;

assign P3417=A2417;

ninexnine_unit ninexnine_unit_1576(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20427)
);

ninexnine_unit ninexnine_unit_1577(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21427)
);

ninexnine_unit ninexnine_unit_1578(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22427)
);

ninexnine_unit ninexnine_unit_1579(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23427)
);

ninexnine_unit ninexnine_unit_1580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24427)
);

ninexnine_unit ninexnine_unit_1581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25427)
);

ninexnine_unit ninexnine_unit_1582(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26427)
);

ninexnine_unit ninexnine_unit_1583(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27427)
);

assign C2427=c20427+c21427+c22427+c23427+c24427+c25427+c26427+c27427;
assign A2427=(C2427>=0)?1:0;

assign P3427=A2427;

ninexnine_unit ninexnine_unit_1584(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20437)
);

ninexnine_unit ninexnine_unit_1585(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21437)
);

ninexnine_unit ninexnine_unit_1586(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22437)
);

ninexnine_unit ninexnine_unit_1587(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23437)
);

ninexnine_unit ninexnine_unit_1588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24437)
);

ninexnine_unit ninexnine_unit_1589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25437)
);

ninexnine_unit ninexnine_unit_1590(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26437)
);

ninexnine_unit ninexnine_unit_1591(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27437)
);

assign C2437=c20437+c21437+c22437+c23437+c24437+c25437+c26437+c27437;
assign A2437=(C2437>=0)?1:0;

assign P3437=A2437;

ninexnine_unit ninexnine_unit_1592(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20447)
);

ninexnine_unit ninexnine_unit_1593(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21447)
);

ninexnine_unit ninexnine_unit_1594(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22447)
);

ninexnine_unit ninexnine_unit_1595(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23447)
);

ninexnine_unit ninexnine_unit_1596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24447)
);

ninexnine_unit ninexnine_unit_1597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25447)
);

ninexnine_unit ninexnine_unit_1598(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26447)
);

ninexnine_unit ninexnine_unit_1599(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27447)
);

assign C2447=c20447+c21447+c22447+c23447+c24447+c25447+c26447+c27447;
assign A2447=(C2447>=0)?1:0;

assign P3447=A2447;

ninexnine_unit ninexnine_unit_1600(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20008)
);

ninexnine_unit ninexnine_unit_1601(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21008)
);

ninexnine_unit ninexnine_unit_1602(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22008)
);

ninexnine_unit ninexnine_unit_1603(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23008)
);

ninexnine_unit ninexnine_unit_1604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24008)
);

ninexnine_unit ninexnine_unit_1605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25008)
);

ninexnine_unit ninexnine_unit_1606(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26008)
);

ninexnine_unit ninexnine_unit_1607(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27008)
);

assign C2008=c20008+c21008+c22008+c23008+c24008+c25008+c26008+c27008;
assign A2008=(C2008>=0)?1:0;

assign P3008=A2008;

ninexnine_unit ninexnine_unit_1608(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20018)
);

ninexnine_unit ninexnine_unit_1609(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21018)
);

ninexnine_unit ninexnine_unit_1610(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22018)
);

ninexnine_unit ninexnine_unit_1611(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23018)
);

ninexnine_unit ninexnine_unit_1612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24018)
);

ninexnine_unit ninexnine_unit_1613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25018)
);

ninexnine_unit ninexnine_unit_1614(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26018)
);

ninexnine_unit ninexnine_unit_1615(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27018)
);

assign C2018=c20018+c21018+c22018+c23018+c24018+c25018+c26018+c27018;
assign A2018=(C2018>=0)?1:0;

assign P3018=A2018;

ninexnine_unit ninexnine_unit_1616(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20028)
);

ninexnine_unit ninexnine_unit_1617(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21028)
);

ninexnine_unit ninexnine_unit_1618(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22028)
);

ninexnine_unit ninexnine_unit_1619(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23028)
);

ninexnine_unit ninexnine_unit_1620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24028)
);

ninexnine_unit ninexnine_unit_1621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25028)
);

ninexnine_unit ninexnine_unit_1622(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26028)
);

ninexnine_unit ninexnine_unit_1623(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27028)
);

assign C2028=c20028+c21028+c22028+c23028+c24028+c25028+c26028+c27028;
assign A2028=(C2028>=0)?1:0;

assign P3028=A2028;

ninexnine_unit ninexnine_unit_1624(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20038)
);

ninexnine_unit ninexnine_unit_1625(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21038)
);

ninexnine_unit ninexnine_unit_1626(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22038)
);

ninexnine_unit ninexnine_unit_1627(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23038)
);

ninexnine_unit ninexnine_unit_1628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24038)
);

ninexnine_unit ninexnine_unit_1629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25038)
);

ninexnine_unit ninexnine_unit_1630(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26038)
);

ninexnine_unit ninexnine_unit_1631(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27038)
);

assign C2038=c20038+c21038+c22038+c23038+c24038+c25038+c26038+c27038;
assign A2038=(C2038>=0)?1:0;

assign P3038=A2038;

ninexnine_unit ninexnine_unit_1632(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20048)
);

ninexnine_unit ninexnine_unit_1633(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21048)
);

ninexnine_unit ninexnine_unit_1634(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22048)
);

ninexnine_unit ninexnine_unit_1635(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23048)
);

ninexnine_unit ninexnine_unit_1636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24048)
);

ninexnine_unit ninexnine_unit_1637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25048)
);

ninexnine_unit ninexnine_unit_1638(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26048)
);

ninexnine_unit ninexnine_unit_1639(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27048)
);

assign C2048=c20048+c21048+c22048+c23048+c24048+c25048+c26048+c27048;
assign A2048=(C2048>=0)?1:0;

assign P3048=A2048;

ninexnine_unit ninexnine_unit_1640(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20108)
);

ninexnine_unit ninexnine_unit_1641(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21108)
);

ninexnine_unit ninexnine_unit_1642(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22108)
);

ninexnine_unit ninexnine_unit_1643(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23108)
);

ninexnine_unit ninexnine_unit_1644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24108)
);

ninexnine_unit ninexnine_unit_1645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25108)
);

ninexnine_unit ninexnine_unit_1646(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26108)
);

ninexnine_unit ninexnine_unit_1647(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27108)
);

assign C2108=c20108+c21108+c22108+c23108+c24108+c25108+c26108+c27108;
assign A2108=(C2108>=0)?1:0;

assign P3108=A2108;

ninexnine_unit ninexnine_unit_1648(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20118)
);

ninexnine_unit ninexnine_unit_1649(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21118)
);

ninexnine_unit ninexnine_unit_1650(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22118)
);

ninexnine_unit ninexnine_unit_1651(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23118)
);

ninexnine_unit ninexnine_unit_1652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24118)
);

ninexnine_unit ninexnine_unit_1653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25118)
);

ninexnine_unit ninexnine_unit_1654(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26118)
);

ninexnine_unit ninexnine_unit_1655(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27118)
);

assign C2118=c20118+c21118+c22118+c23118+c24118+c25118+c26118+c27118;
assign A2118=(C2118>=0)?1:0;

assign P3118=A2118;

ninexnine_unit ninexnine_unit_1656(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20128)
);

ninexnine_unit ninexnine_unit_1657(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21128)
);

ninexnine_unit ninexnine_unit_1658(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22128)
);

ninexnine_unit ninexnine_unit_1659(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23128)
);

ninexnine_unit ninexnine_unit_1660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24128)
);

ninexnine_unit ninexnine_unit_1661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25128)
);

ninexnine_unit ninexnine_unit_1662(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26128)
);

ninexnine_unit ninexnine_unit_1663(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27128)
);

assign C2128=c20128+c21128+c22128+c23128+c24128+c25128+c26128+c27128;
assign A2128=(C2128>=0)?1:0;

assign P3128=A2128;

ninexnine_unit ninexnine_unit_1664(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20138)
);

ninexnine_unit ninexnine_unit_1665(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21138)
);

ninexnine_unit ninexnine_unit_1666(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22138)
);

ninexnine_unit ninexnine_unit_1667(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23138)
);

ninexnine_unit ninexnine_unit_1668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24138)
);

ninexnine_unit ninexnine_unit_1669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25138)
);

ninexnine_unit ninexnine_unit_1670(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26138)
);

ninexnine_unit ninexnine_unit_1671(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27138)
);

assign C2138=c20138+c21138+c22138+c23138+c24138+c25138+c26138+c27138;
assign A2138=(C2138>=0)?1:0;

assign P3138=A2138;

ninexnine_unit ninexnine_unit_1672(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20148)
);

ninexnine_unit ninexnine_unit_1673(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21148)
);

ninexnine_unit ninexnine_unit_1674(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22148)
);

ninexnine_unit ninexnine_unit_1675(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23148)
);

ninexnine_unit ninexnine_unit_1676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24148)
);

ninexnine_unit ninexnine_unit_1677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25148)
);

ninexnine_unit ninexnine_unit_1678(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26148)
);

ninexnine_unit ninexnine_unit_1679(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27148)
);

assign C2148=c20148+c21148+c22148+c23148+c24148+c25148+c26148+c27148;
assign A2148=(C2148>=0)?1:0;

assign P3148=A2148;

ninexnine_unit ninexnine_unit_1680(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20208)
);

ninexnine_unit ninexnine_unit_1681(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21208)
);

ninexnine_unit ninexnine_unit_1682(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22208)
);

ninexnine_unit ninexnine_unit_1683(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23208)
);

ninexnine_unit ninexnine_unit_1684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24208)
);

ninexnine_unit ninexnine_unit_1685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25208)
);

ninexnine_unit ninexnine_unit_1686(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26208)
);

ninexnine_unit ninexnine_unit_1687(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27208)
);

assign C2208=c20208+c21208+c22208+c23208+c24208+c25208+c26208+c27208;
assign A2208=(C2208>=0)?1:0;

assign P3208=A2208;

ninexnine_unit ninexnine_unit_1688(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20218)
);

ninexnine_unit ninexnine_unit_1689(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21218)
);

ninexnine_unit ninexnine_unit_1690(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22218)
);

ninexnine_unit ninexnine_unit_1691(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23218)
);

ninexnine_unit ninexnine_unit_1692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24218)
);

ninexnine_unit ninexnine_unit_1693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25218)
);

ninexnine_unit ninexnine_unit_1694(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26218)
);

ninexnine_unit ninexnine_unit_1695(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27218)
);

assign C2218=c20218+c21218+c22218+c23218+c24218+c25218+c26218+c27218;
assign A2218=(C2218>=0)?1:0;

assign P3218=A2218;

ninexnine_unit ninexnine_unit_1696(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20228)
);

ninexnine_unit ninexnine_unit_1697(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21228)
);

ninexnine_unit ninexnine_unit_1698(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22228)
);

ninexnine_unit ninexnine_unit_1699(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23228)
);

ninexnine_unit ninexnine_unit_1700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24228)
);

ninexnine_unit ninexnine_unit_1701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25228)
);

ninexnine_unit ninexnine_unit_1702(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26228)
);

ninexnine_unit ninexnine_unit_1703(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27228)
);

assign C2228=c20228+c21228+c22228+c23228+c24228+c25228+c26228+c27228;
assign A2228=(C2228>=0)?1:0;

assign P3228=A2228;

ninexnine_unit ninexnine_unit_1704(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20238)
);

ninexnine_unit ninexnine_unit_1705(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21238)
);

ninexnine_unit ninexnine_unit_1706(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22238)
);

ninexnine_unit ninexnine_unit_1707(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23238)
);

ninexnine_unit ninexnine_unit_1708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24238)
);

ninexnine_unit ninexnine_unit_1709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25238)
);

ninexnine_unit ninexnine_unit_1710(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26238)
);

ninexnine_unit ninexnine_unit_1711(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27238)
);

assign C2238=c20238+c21238+c22238+c23238+c24238+c25238+c26238+c27238;
assign A2238=(C2238>=0)?1:0;

assign P3238=A2238;

ninexnine_unit ninexnine_unit_1712(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20248)
);

ninexnine_unit ninexnine_unit_1713(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21248)
);

ninexnine_unit ninexnine_unit_1714(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22248)
);

ninexnine_unit ninexnine_unit_1715(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23248)
);

ninexnine_unit ninexnine_unit_1716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24248)
);

ninexnine_unit ninexnine_unit_1717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25248)
);

ninexnine_unit ninexnine_unit_1718(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26248)
);

ninexnine_unit ninexnine_unit_1719(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27248)
);

assign C2248=c20248+c21248+c22248+c23248+c24248+c25248+c26248+c27248;
assign A2248=(C2248>=0)?1:0;

assign P3248=A2248;

ninexnine_unit ninexnine_unit_1720(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20308)
);

ninexnine_unit ninexnine_unit_1721(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21308)
);

ninexnine_unit ninexnine_unit_1722(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22308)
);

ninexnine_unit ninexnine_unit_1723(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23308)
);

ninexnine_unit ninexnine_unit_1724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24308)
);

ninexnine_unit ninexnine_unit_1725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25308)
);

ninexnine_unit ninexnine_unit_1726(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26308)
);

ninexnine_unit ninexnine_unit_1727(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27308)
);

assign C2308=c20308+c21308+c22308+c23308+c24308+c25308+c26308+c27308;
assign A2308=(C2308>=0)?1:0;

assign P3308=A2308;

ninexnine_unit ninexnine_unit_1728(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20318)
);

ninexnine_unit ninexnine_unit_1729(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21318)
);

ninexnine_unit ninexnine_unit_1730(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22318)
);

ninexnine_unit ninexnine_unit_1731(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23318)
);

ninexnine_unit ninexnine_unit_1732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24318)
);

ninexnine_unit ninexnine_unit_1733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25318)
);

ninexnine_unit ninexnine_unit_1734(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26318)
);

ninexnine_unit ninexnine_unit_1735(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27318)
);

assign C2318=c20318+c21318+c22318+c23318+c24318+c25318+c26318+c27318;
assign A2318=(C2318>=0)?1:0;

assign P3318=A2318;

ninexnine_unit ninexnine_unit_1736(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20328)
);

ninexnine_unit ninexnine_unit_1737(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21328)
);

ninexnine_unit ninexnine_unit_1738(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22328)
);

ninexnine_unit ninexnine_unit_1739(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23328)
);

ninexnine_unit ninexnine_unit_1740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24328)
);

ninexnine_unit ninexnine_unit_1741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25328)
);

ninexnine_unit ninexnine_unit_1742(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26328)
);

ninexnine_unit ninexnine_unit_1743(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27328)
);

assign C2328=c20328+c21328+c22328+c23328+c24328+c25328+c26328+c27328;
assign A2328=(C2328>=0)?1:0;

assign P3328=A2328;

ninexnine_unit ninexnine_unit_1744(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20338)
);

ninexnine_unit ninexnine_unit_1745(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21338)
);

ninexnine_unit ninexnine_unit_1746(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22338)
);

ninexnine_unit ninexnine_unit_1747(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23338)
);

ninexnine_unit ninexnine_unit_1748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24338)
);

ninexnine_unit ninexnine_unit_1749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25338)
);

ninexnine_unit ninexnine_unit_1750(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26338)
);

ninexnine_unit ninexnine_unit_1751(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27338)
);

assign C2338=c20338+c21338+c22338+c23338+c24338+c25338+c26338+c27338;
assign A2338=(C2338>=0)?1:0;

assign P3338=A2338;

ninexnine_unit ninexnine_unit_1752(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20348)
);

ninexnine_unit ninexnine_unit_1753(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21348)
);

ninexnine_unit ninexnine_unit_1754(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22348)
);

ninexnine_unit ninexnine_unit_1755(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23348)
);

ninexnine_unit ninexnine_unit_1756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24348)
);

ninexnine_unit ninexnine_unit_1757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25348)
);

ninexnine_unit ninexnine_unit_1758(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26348)
);

ninexnine_unit ninexnine_unit_1759(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27348)
);

assign C2348=c20348+c21348+c22348+c23348+c24348+c25348+c26348+c27348;
assign A2348=(C2348>=0)?1:0;

assign P3348=A2348;

ninexnine_unit ninexnine_unit_1760(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20408)
);

ninexnine_unit ninexnine_unit_1761(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21408)
);

ninexnine_unit ninexnine_unit_1762(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22408)
);

ninexnine_unit ninexnine_unit_1763(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23408)
);

ninexnine_unit ninexnine_unit_1764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24408)
);

ninexnine_unit ninexnine_unit_1765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25408)
);

ninexnine_unit ninexnine_unit_1766(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26408)
);

ninexnine_unit ninexnine_unit_1767(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27408)
);

assign C2408=c20408+c21408+c22408+c23408+c24408+c25408+c26408+c27408;
assign A2408=(C2408>=0)?1:0;

assign P3408=A2408;

ninexnine_unit ninexnine_unit_1768(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20418)
);

ninexnine_unit ninexnine_unit_1769(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21418)
);

ninexnine_unit ninexnine_unit_1770(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22418)
);

ninexnine_unit ninexnine_unit_1771(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23418)
);

ninexnine_unit ninexnine_unit_1772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24418)
);

ninexnine_unit ninexnine_unit_1773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25418)
);

ninexnine_unit ninexnine_unit_1774(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26418)
);

ninexnine_unit ninexnine_unit_1775(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27418)
);

assign C2418=c20418+c21418+c22418+c23418+c24418+c25418+c26418+c27418;
assign A2418=(C2418>=0)?1:0;

assign P3418=A2418;

ninexnine_unit ninexnine_unit_1776(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20428)
);

ninexnine_unit ninexnine_unit_1777(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21428)
);

ninexnine_unit ninexnine_unit_1778(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22428)
);

ninexnine_unit ninexnine_unit_1779(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23428)
);

ninexnine_unit ninexnine_unit_1780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24428)
);

ninexnine_unit ninexnine_unit_1781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25428)
);

ninexnine_unit ninexnine_unit_1782(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26428)
);

ninexnine_unit ninexnine_unit_1783(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27428)
);

assign C2428=c20428+c21428+c22428+c23428+c24428+c25428+c26428+c27428;
assign A2428=(C2428>=0)?1:0;

assign P3428=A2428;

ninexnine_unit ninexnine_unit_1784(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20438)
);

ninexnine_unit ninexnine_unit_1785(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21438)
);

ninexnine_unit ninexnine_unit_1786(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22438)
);

ninexnine_unit ninexnine_unit_1787(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23438)
);

ninexnine_unit ninexnine_unit_1788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24438)
);

ninexnine_unit ninexnine_unit_1789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25438)
);

ninexnine_unit ninexnine_unit_1790(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26438)
);

ninexnine_unit ninexnine_unit_1791(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27438)
);

assign C2438=c20438+c21438+c22438+c23438+c24438+c25438+c26438+c27438;
assign A2438=(C2438>=0)?1:0;

assign P3438=A2438;

ninexnine_unit ninexnine_unit_1792(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20448)
);

ninexnine_unit ninexnine_unit_1793(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21448)
);

ninexnine_unit ninexnine_unit_1794(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22448)
);

ninexnine_unit ninexnine_unit_1795(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23448)
);

ninexnine_unit ninexnine_unit_1796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24448)
);

ninexnine_unit ninexnine_unit_1797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25448)
);

ninexnine_unit ninexnine_unit_1798(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26448)
);

ninexnine_unit ninexnine_unit_1799(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27448)
);

assign C2448=c20448+c21448+c22448+c23448+c24448+c25448+c26448+c27448;
assign A2448=(C2448>=0)?1:0;

assign P3448=A2448;

ninexnine_unit ninexnine_unit_1800(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20009)
);

ninexnine_unit ninexnine_unit_1801(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21009)
);

ninexnine_unit ninexnine_unit_1802(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22009)
);

ninexnine_unit ninexnine_unit_1803(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23009)
);

ninexnine_unit ninexnine_unit_1804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24009)
);

ninexnine_unit ninexnine_unit_1805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25009)
);

ninexnine_unit ninexnine_unit_1806(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26009)
);

ninexnine_unit ninexnine_unit_1807(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27009)
);

assign C2009=c20009+c21009+c22009+c23009+c24009+c25009+c26009+c27009;
assign A2009=(C2009>=0)?1:0;

assign P3009=A2009;

ninexnine_unit ninexnine_unit_1808(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20019)
);

ninexnine_unit ninexnine_unit_1809(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21019)
);

ninexnine_unit ninexnine_unit_1810(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22019)
);

ninexnine_unit ninexnine_unit_1811(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23019)
);

ninexnine_unit ninexnine_unit_1812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24019)
);

ninexnine_unit ninexnine_unit_1813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25019)
);

ninexnine_unit ninexnine_unit_1814(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26019)
);

ninexnine_unit ninexnine_unit_1815(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27019)
);

assign C2019=c20019+c21019+c22019+c23019+c24019+c25019+c26019+c27019;
assign A2019=(C2019>=0)?1:0;

assign P3019=A2019;

ninexnine_unit ninexnine_unit_1816(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20029)
);

ninexnine_unit ninexnine_unit_1817(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21029)
);

ninexnine_unit ninexnine_unit_1818(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22029)
);

ninexnine_unit ninexnine_unit_1819(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23029)
);

ninexnine_unit ninexnine_unit_1820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24029)
);

ninexnine_unit ninexnine_unit_1821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25029)
);

ninexnine_unit ninexnine_unit_1822(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26029)
);

ninexnine_unit ninexnine_unit_1823(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27029)
);

assign C2029=c20029+c21029+c22029+c23029+c24029+c25029+c26029+c27029;
assign A2029=(C2029>=0)?1:0;

assign P3029=A2029;

ninexnine_unit ninexnine_unit_1824(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20039)
);

ninexnine_unit ninexnine_unit_1825(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21039)
);

ninexnine_unit ninexnine_unit_1826(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22039)
);

ninexnine_unit ninexnine_unit_1827(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23039)
);

ninexnine_unit ninexnine_unit_1828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24039)
);

ninexnine_unit ninexnine_unit_1829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25039)
);

ninexnine_unit ninexnine_unit_1830(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26039)
);

ninexnine_unit ninexnine_unit_1831(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27039)
);

assign C2039=c20039+c21039+c22039+c23039+c24039+c25039+c26039+c27039;
assign A2039=(C2039>=0)?1:0;

assign P3039=A2039;

ninexnine_unit ninexnine_unit_1832(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20049)
);

ninexnine_unit ninexnine_unit_1833(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21049)
);

ninexnine_unit ninexnine_unit_1834(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22049)
);

ninexnine_unit ninexnine_unit_1835(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23049)
);

ninexnine_unit ninexnine_unit_1836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24049)
);

ninexnine_unit ninexnine_unit_1837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25049)
);

ninexnine_unit ninexnine_unit_1838(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26049)
);

ninexnine_unit ninexnine_unit_1839(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27049)
);

assign C2049=c20049+c21049+c22049+c23049+c24049+c25049+c26049+c27049;
assign A2049=(C2049>=0)?1:0;

assign P3049=A2049;

ninexnine_unit ninexnine_unit_1840(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20109)
);

ninexnine_unit ninexnine_unit_1841(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21109)
);

ninexnine_unit ninexnine_unit_1842(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22109)
);

ninexnine_unit ninexnine_unit_1843(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23109)
);

ninexnine_unit ninexnine_unit_1844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24109)
);

ninexnine_unit ninexnine_unit_1845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25109)
);

ninexnine_unit ninexnine_unit_1846(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26109)
);

ninexnine_unit ninexnine_unit_1847(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27109)
);

assign C2109=c20109+c21109+c22109+c23109+c24109+c25109+c26109+c27109;
assign A2109=(C2109>=0)?1:0;

assign P3109=A2109;

ninexnine_unit ninexnine_unit_1848(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20119)
);

ninexnine_unit ninexnine_unit_1849(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21119)
);

ninexnine_unit ninexnine_unit_1850(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22119)
);

ninexnine_unit ninexnine_unit_1851(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23119)
);

ninexnine_unit ninexnine_unit_1852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24119)
);

ninexnine_unit ninexnine_unit_1853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25119)
);

ninexnine_unit ninexnine_unit_1854(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26119)
);

ninexnine_unit ninexnine_unit_1855(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27119)
);

assign C2119=c20119+c21119+c22119+c23119+c24119+c25119+c26119+c27119;
assign A2119=(C2119>=0)?1:0;

assign P3119=A2119;

ninexnine_unit ninexnine_unit_1856(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20129)
);

ninexnine_unit ninexnine_unit_1857(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21129)
);

ninexnine_unit ninexnine_unit_1858(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22129)
);

ninexnine_unit ninexnine_unit_1859(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23129)
);

ninexnine_unit ninexnine_unit_1860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24129)
);

ninexnine_unit ninexnine_unit_1861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25129)
);

ninexnine_unit ninexnine_unit_1862(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26129)
);

ninexnine_unit ninexnine_unit_1863(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27129)
);

assign C2129=c20129+c21129+c22129+c23129+c24129+c25129+c26129+c27129;
assign A2129=(C2129>=0)?1:0;

assign P3129=A2129;

ninexnine_unit ninexnine_unit_1864(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20139)
);

ninexnine_unit ninexnine_unit_1865(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21139)
);

ninexnine_unit ninexnine_unit_1866(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22139)
);

ninexnine_unit ninexnine_unit_1867(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23139)
);

ninexnine_unit ninexnine_unit_1868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24139)
);

ninexnine_unit ninexnine_unit_1869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25139)
);

ninexnine_unit ninexnine_unit_1870(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26139)
);

ninexnine_unit ninexnine_unit_1871(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27139)
);

assign C2139=c20139+c21139+c22139+c23139+c24139+c25139+c26139+c27139;
assign A2139=(C2139>=0)?1:0;

assign P3139=A2139;

ninexnine_unit ninexnine_unit_1872(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20149)
);

ninexnine_unit ninexnine_unit_1873(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21149)
);

ninexnine_unit ninexnine_unit_1874(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22149)
);

ninexnine_unit ninexnine_unit_1875(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23149)
);

ninexnine_unit ninexnine_unit_1876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24149)
);

ninexnine_unit ninexnine_unit_1877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25149)
);

ninexnine_unit ninexnine_unit_1878(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26149)
);

ninexnine_unit ninexnine_unit_1879(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27149)
);

assign C2149=c20149+c21149+c22149+c23149+c24149+c25149+c26149+c27149;
assign A2149=(C2149>=0)?1:0;

assign P3149=A2149;

ninexnine_unit ninexnine_unit_1880(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20209)
);

ninexnine_unit ninexnine_unit_1881(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21209)
);

ninexnine_unit ninexnine_unit_1882(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22209)
);

ninexnine_unit ninexnine_unit_1883(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23209)
);

ninexnine_unit ninexnine_unit_1884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24209)
);

ninexnine_unit ninexnine_unit_1885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25209)
);

ninexnine_unit ninexnine_unit_1886(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26209)
);

ninexnine_unit ninexnine_unit_1887(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27209)
);

assign C2209=c20209+c21209+c22209+c23209+c24209+c25209+c26209+c27209;
assign A2209=(C2209>=0)?1:0;

assign P3209=A2209;

ninexnine_unit ninexnine_unit_1888(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20219)
);

ninexnine_unit ninexnine_unit_1889(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21219)
);

ninexnine_unit ninexnine_unit_1890(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22219)
);

ninexnine_unit ninexnine_unit_1891(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23219)
);

ninexnine_unit ninexnine_unit_1892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24219)
);

ninexnine_unit ninexnine_unit_1893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25219)
);

ninexnine_unit ninexnine_unit_1894(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26219)
);

ninexnine_unit ninexnine_unit_1895(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27219)
);

assign C2219=c20219+c21219+c22219+c23219+c24219+c25219+c26219+c27219;
assign A2219=(C2219>=0)?1:0;

assign P3219=A2219;

ninexnine_unit ninexnine_unit_1896(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20229)
);

ninexnine_unit ninexnine_unit_1897(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21229)
);

ninexnine_unit ninexnine_unit_1898(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22229)
);

ninexnine_unit ninexnine_unit_1899(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23229)
);

ninexnine_unit ninexnine_unit_1900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24229)
);

ninexnine_unit ninexnine_unit_1901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25229)
);

ninexnine_unit ninexnine_unit_1902(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26229)
);

ninexnine_unit ninexnine_unit_1903(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27229)
);

assign C2229=c20229+c21229+c22229+c23229+c24229+c25229+c26229+c27229;
assign A2229=(C2229>=0)?1:0;

assign P3229=A2229;

ninexnine_unit ninexnine_unit_1904(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20239)
);

ninexnine_unit ninexnine_unit_1905(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21239)
);

ninexnine_unit ninexnine_unit_1906(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22239)
);

ninexnine_unit ninexnine_unit_1907(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23239)
);

ninexnine_unit ninexnine_unit_1908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24239)
);

ninexnine_unit ninexnine_unit_1909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25239)
);

ninexnine_unit ninexnine_unit_1910(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26239)
);

ninexnine_unit ninexnine_unit_1911(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27239)
);

assign C2239=c20239+c21239+c22239+c23239+c24239+c25239+c26239+c27239;
assign A2239=(C2239>=0)?1:0;

assign P3239=A2239;

ninexnine_unit ninexnine_unit_1912(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20249)
);

ninexnine_unit ninexnine_unit_1913(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21249)
);

ninexnine_unit ninexnine_unit_1914(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22249)
);

ninexnine_unit ninexnine_unit_1915(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23249)
);

ninexnine_unit ninexnine_unit_1916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24249)
);

ninexnine_unit ninexnine_unit_1917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25249)
);

ninexnine_unit ninexnine_unit_1918(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26249)
);

ninexnine_unit ninexnine_unit_1919(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27249)
);

assign C2249=c20249+c21249+c22249+c23249+c24249+c25249+c26249+c27249;
assign A2249=(C2249>=0)?1:0;

assign P3249=A2249;

ninexnine_unit ninexnine_unit_1920(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20309)
);

ninexnine_unit ninexnine_unit_1921(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21309)
);

ninexnine_unit ninexnine_unit_1922(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22309)
);

ninexnine_unit ninexnine_unit_1923(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23309)
);

ninexnine_unit ninexnine_unit_1924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24309)
);

ninexnine_unit ninexnine_unit_1925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25309)
);

ninexnine_unit ninexnine_unit_1926(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26309)
);

ninexnine_unit ninexnine_unit_1927(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27309)
);

assign C2309=c20309+c21309+c22309+c23309+c24309+c25309+c26309+c27309;
assign A2309=(C2309>=0)?1:0;

assign P3309=A2309;

ninexnine_unit ninexnine_unit_1928(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20319)
);

ninexnine_unit ninexnine_unit_1929(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21319)
);

ninexnine_unit ninexnine_unit_1930(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22319)
);

ninexnine_unit ninexnine_unit_1931(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23319)
);

ninexnine_unit ninexnine_unit_1932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24319)
);

ninexnine_unit ninexnine_unit_1933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25319)
);

ninexnine_unit ninexnine_unit_1934(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26319)
);

ninexnine_unit ninexnine_unit_1935(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27319)
);

assign C2319=c20319+c21319+c22319+c23319+c24319+c25319+c26319+c27319;
assign A2319=(C2319>=0)?1:0;

assign P3319=A2319;

ninexnine_unit ninexnine_unit_1936(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20329)
);

ninexnine_unit ninexnine_unit_1937(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21329)
);

ninexnine_unit ninexnine_unit_1938(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22329)
);

ninexnine_unit ninexnine_unit_1939(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23329)
);

ninexnine_unit ninexnine_unit_1940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24329)
);

ninexnine_unit ninexnine_unit_1941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25329)
);

ninexnine_unit ninexnine_unit_1942(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26329)
);

ninexnine_unit ninexnine_unit_1943(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27329)
);

assign C2329=c20329+c21329+c22329+c23329+c24329+c25329+c26329+c27329;
assign A2329=(C2329>=0)?1:0;

assign P3329=A2329;

ninexnine_unit ninexnine_unit_1944(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20339)
);

ninexnine_unit ninexnine_unit_1945(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21339)
);

ninexnine_unit ninexnine_unit_1946(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22339)
);

ninexnine_unit ninexnine_unit_1947(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23339)
);

ninexnine_unit ninexnine_unit_1948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24339)
);

ninexnine_unit ninexnine_unit_1949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25339)
);

ninexnine_unit ninexnine_unit_1950(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26339)
);

ninexnine_unit ninexnine_unit_1951(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27339)
);

assign C2339=c20339+c21339+c22339+c23339+c24339+c25339+c26339+c27339;
assign A2339=(C2339>=0)?1:0;

assign P3339=A2339;

ninexnine_unit ninexnine_unit_1952(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20349)
);

ninexnine_unit ninexnine_unit_1953(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21349)
);

ninexnine_unit ninexnine_unit_1954(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22349)
);

ninexnine_unit ninexnine_unit_1955(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23349)
);

ninexnine_unit ninexnine_unit_1956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24349)
);

ninexnine_unit ninexnine_unit_1957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25349)
);

ninexnine_unit ninexnine_unit_1958(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26349)
);

ninexnine_unit ninexnine_unit_1959(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27349)
);

assign C2349=c20349+c21349+c22349+c23349+c24349+c25349+c26349+c27349;
assign A2349=(C2349>=0)?1:0;

assign P3349=A2349;

ninexnine_unit ninexnine_unit_1960(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20409)
);

ninexnine_unit ninexnine_unit_1961(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21409)
);

ninexnine_unit ninexnine_unit_1962(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22409)
);

ninexnine_unit ninexnine_unit_1963(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23409)
);

ninexnine_unit ninexnine_unit_1964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24409)
);

ninexnine_unit ninexnine_unit_1965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25409)
);

ninexnine_unit ninexnine_unit_1966(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26409)
);

ninexnine_unit ninexnine_unit_1967(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27409)
);

assign C2409=c20409+c21409+c22409+c23409+c24409+c25409+c26409+c27409;
assign A2409=(C2409>=0)?1:0;

assign P3409=A2409;

ninexnine_unit ninexnine_unit_1968(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20419)
);

ninexnine_unit ninexnine_unit_1969(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21419)
);

ninexnine_unit ninexnine_unit_1970(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22419)
);

ninexnine_unit ninexnine_unit_1971(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23419)
);

ninexnine_unit ninexnine_unit_1972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24419)
);

ninexnine_unit ninexnine_unit_1973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25419)
);

ninexnine_unit ninexnine_unit_1974(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26419)
);

ninexnine_unit ninexnine_unit_1975(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27419)
);

assign C2419=c20419+c21419+c22419+c23419+c24419+c25419+c26419+c27419;
assign A2419=(C2419>=0)?1:0;

assign P3419=A2419;

ninexnine_unit ninexnine_unit_1976(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20429)
);

ninexnine_unit ninexnine_unit_1977(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21429)
);

ninexnine_unit ninexnine_unit_1978(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22429)
);

ninexnine_unit ninexnine_unit_1979(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23429)
);

ninexnine_unit ninexnine_unit_1980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24429)
);

ninexnine_unit ninexnine_unit_1981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25429)
);

ninexnine_unit ninexnine_unit_1982(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26429)
);

ninexnine_unit ninexnine_unit_1983(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27429)
);

assign C2429=c20429+c21429+c22429+c23429+c24429+c25429+c26429+c27429;
assign A2429=(C2429>=0)?1:0;

assign P3429=A2429;

ninexnine_unit ninexnine_unit_1984(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20439)
);

ninexnine_unit ninexnine_unit_1985(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21439)
);

ninexnine_unit ninexnine_unit_1986(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22439)
);

ninexnine_unit ninexnine_unit_1987(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23439)
);

ninexnine_unit ninexnine_unit_1988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24439)
);

ninexnine_unit ninexnine_unit_1989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25439)
);

ninexnine_unit ninexnine_unit_1990(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26439)
);

ninexnine_unit ninexnine_unit_1991(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27439)
);

assign C2439=c20439+c21439+c22439+c23439+c24439+c25439+c26439+c27439;
assign A2439=(C2439>=0)?1:0;

assign P3439=A2439;

ninexnine_unit ninexnine_unit_1992(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20449)
);

ninexnine_unit ninexnine_unit_1993(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21449)
);

ninexnine_unit ninexnine_unit_1994(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22449)
);

ninexnine_unit ninexnine_unit_1995(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23449)
);

ninexnine_unit ninexnine_unit_1996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24449)
);

ninexnine_unit ninexnine_unit_1997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25449)
);

ninexnine_unit ninexnine_unit_1998(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26449)
);

ninexnine_unit ninexnine_unit_1999(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27449)
);

assign C2449=c20449+c21449+c22449+c23449+c24449+c25449+c26449+c27449;
assign A2449=(C2449>=0)?1:0;

assign P3449=A2449;

ninexnine_unit ninexnine_unit_2000(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2000A)
);

ninexnine_unit ninexnine_unit_2001(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2100A)
);

ninexnine_unit ninexnine_unit_2002(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2200A)
);

ninexnine_unit ninexnine_unit_2003(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2300A)
);

ninexnine_unit ninexnine_unit_2004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2400A)
);

ninexnine_unit ninexnine_unit_2005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2500A)
);

ninexnine_unit ninexnine_unit_2006(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2600A)
);

ninexnine_unit ninexnine_unit_2007(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2700A)
);

assign C200A=c2000A+c2100A+c2200A+c2300A+c2400A+c2500A+c2600A+c2700A;
assign A200A=(C200A>=0)?1:0;

assign P300A=A200A;

ninexnine_unit ninexnine_unit_2008(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2001A)
);

ninexnine_unit ninexnine_unit_2009(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2101A)
);

ninexnine_unit ninexnine_unit_2010(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2201A)
);

ninexnine_unit ninexnine_unit_2011(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2301A)
);

ninexnine_unit ninexnine_unit_2012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2401A)
);

ninexnine_unit ninexnine_unit_2013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2501A)
);

ninexnine_unit ninexnine_unit_2014(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2601A)
);

ninexnine_unit ninexnine_unit_2015(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2701A)
);

assign C201A=c2001A+c2101A+c2201A+c2301A+c2401A+c2501A+c2601A+c2701A;
assign A201A=(C201A>=0)?1:0;

assign P301A=A201A;

ninexnine_unit ninexnine_unit_2016(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2002A)
);

ninexnine_unit ninexnine_unit_2017(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2102A)
);

ninexnine_unit ninexnine_unit_2018(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2202A)
);

ninexnine_unit ninexnine_unit_2019(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2302A)
);

ninexnine_unit ninexnine_unit_2020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2402A)
);

ninexnine_unit ninexnine_unit_2021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2502A)
);

ninexnine_unit ninexnine_unit_2022(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2602A)
);

ninexnine_unit ninexnine_unit_2023(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2702A)
);

assign C202A=c2002A+c2102A+c2202A+c2302A+c2402A+c2502A+c2602A+c2702A;
assign A202A=(C202A>=0)?1:0;

assign P302A=A202A;

ninexnine_unit ninexnine_unit_2024(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2003A)
);

ninexnine_unit ninexnine_unit_2025(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2103A)
);

ninexnine_unit ninexnine_unit_2026(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2203A)
);

ninexnine_unit ninexnine_unit_2027(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2303A)
);

ninexnine_unit ninexnine_unit_2028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2403A)
);

ninexnine_unit ninexnine_unit_2029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2503A)
);

ninexnine_unit ninexnine_unit_2030(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2603A)
);

ninexnine_unit ninexnine_unit_2031(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2703A)
);

assign C203A=c2003A+c2103A+c2203A+c2303A+c2403A+c2503A+c2603A+c2703A;
assign A203A=(C203A>=0)?1:0;

assign P303A=A203A;

ninexnine_unit ninexnine_unit_2032(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2004A)
);

ninexnine_unit ninexnine_unit_2033(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2104A)
);

ninexnine_unit ninexnine_unit_2034(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2204A)
);

ninexnine_unit ninexnine_unit_2035(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2304A)
);

ninexnine_unit ninexnine_unit_2036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2404A)
);

ninexnine_unit ninexnine_unit_2037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2504A)
);

ninexnine_unit ninexnine_unit_2038(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2604A)
);

ninexnine_unit ninexnine_unit_2039(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2704A)
);

assign C204A=c2004A+c2104A+c2204A+c2304A+c2404A+c2504A+c2604A+c2704A;
assign A204A=(C204A>=0)?1:0;

assign P304A=A204A;

ninexnine_unit ninexnine_unit_2040(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2010A)
);

ninexnine_unit ninexnine_unit_2041(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2110A)
);

ninexnine_unit ninexnine_unit_2042(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2210A)
);

ninexnine_unit ninexnine_unit_2043(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2310A)
);

ninexnine_unit ninexnine_unit_2044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2410A)
);

ninexnine_unit ninexnine_unit_2045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2510A)
);

ninexnine_unit ninexnine_unit_2046(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2610A)
);

ninexnine_unit ninexnine_unit_2047(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2710A)
);

assign C210A=c2010A+c2110A+c2210A+c2310A+c2410A+c2510A+c2610A+c2710A;
assign A210A=(C210A>=0)?1:0;

assign P310A=A210A;

ninexnine_unit ninexnine_unit_2048(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2011A)
);

ninexnine_unit ninexnine_unit_2049(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2111A)
);

ninexnine_unit ninexnine_unit_2050(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2211A)
);

ninexnine_unit ninexnine_unit_2051(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2311A)
);

ninexnine_unit ninexnine_unit_2052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2411A)
);

ninexnine_unit ninexnine_unit_2053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2511A)
);

ninexnine_unit ninexnine_unit_2054(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2611A)
);

ninexnine_unit ninexnine_unit_2055(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2711A)
);

assign C211A=c2011A+c2111A+c2211A+c2311A+c2411A+c2511A+c2611A+c2711A;
assign A211A=(C211A>=0)?1:0;

assign P311A=A211A;

ninexnine_unit ninexnine_unit_2056(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2012A)
);

ninexnine_unit ninexnine_unit_2057(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2112A)
);

ninexnine_unit ninexnine_unit_2058(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2212A)
);

ninexnine_unit ninexnine_unit_2059(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2312A)
);

ninexnine_unit ninexnine_unit_2060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2412A)
);

ninexnine_unit ninexnine_unit_2061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2512A)
);

ninexnine_unit ninexnine_unit_2062(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2612A)
);

ninexnine_unit ninexnine_unit_2063(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2712A)
);

assign C212A=c2012A+c2112A+c2212A+c2312A+c2412A+c2512A+c2612A+c2712A;
assign A212A=(C212A>=0)?1:0;

assign P312A=A212A;

ninexnine_unit ninexnine_unit_2064(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2013A)
);

ninexnine_unit ninexnine_unit_2065(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2113A)
);

ninexnine_unit ninexnine_unit_2066(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2213A)
);

ninexnine_unit ninexnine_unit_2067(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2313A)
);

ninexnine_unit ninexnine_unit_2068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2413A)
);

ninexnine_unit ninexnine_unit_2069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2513A)
);

ninexnine_unit ninexnine_unit_2070(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2613A)
);

ninexnine_unit ninexnine_unit_2071(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2713A)
);

assign C213A=c2013A+c2113A+c2213A+c2313A+c2413A+c2513A+c2613A+c2713A;
assign A213A=(C213A>=0)?1:0;

assign P313A=A213A;

ninexnine_unit ninexnine_unit_2072(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2014A)
);

ninexnine_unit ninexnine_unit_2073(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2114A)
);

ninexnine_unit ninexnine_unit_2074(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2214A)
);

ninexnine_unit ninexnine_unit_2075(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2314A)
);

ninexnine_unit ninexnine_unit_2076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2414A)
);

ninexnine_unit ninexnine_unit_2077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2514A)
);

ninexnine_unit ninexnine_unit_2078(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2614A)
);

ninexnine_unit ninexnine_unit_2079(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2714A)
);

assign C214A=c2014A+c2114A+c2214A+c2314A+c2414A+c2514A+c2614A+c2714A;
assign A214A=(C214A>=0)?1:0;

assign P314A=A214A;

ninexnine_unit ninexnine_unit_2080(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2020A)
);

ninexnine_unit ninexnine_unit_2081(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2120A)
);

ninexnine_unit ninexnine_unit_2082(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2220A)
);

ninexnine_unit ninexnine_unit_2083(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2320A)
);

ninexnine_unit ninexnine_unit_2084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2420A)
);

ninexnine_unit ninexnine_unit_2085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2520A)
);

ninexnine_unit ninexnine_unit_2086(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2620A)
);

ninexnine_unit ninexnine_unit_2087(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2720A)
);

assign C220A=c2020A+c2120A+c2220A+c2320A+c2420A+c2520A+c2620A+c2720A;
assign A220A=(C220A>=0)?1:0;

assign P320A=A220A;

ninexnine_unit ninexnine_unit_2088(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2021A)
);

ninexnine_unit ninexnine_unit_2089(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2121A)
);

ninexnine_unit ninexnine_unit_2090(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2221A)
);

ninexnine_unit ninexnine_unit_2091(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2321A)
);

ninexnine_unit ninexnine_unit_2092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2421A)
);

ninexnine_unit ninexnine_unit_2093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2521A)
);

ninexnine_unit ninexnine_unit_2094(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2621A)
);

ninexnine_unit ninexnine_unit_2095(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2721A)
);

assign C221A=c2021A+c2121A+c2221A+c2321A+c2421A+c2521A+c2621A+c2721A;
assign A221A=(C221A>=0)?1:0;

assign P321A=A221A;

ninexnine_unit ninexnine_unit_2096(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2022A)
);

ninexnine_unit ninexnine_unit_2097(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2122A)
);

ninexnine_unit ninexnine_unit_2098(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2222A)
);

ninexnine_unit ninexnine_unit_2099(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2322A)
);

ninexnine_unit ninexnine_unit_2100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2422A)
);

ninexnine_unit ninexnine_unit_2101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2522A)
);

ninexnine_unit ninexnine_unit_2102(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2622A)
);

ninexnine_unit ninexnine_unit_2103(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2722A)
);

assign C222A=c2022A+c2122A+c2222A+c2322A+c2422A+c2522A+c2622A+c2722A;
assign A222A=(C222A>=0)?1:0;

assign P322A=A222A;

ninexnine_unit ninexnine_unit_2104(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2023A)
);

ninexnine_unit ninexnine_unit_2105(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2123A)
);

ninexnine_unit ninexnine_unit_2106(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2223A)
);

ninexnine_unit ninexnine_unit_2107(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2323A)
);

ninexnine_unit ninexnine_unit_2108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2423A)
);

ninexnine_unit ninexnine_unit_2109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2523A)
);

ninexnine_unit ninexnine_unit_2110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2623A)
);

ninexnine_unit ninexnine_unit_2111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2723A)
);

assign C223A=c2023A+c2123A+c2223A+c2323A+c2423A+c2523A+c2623A+c2723A;
assign A223A=(C223A>=0)?1:0;

assign P323A=A223A;

ninexnine_unit ninexnine_unit_2112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2024A)
);

ninexnine_unit ninexnine_unit_2113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2124A)
);

ninexnine_unit ninexnine_unit_2114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2224A)
);

ninexnine_unit ninexnine_unit_2115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2324A)
);

ninexnine_unit ninexnine_unit_2116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2424A)
);

ninexnine_unit ninexnine_unit_2117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2524A)
);

ninexnine_unit ninexnine_unit_2118(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2624A)
);

ninexnine_unit ninexnine_unit_2119(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2724A)
);

assign C224A=c2024A+c2124A+c2224A+c2324A+c2424A+c2524A+c2624A+c2724A;
assign A224A=(C224A>=0)?1:0;

assign P324A=A224A;

ninexnine_unit ninexnine_unit_2120(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2030A)
);

ninexnine_unit ninexnine_unit_2121(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2130A)
);

ninexnine_unit ninexnine_unit_2122(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2230A)
);

ninexnine_unit ninexnine_unit_2123(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2330A)
);

ninexnine_unit ninexnine_unit_2124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2430A)
);

ninexnine_unit ninexnine_unit_2125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2530A)
);

ninexnine_unit ninexnine_unit_2126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2630A)
);

ninexnine_unit ninexnine_unit_2127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2730A)
);

assign C230A=c2030A+c2130A+c2230A+c2330A+c2430A+c2530A+c2630A+c2730A;
assign A230A=(C230A>=0)?1:0;

assign P330A=A230A;

ninexnine_unit ninexnine_unit_2128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2031A)
);

ninexnine_unit ninexnine_unit_2129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2131A)
);

ninexnine_unit ninexnine_unit_2130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2231A)
);

ninexnine_unit ninexnine_unit_2131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2331A)
);

ninexnine_unit ninexnine_unit_2132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2431A)
);

ninexnine_unit ninexnine_unit_2133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2531A)
);

ninexnine_unit ninexnine_unit_2134(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2631A)
);

ninexnine_unit ninexnine_unit_2135(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2731A)
);

assign C231A=c2031A+c2131A+c2231A+c2331A+c2431A+c2531A+c2631A+c2731A;
assign A231A=(C231A>=0)?1:0;

assign P331A=A231A;

ninexnine_unit ninexnine_unit_2136(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2032A)
);

ninexnine_unit ninexnine_unit_2137(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2132A)
);

ninexnine_unit ninexnine_unit_2138(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2232A)
);

ninexnine_unit ninexnine_unit_2139(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2332A)
);

ninexnine_unit ninexnine_unit_2140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2432A)
);

ninexnine_unit ninexnine_unit_2141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2532A)
);

ninexnine_unit ninexnine_unit_2142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2632A)
);

ninexnine_unit ninexnine_unit_2143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2732A)
);

assign C232A=c2032A+c2132A+c2232A+c2332A+c2432A+c2532A+c2632A+c2732A;
assign A232A=(C232A>=0)?1:0;

assign P332A=A232A;

ninexnine_unit ninexnine_unit_2144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2033A)
);

ninexnine_unit ninexnine_unit_2145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2133A)
);

ninexnine_unit ninexnine_unit_2146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2233A)
);

ninexnine_unit ninexnine_unit_2147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2333A)
);

ninexnine_unit ninexnine_unit_2148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2433A)
);

ninexnine_unit ninexnine_unit_2149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2533A)
);

ninexnine_unit ninexnine_unit_2150(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2633A)
);

ninexnine_unit ninexnine_unit_2151(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2733A)
);

assign C233A=c2033A+c2133A+c2233A+c2333A+c2433A+c2533A+c2633A+c2733A;
assign A233A=(C233A>=0)?1:0;

assign P333A=A233A;

ninexnine_unit ninexnine_unit_2152(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2034A)
);

ninexnine_unit ninexnine_unit_2153(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2134A)
);

ninexnine_unit ninexnine_unit_2154(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2234A)
);

ninexnine_unit ninexnine_unit_2155(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2334A)
);

ninexnine_unit ninexnine_unit_2156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2434A)
);

ninexnine_unit ninexnine_unit_2157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2534A)
);

ninexnine_unit ninexnine_unit_2158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2634A)
);

ninexnine_unit ninexnine_unit_2159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2734A)
);

assign C234A=c2034A+c2134A+c2234A+c2334A+c2434A+c2534A+c2634A+c2734A;
assign A234A=(C234A>=0)?1:0;

assign P334A=A234A;

ninexnine_unit ninexnine_unit_2160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2040A)
);

ninexnine_unit ninexnine_unit_2161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2140A)
);

ninexnine_unit ninexnine_unit_2162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2240A)
);

ninexnine_unit ninexnine_unit_2163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2340A)
);

ninexnine_unit ninexnine_unit_2164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2440A)
);

ninexnine_unit ninexnine_unit_2165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2540A)
);

ninexnine_unit ninexnine_unit_2166(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2640A)
);

ninexnine_unit ninexnine_unit_2167(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2740A)
);

assign C240A=c2040A+c2140A+c2240A+c2340A+c2440A+c2540A+c2640A+c2740A;
assign A240A=(C240A>=0)?1:0;

assign P340A=A240A;

ninexnine_unit ninexnine_unit_2168(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2041A)
);

ninexnine_unit ninexnine_unit_2169(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2141A)
);

ninexnine_unit ninexnine_unit_2170(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2241A)
);

ninexnine_unit ninexnine_unit_2171(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2341A)
);

ninexnine_unit ninexnine_unit_2172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2441A)
);

ninexnine_unit ninexnine_unit_2173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2541A)
);

ninexnine_unit ninexnine_unit_2174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2641A)
);

ninexnine_unit ninexnine_unit_2175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2741A)
);

assign C241A=c2041A+c2141A+c2241A+c2341A+c2441A+c2541A+c2641A+c2741A;
assign A241A=(C241A>=0)?1:0;

assign P341A=A241A;

ninexnine_unit ninexnine_unit_2176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2042A)
);

ninexnine_unit ninexnine_unit_2177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2142A)
);

ninexnine_unit ninexnine_unit_2178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2242A)
);

ninexnine_unit ninexnine_unit_2179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2342A)
);

ninexnine_unit ninexnine_unit_2180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2442A)
);

ninexnine_unit ninexnine_unit_2181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2542A)
);

ninexnine_unit ninexnine_unit_2182(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2642A)
);

ninexnine_unit ninexnine_unit_2183(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2742A)
);

assign C242A=c2042A+c2142A+c2242A+c2342A+c2442A+c2542A+c2642A+c2742A;
assign A242A=(C242A>=0)?1:0;

assign P342A=A242A;

ninexnine_unit ninexnine_unit_2184(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2043A)
);

ninexnine_unit ninexnine_unit_2185(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2143A)
);

ninexnine_unit ninexnine_unit_2186(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2243A)
);

ninexnine_unit ninexnine_unit_2187(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2343A)
);

ninexnine_unit ninexnine_unit_2188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2443A)
);

ninexnine_unit ninexnine_unit_2189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2543A)
);

ninexnine_unit ninexnine_unit_2190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2643A)
);

ninexnine_unit ninexnine_unit_2191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2743A)
);

assign C243A=c2043A+c2143A+c2243A+c2343A+c2443A+c2543A+c2643A+c2743A;
assign A243A=(C243A>=0)?1:0;

assign P343A=A243A;

ninexnine_unit ninexnine_unit_2192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2044A)
);

ninexnine_unit ninexnine_unit_2193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2144A)
);

ninexnine_unit ninexnine_unit_2194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2244A)
);

ninexnine_unit ninexnine_unit_2195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2344A)
);

ninexnine_unit ninexnine_unit_2196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2444A)
);

ninexnine_unit ninexnine_unit_2197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2544A)
);

ninexnine_unit ninexnine_unit_2198(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2644A)
);

ninexnine_unit ninexnine_unit_2199(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2744A)
);

assign C244A=c2044A+c2144A+c2244A+c2344A+c2444A+c2544A+c2644A+c2744A;
assign A244A=(C244A>=0)?1:0;

assign P344A=A244A;

ninexnine_unit ninexnine_unit_2200(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2000B)
);

ninexnine_unit ninexnine_unit_2201(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2100B)
);

ninexnine_unit ninexnine_unit_2202(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2200B)
);

ninexnine_unit ninexnine_unit_2203(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2300B)
);

ninexnine_unit ninexnine_unit_2204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2400B)
);

ninexnine_unit ninexnine_unit_2205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2500B)
);

ninexnine_unit ninexnine_unit_2206(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2600B)
);

ninexnine_unit ninexnine_unit_2207(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2700B)
);

assign C200B=c2000B+c2100B+c2200B+c2300B+c2400B+c2500B+c2600B+c2700B;
assign A200B=(C200B>=0)?1:0;

assign P300B=A200B;

ninexnine_unit ninexnine_unit_2208(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2001B)
);

ninexnine_unit ninexnine_unit_2209(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2101B)
);

ninexnine_unit ninexnine_unit_2210(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2201B)
);

ninexnine_unit ninexnine_unit_2211(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2301B)
);

ninexnine_unit ninexnine_unit_2212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2401B)
);

ninexnine_unit ninexnine_unit_2213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2501B)
);

ninexnine_unit ninexnine_unit_2214(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2601B)
);

ninexnine_unit ninexnine_unit_2215(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2701B)
);

assign C201B=c2001B+c2101B+c2201B+c2301B+c2401B+c2501B+c2601B+c2701B;
assign A201B=(C201B>=0)?1:0;

assign P301B=A201B;

ninexnine_unit ninexnine_unit_2216(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2002B)
);

ninexnine_unit ninexnine_unit_2217(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2102B)
);

ninexnine_unit ninexnine_unit_2218(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2202B)
);

ninexnine_unit ninexnine_unit_2219(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2302B)
);

ninexnine_unit ninexnine_unit_2220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2402B)
);

ninexnine_unit ninexnine_unit_2221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2502B)
);

ninexnine_unit ninexnine_unit_2222(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2602B)
);

ninexnine_unit ninexnine_unit_2223(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2702B)
);

assign C202B=c2002B+c2102B+c2202B+c2302B+c2402B+c2502B+c2602B+c2702B;
assign A202B=(C202B>=0)?1:0;

assign P302B=A202B;

ninexnine_unit ninexnine_unit_2224(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2003B)
);

ninexnine_unit ninexnine_unit_2225(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2103B)
);

ninexnine_unit ninexnine_unit_2226(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2203B)
);

ninexnine_unit ninexnine_unit_2227(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2303B)
);

ninexnine_unit ninexnine_unit_2228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2403B)
);

ninexnine_unit ninexnine_unit_2229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2503B)
);

ninexnine_unit ninexnine_unit_2230(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2603B)
);

ninexnine_unit ninexnine_unit_2231(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2703B)
);

assign C203B=c2003B+c2103B+c2203B+c2303B+c2403B+c2503B+c2603B+c2703B;
assign A203B=(C203B>=0)?1:0;

assign P303B=A203B;

ninexnine_unit ninexnine_unit_2232(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2004B)
);

ninexnine_unit ninexnine_unit_2233(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2104B)
);

ninexnine_unit ninexnine_unit_2234(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2204B)
);

ninexnine_unit ninexnine_unit_2235(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2304B)
);

ninexnine_unit ninexnine_unit_2236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2404B)
);

ninexnine_unit ninexnine_unit_2237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2504B)
);

ninexnine_unit ninexnine_unit_2238(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2604B)
);

ninexnine_unit ninexnine_unit_2239(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2704B)
);

assign C204B=c2004B+c2104B+c2204B+c2304B+c2404B+c2504B+c2604B+c2704B;
assign A204B=(C204B>=0)?1:0;

assign P304B=A204B;

ninexnine_unit ninexnine_unit_2240(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2010B)
);

ninexnine_unit ninexnine_unit_2241(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2110B)
);

ninexnine_unit ninexnine_unit_2242(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2210B)
);

ninexnine_unit ninexnine_unit_2243(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2310B)
);

ninexnine_unit ninexnine_unit_2244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2410B)
);

ninexnine_unit ninexnine_unit_2245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2510B)
);

ninexnine_unit ninexnine_unit_2246(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2610B)
);

ninexnine_unit ninexnine_unit_2247(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2710B)
);

assign C210B=c2010B+c2110B+c2210B+c2310B+c2410B+c2510B+c2610B+c2710B;
assign A210B=(C210B>=0)?1:0;

assign P310B=A210B;

ninexnine_unit ninexnine_unit_2248(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2011B)
);

ninexnine_unit ninexnine_unit_2249(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2111B)
);

ninexnine_unit ninexnine_unit_2250(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2211B)
);

ninexnine_unit ninexnine_unit_2251(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2311B)
);

ninexnine_unit ninexnine_unit_2252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2411B)
);

ninexnine_unit ninexnine_unit_2253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2511B)
);

ninexnine_unit ninexnine_unit_2254(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2611B)
);

ninexnine_unit ninexnine_unit_2255(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2711B)
);

assign C211B=c2011B+c2111B+c2211B+c2311B+c2411B+c2511B+c2611B+c2711B;
assign A211B=(C211B>=0)?1:0;

assign P311B=A211B;

ninexnine_unit ninexnine_unit_2256(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2012B)
);

ninexnine_unit ninexnine_unit_2257(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2112B)
);

ninexnine_unit ninexnine_unit_2258(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2212B)
);

ninexnine_unit ninexnine_unit_2259(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2312B)
);

ninexnine_unit ninexnine_unit_2260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2412B)
);

ninexnine_unit ninexnine_unit_2261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2512B)
);

ninexnine_unit ninexnine_unit_2262(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2612B)
);

ninexnine_unit ninexnine_unit_2263(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2712B)
);

assign C212B=c2012B+c2112B+c2212B+c2312B+c2412B+c2512B+c2612B+c2712B;
assign A212B=(C212B>=0)?1:0;

assign P312B=A212B;

ninexnine_unit ninexnine_unit_2264(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2013B)
);

ninexnine_unit ninexnine_unit_2265(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2113B)
);

ninexnine_unit ninexnine_unit_2266(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2213B)
);

ninexnine_unit ninexnine_unit_2267(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2313B)
);

ninexnine_unit ninexnine_unit_2268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2413B)
);

ninexnine_unit ninexnine_unit_2269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2513B)
);

ninexnine_unit ninexnine_unit_2270(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2613B)
);

ninexnine_unit ninexnine_unit_2271(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2713B)
);

assign C213B=c2013B+c2113B+c2213B+c2313B+c2413B+c2513B+c2613B+c2713B;
assign A213B=(C213B>=0)?1:0;

assign P313B=A213B;

ninexnine_unit ninexnine_unit_2272(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2014B)
);

ninexnine_unit ninexnine_unit_2273(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2114B)
);

ninexnine_unit ninexnine_unit_2274(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2214B)
);

ninexnine_unit ninexnine_unit_2275(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2314B)
);

ninexnine_unit ninexnine_unit_2276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2414B)
);

ninexnine_unit ninexnine_unit_2277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2514B)
);

ninexnine_unit ninexnine_unit_2278(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2614B)
);

ninexnine_unit ninexnine_unit_2279(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2714B)
);

assign C214B=c2014B+c2114B+c2214B+c2314B+c2414B+c2514B+c2614B+c2714B;
assign A214B=(C214B>=0)?1:0;

assign P314B=A214B;

ninexnine_unit ninexnine_unit_2280(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2020B)
);

ninexnine_unit ninexnine_unit_2281(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2120B)
);

ninexnine_unit ninexnine_unit_2282(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2220B)
);

ninexnine_unit ninexnine_unit_2283(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2320B)
);

ninexnine_unit ninexnine_unit_2284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2420B)
);

ninexnine_unit ninexnine_unit_2285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2520B)
);

ninexnine_unit ninexnine_unit_2286(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2620B)
);

ninexnine_unit ninexnine_unit_2287(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2720B)
);

assign C220B=c2020B+c2120B+c2220B+c2320B+c2420B+c2520B+c2620B+c2720B;
assign A220B=(C220B>=0)?1:0;

assign P320B=A220B;

ninexnine_unit ninexnine_unit_2288(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2021B)
);

ninexnine_unit ninexnine_unit_2289(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2121B)
);

ninexnine_unit ninexnine_unit_2290(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2221B)
);

ninexnine_unit ninexnine_unit_2291(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2321B)
);

ninexnine_unit ninexnine_unit_2292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2421B)
);

ninexnine_unit ninexnine_unit_2293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2521B)
);

ninexnine_unit ninexnine_unit_2294(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2621B)
);

ninexnine_unit ninexnine_unit_2295(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2721B)
);

assign C221B=c2021B+c2121B+c2221B+c2321B+c2421B+c2521B+c2621B+c2721B;
assign A221B=(C221B>=0)?1:0;

assign P321B=A221B;

ninexnine_unit ninexnine_unit_2296(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2022B)
);

ninexnine_unit ninexnine_unit_2297(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2122B)
);

ninexnine_unit ninexnine_unit_2298(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2222B)
);

ninexnine_unit ninexnine_unit_2299(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2322B)
);

ninexnine_unit ninexnine_unit_2300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2422B)
);

ninexnine_unit ninexnine_unit_2301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2522B)
);

ninexnine_unit ninexnine_unit_2302(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2622B)
);

ninexnine_unit ninexnine_unit_2303(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2722B)
);

assign C222B=c2022B+c2122B+c2222B+c2322B+c2422B+c2522B+c2622B+c2722B;
assign A222B=(C222B>=0)?1:0;

assign P322B=A222B;

ninexnine_unit ninexnine_unit_2304(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2023B)
);

ninexnine_unit ninexnine_unit_2305(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2123B)
);

ninexnine_unit ninexnine_unit_2306(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2223B)
);

ninexnine_unit ninexnine_unit_2307(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2323B)
);

ninexnine_unit ninexnine_unit_2308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2423B)
);

ninexnine_unit ninexnine_unit_2309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2523B)
);

ninexnine_unit ninexnine_unit_2310(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2623B)
);

ninexnine_unit ninexnine_unit_2311(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2723B)
);

assign C223B=c2023B+c2123B+c2223B+c2323B+c2423B+c2523B+c2623B+c2723B;
assign A223B=(C223B>=0)?1:0;

assign P323B=A223B;

ninexnine_unit ninexnine_unit_2312(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2024B)
);

ninexnine_unit ninexnine_unit_2313(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2124B)
);

ninexnine_unit ninexnine_unit_2314(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2224B)
);

ninexnine_unit ninexnine_unit_2315(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2324B)
);

ninexnine_unit ninexnine_unit_2316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2424B)
);

ninexnine_unit ninexnine_unit_2317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2524B)
);

ninexnine_unit ninexnine_unit_2318(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2624B)
);

ninexnine_unit ninexnine_unit_2319(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2724B)
);

assign C224B=c2024B+c2124B+c2224B+c2324B+c2424B+c2524B+c2624B+c2724B;
assign A224B=(C224B>=0)?1:0;

assign P324B=A224B;

ninexnine_unit ninexnine_unit_2320(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2030B)
);

ninexnine_unit ninexnine_unit_2321(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2130B)
);

ninexnine_unit ninexnine_unit_2322(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2230B)
);

ninexnine_unit ninexnine_unit_2323(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2330B)
);

ninexnine_unit ninexnine_unit_2324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2430B)
);

ninexnine_unit ninexnine_unit_2325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2530B)
);

ninexnine_unit ninexnine_unit_2326(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2630B)
);

ninexnine_unit ninexnine_unit_2327(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2730B)
);

assign C230B=c2030B+c2130B+c2230B+c2330B+c2430B+c2530B+c2630B+c2730B;
assign A230B=(C230B>=0)?1:0;

assign P330B=A230B;

ninexnine_unit ninexnine_unit_2328(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2031B)
);

ninexnine_unit ninexnine_unit_2329(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2131B)
);

ninexnine_unit ninexnine_unit_2330(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2231B)
);

ninexnine_unit ninexnine_unit_2331(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2331B)
);

ninexnine_unit ninexnine_unit_2332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2431B)
);

ninexnine_unit ninexnine_unit_2333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2531B)
);

ninexnine_unit ninexnine_unit_2334(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2631B)
);

ninexnine_unit ninexnine_unit_2335(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2731B)
);

assign C231B=c2031B+c2131B+c2231B+c2331B+c2431B+c2531B+c2631B+c2731B;
assign A231B=(C231B>=0)?1:0;

assign P331B=A231B;

ninexnine_unit ninexnine_unit_2336(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2032B)
);

ninexnine_unit ninexnine_unit_2337(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2132B)
);

ninexnine_unit ninexnine_unit_2338(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2232B)
);

ninexnine_unit ninexnine_unit_2339(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2332B)
);

ninexnine_unit ninexnine_unit_2340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2432B)
);

ninexnine_unit ninexnine_unit_2341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2532B)
);

ninexnine_unit ninexnine_unit_2342(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2632B)
);

ninexnine_unit ninexnine_unit_2343(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2732B)
);

assign C232B=c2032B+c2132B+c2232B+c2332B+c2432B+c2532B+c2632B+c2732B;
assign A232B=(C232B>=0)?1:0;

assign P332B=A232B;

ninexnine_unit ninexnine_unit_2344(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2033B)
);

ninexnine_unit ninexnine_unit_2345(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2133B)
);

ninexnine_unit ninexnine_unit_2346(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2233B)
);

ninexnine_unit ninexnine_unit_2347(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2333B)
);

ninexnine_unit ninexnine_unit_2348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2433B)
);

ninexnine_unit ninexnine_unit_2349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2533B)
);

ninexnine_unit ninexnine_unit_2350(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2633B)
);

ninexnine_unit ninexnine_unit_2351(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2733B)
);

assign C233B=c2033B+c2133B+c2233B+c2333B+c2433B+c2533B+c2633B+c2733B;
assign A233B=(C233B>=0)?1:0;

assign P333B=A233B;

ninexnine_unit ninexnine_unit_2352(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2034B)
);

ninexnine_unit ninexnine_unit_2353(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2134B)
);

ninexnine_unit ninexnine_unit_2354(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2234B)
);

ninexnine_unit ninexnine_unit_2355(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2334B)
);

ninexnine_unit ninexnine_unit_2356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2434B)
);

ninexnine_unit ninexnine_unit_2357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2534B)
);

ninexnine_unit ninexnine_unit_2358(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2634B)
);

ninexnine_unit ninexnine_unit_2359(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2734B)
);

assign C234B=c2034B+c2134B+c2234B+c2334B+c2434B+c2534B+c2634B+c2734B;
assign A234B=(C234B>=0)?1:0;

assign P334B=A234B;

ninexnine_unit ninexnine_unit_2360(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2040B)
);

ninexnine_unit ninexnine_unit_2361(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2140B)
);

ninexnine_unit ninexnine_unit_2362(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2240B)
);

ninexnine_unit ninexnine_unit_2363(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2340B)
);

ninexnine_unit ninexnine_unit_2364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2440B)
);

ninexnine_unit ninexnine_unit_2365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2540B)
);

ninexnine_unit ninexnine_unit_2366(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2640B)
);

ninexnine_unit ninexnine_unit_2367(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2740B)
);

assign C240B=c2040B+c2140B+c2240B+c2340B+c2440B+c2540B+c2640B+c2740B;
assign A240B=(C240B>=0)?1:0;

assign P340B=A240B;

ninexnine_unit ninexnine_unit_2368(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2041B)
);

ninexnine_unit ninexnine_unit_2369(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2141B)
);

ninexnine_unit ninexnine_unit_2370(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2241B)
);

ninexnine_unit ninexnine_unit_2371(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2341B)
);

ninexnine_unit ninexnine_unit_2372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2441B)
);

ninexnine_unit ninexnine_unit_2373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2541B)
);

ninexnine_unit ninexnine_unit_2374(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2641B)
);

ninexnine_unit ninexnine_unit_2375(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2741B)
);

assign C241B=c2041B+c2141B+c2241B+c2341B+c2441B+c2541B+c2641B+c2741B;
assign A241B=(C241B>=0)?1:0;

assign P341B=A241B;

ninexnine_unit ninexnine_unit_2376(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2042B)
);

ninexnine_unit ninexnine_unit_2377(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2142B)
);

ninexnine_unit ninexnine_unit_2378(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2242B)
);

ninexnine_unit ninexnine_unit_2379(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2342B)
);

ninexnine_unit ninexnine_unit_2380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2442B)
);

ninexnine_unit ninexnine_unit_2381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2542B)
);

ninexnine_unit ninexnine_unit_2382(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2642B)
);

ninexnine_unit ninexnine_unit_2383(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2742B)
);

assign C242B=c2042B+c2142B+c2242B+c2342B+c2442B+c2542B+c2642B+c2742B;
assign A242B=(C242B>=0)?1:0;

assign P342B=A242B;

ninexnine_unit ninexnine_unit_2384(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2043B)
);

ninexnine_unit ninexnine_unit_2385(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2143B)
);

ninexnine_unit ninexnine_unit_2386(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2243B)
);

ninexnine_unit ninexnine_unit_2387(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2343B)
);

ninexnine_unit ninexnine_unit_2388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2443B)
);

ninexnine_unit ninexnine_unit_2389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2543B)
);

ninexnine_unit ninexnine_unit_2390(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2643B)
);

ninexnine_unit ninexnine_unit_2391(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2743B)
);

assign C243B=c2043B+c2143B+c2243B+c2343B+c2443B+c2543B+c2643B+c2743B;
assign A243B=(C243B>=0)?1:0;

assign P343B=A243B;

ninexnine_unit ninexnine_unit_2392(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2044B)
);

ninexnine_unit ninexnine_unit_2393(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2144B)
);

ninexnine_unit ninexnine_unit_2394(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2244B)
);

ninexnine_unit ninexnine_unit_2395(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2344B)
);

ninexnine_unit ninexnine_unit_2396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2444B)
);

ninexnine_unit ninexnine_unit_2397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2544B)
);

ninexnine_unit ninexnine_unit_2398(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2644B)
);

ninexnine_unit ninexnine_unit_2399(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2744B)
);

assign C244B=c2044B+c2144B+c2244B+c2344B+c2444B+c2544B+c2644B+c2744B;
assign A244B=(C244B>=0)?1:0;

assign P344B=A244B;

ninexnine_unit ninexnine_unit_2400(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2000C)
);

ninexnine_unit ninexnine_unit_2401(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2100C)
);

ninexnine_unit ninexnine_unit_2402(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2200C)
);

ninexnine_unit ninexnine_unit_2403(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2300C)
);

ninexnine_unit ninexnine_unit_2404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2400C)
);

ninexnine_unit ninexnine_unit_2405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2500C)
);

ninexnine_unit ninexnine_unit_2406(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2600C)
);

ninexnine_unit ninexnine_unit_2407(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2700C)
);

assign C200C=c2000C+c2100C+c2200C+c2300C+c2400C+c2500C+c2600C+c2700C;
assign A200C=(C200C>=0)?1:0;

assign P300C=A200C;

ninexnine_unit ninexnine_unit_2408(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2001C)
);

ninexnine_unit ninexnine_unit_2409(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2101C)
);

ninexnine_unit ninexnine_unit_2410(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2201C)
);

ninexnine_unit ninexnine_unit_2411(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2301C)
);

ninexnine_unit ninexnine_unit_2412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2401C)
);

ninexnine_unit ninexnine_unit_2413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2501C)
);

ninexnine_unit ninexnine_unit_2414(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2601C)
);

ninexnine_unit ninexnine_unit_2415(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2701C)
);

assign C201C=c2001C+c2101C+c2201C+c2301C+c2401C+c2501C+c2601C+c2701C;
assign A201C=(C201C>=0)?1:0;

assign P301C=A201C;

ninexnine_unit ninexnine_unit_2416(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2002C)
);

ninexnine_unit ninexnine_unit_2417(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2102C)
);

ninexnine_unit ninexnine_unit_2418(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2202C)
);

ninexnine_unit ninexnine_unit_2419(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2302C)
);

ninexnine_unit ninexnine_unit_2420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2402C)
);

ninexnine_unit ninexnine_unit_2421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2502C)
);

ninexnine_unit ninexnine_unit_2422(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2602C)
);

ninexnine_unit ninexnine_unit_2423(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2702C)
);

assign C202C=c2002C+c2102C+c2202C+c2302C+c2402C+c2502C+c2602C+c2702C;
assign A202C=(C202C>=0)?1:0;

assign P302C=A202C;

ninexnine_unit ninexnine_unit_2424(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2003C)
);

ninexnine_unit ninexnine_unit_2425(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2103C)
);

ninexnine_unit ninexnine_unit_2426(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2203C)
);

ninexnine_unit ninexnine_unit_2427(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2303C)
);

ninexnine_unit ninexnine_unit_2428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2403C)
);

ninexnine_unit ninexnine_unit_2429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2503C)
);

ninexnine_unit ninexnine_unit_2430(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2603C)
);

ninexnine_unit ninexnine_unit_2431(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2703C)
);

assign C203C=c2003C+c2103C+c2203C+c2303C+c2403C+c2503C+c2603C+c2703C;
assign A203C=(C203C>=0)?1:0;

assign P303C=A203C;

ninexnine_unit ninexnine_unit_2432(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2004C)
);

ninexnine_unit ninexnine_unit_2433(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2104C)
);

ninexnine_unit ninexnine_unit_2434(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2204C)
);

ninexnine_unit ninexnine_unit_2435(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2304C)
);

ninexnine_unit ninexnine_unit_2436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2404C)
);

ninexnine_unit ninexnine_unit_2437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2504C)
);

ninexnine_unit ninexnine_unit_2438(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2604C)
);

ninexnine_unit ninexnine_unit_2439(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2704C)
);

assign C204C=c2004C+c2104C+c2204C+c2304C+c2404C+c2504C+c2604C+c2704C;
assign A204C=(C204C>=0)?1:0;

assign P304C=A204C;

ninexnine_unit ninexnine_unit_2440(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2010C)
);

ninexnine_unit ninexnine_unit_2441(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2110C)
);

ninexnine_unit ninexnine_unit_2442(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2210C)
);

ninexnine_unit ninexnine_unit_2443(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2310C)
);

ninexnine_unit ninexnine_unit_2444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2410C)
);

ninexnine_unit ninexnine_unit_2445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2510C)
);

ninexnine_unit ninexnine_unit_2446(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2610C)
);

ninexnine_unit ninexnine_unit_2447(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2710C)
);

assign C210C=c2010C+c2110C+c2210C+c2310C+c2410C+c2510C+c2610C+c2710C;
assign A210C=(C210C>=0)?1:0;

assign P310C=A210C;

ninexnine_unit ninexnine_unit_2448(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2011C)
);

ninexnine_unit ninexnine_unit_2449(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2111C)
);

ninexnine_unit ninexnine_unit_2450(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2211C)
);

ninexnine_unit ninexnine_unit_2451(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2311C)
);

ninexnine_unit ninexnine_unit_2452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2411C)
);

ninexnine_unit ninexnine_unit_2453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2511C)
);

ninexnine_unit ninexnine_unit_2454(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2611C)
);

ninexnine_unit ninexnine_unit_2455(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2711C)
);

assign C211C=c2011C+c2111C+c2211C+c2311C+c2411C+c2511C+c2611C+c2711C;
assign A211C=(C211C>=0)?1:0;

assign P311C=A211C;

ninexnine_unit ninexnine_unit_2456(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2012C)
);

ninexnine_unit ninexnine_unit_2457(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2112C)
);

ninexnine_unit ninexnine_unit_2458(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2212C)
);

ninexnine_unit ninexnine_unit_2459(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2312C)
);

ninexnine_unit ninexnine_unit_2460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2412C)
);

ninexnine_unit ninexnine_unit_2461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2512C)
);

ninexnine_unit ninexnine_unit_2462(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2612C)
);

ninexnine_unit ninexnine_unit_2463(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2712C)
);

assign C212C=c2012C+c2112C+c2212C+c2312C+c2412C+c2512C+c2612C+c2712C;
assign A212C=(C212C>=0)?1:0;

assign P312C=A212C;

ninexnine_unit ninexnine_unit_2464(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2013C)
);

ninexnine_unit ninexnine_unit_2465(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2113C)
);

ninexnine_unit ninexnine_unit_2466(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2213C)
);

ninexnine_unit ninexnine_unit_2467(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2313C)
);

ninexnine_unit ninexnine_unit_2468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2413C)
);

ninexnine_unit ninexnine_unit_2469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2513C)
);

ninexnine_unit ninexnine_unit_2470(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2613C)
);

ninexnine_unit ninexnine_unit_2471(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2713C)
);

assign C213C=c2013C+c2113C+c2213C+c2313C+c2413C+c2513C+c2613C+c2713C;
assign A213C=(C213C>=0)?1:0;

assign P313C=A213C;

ninexnine_unit ninexnine_unit_2472(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2014C)
);

ninexnine_unit ninexnine_unit_2473(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2114C)
);

ninexnine_unit ninexnine_unit_2474(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2214C)
);

ninexnine_unit ninexnine_unit_2475(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2314C)
);

ninexnine_unit ninexnine_unit_2476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2414C)
);

ninexnine_unit ninexnine_unit_2477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2514C)
);

ninexnine_unit ninexnine_unit_2478(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2614C)
);

ninexnine_unit ninexnine_unit_2479(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2714C)
);

assign C214C=c2014C+c2114C+c2214C+c2314C+c2414C+c2514C+c2614C+c2714C;
assign A214C=(C214C>=0)?1:0;

assign P314C=A214C;

ninexnine_unit ninexnine_unit_2480(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2020C)
);

ninexnine_unit ninexnine_unit_2481(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2120C)
);

ninexnine_unit ninexnine_unit_2482(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2220C)
);

ninexnine_unit ninexnine_unit_2483(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2320C)
);

ninexnine_unit ninexnine_unit_2484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2420C)
);

ninexnine_unit ninexnine_unit_2485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2520C)
);

ninexnine_unit ninexnine_unit_2486(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2620C)
);

ninexnine_unit ninexnine_unit_2487(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2720C)
);

assign C220C=c2020C+c2120C+c2220C+c2320C+c2420C+c2520C+c2620C+c2720C;
assign A220C=(C220C>=0)?1:0;

assign P320C=A220C;

ninexnine_unit ninexnine_unit_2488(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2021C)
);

ninexnine_unit ninexnine_unit_2489(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2121C)
);

ninexnine_unit ninexnine_unit_2490(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2221C)
);

ninexnine_unit ninexnine_unit_2491(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2321C)
);

ninexnine_unit ninexnine_unit_2492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2421C)
);

ninexnine_unit ninexnine_unit_2493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2521C)
);

ninexnine_unit ninexnine_unit_2494(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2621C)
);

ninexnine_unit ninexnine_unit_2495(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2721C)
);

assign C221C=c2021C+c2121C+c2221C+c2321C+c2421C+c2521C+c2621C+c2721C;
assign A221C=(C221C>=0)?1:0;

assign P321C=A221C;

ninexnine_unit ninexnine_unit_2496(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2022C)
);

ninexnine_unit ninexnine_unit_2497(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2122C)
);

ninexnine_unit ninexnine_unit_2498(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2222C)
);

ninexnine_unit ninexnine_unit_2499(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2322C)
);

ninexnine_unit ninexnine_unit_2500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2422C)
);

ninexnine_unit ninexnine_unit_2501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2522C)
);

ninexnine_unit ninexnine_unit_2502(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2622C)
);

ninexnine_unit ninexnine_unit_2503(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2722C)
);

assign C222C=c2022C+c2122C+c2222C+c2322C+c2422C+c2522C+c2622C+c2722C;
assign A222C=(C222C>=0)?1:0;

assign P322C=A222C;

ninexnine_unit ninexnine_unit_2504(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2023C)
);

ninexnine_unit ninexnine_unit_2505(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2123C)
);

ninexnine_unit ninexnine_unit_2506(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2223C)
);

ninexnine_unit ninexnine_unit_2507(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2323C)
);

ninexnine_unit ninexnine_unit_2508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2423C)
);

ninexnine_unit ninexnine_unit_2509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2523C)
);

ninexnine_unit ninexnine_unit_2510(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2623C)
);

ninexnine_unit ninexnine_unit_2511(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2723C)
);

assign C223C=c2023C+c2123C+c2223C+c2323C+c2423C+c2523C+c2623C+c2723C;
assign A223C=(C223C>=0)?1:0;

assign P323C=A223C;

ninexnine_unit ninexnine_unit_2512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2024C)
);

ninexnine_unit ninexnine_unit_2513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2124C)
);

ninexnine_unit ninexnine_unit_2514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2224C)
);

ninexnine_unit ninexnine_unit_2515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2324C)
);

ninexnine_unit ninexnine_unit_2516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2424C)
);

ninexnine_unit ninexnine_unit_2517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2524C)
);

ninexnine_unit ninexnine_unit_2518(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2624C)
);

ninexnine_unit ninexnine_unit_2519(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2724C)
);

assign C224C=c2024C+c2124C+c2224C+c2324C+c2424C+c2524C+c2624C+c2724C;
assign A224C=(C224C>=0)?1:0;

assign P324C=A224C;

ninexnine_unit ninexnine_unit_2520(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2030C)
);

ninexnine_unit ninexnine_unit_2521(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2130C)
);

ninexnine_unit ninexnine_unit_2522(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2230C)
);

ninexnine_unit ninexnine_unit_2523(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2330C)
);

ninexnine_unit ninexnine_unit_2524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2430C)
);

ninexnine_unit ninexnine_unit_2525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2530C)
);

ninexnine_unit ninexnine_unit_2526(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2630C)
);

ninexnine_unit ninexnine_unit_2527(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2730C)
);

assign C230C=c2030C+c2130C+c2230C+c2330C+c2430C+c2530C+c2630C+c2730C;
assign A230C=(C230C>=0)?1:0;

assign P330C=A230C;

ninexnine_unit ninexnine_unit_2528(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2031C)
);

ninexnine_unit ninexnine_unit_2529(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2131C)
);

ninexnine_unit ninexnine_unit_2530(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2231C)
);

ninexnine_unit ninexnine_unit_2531(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2331C)
);

ninexnine_unit ninexnine_unit_2532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2431C)
);

ninexnine_unit ninexnine_unit_2533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2531C)
);

ninexnine_unit ninexnine_unit_2534(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2631C)
);

ninexnine_unit ninexnine_unit_2535(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2731C)
);

assign C231C=c2031C+c2131C+c2231C+c2331C+c2431C+c2531C+c2631C+c2731C;
assign A231C=(C231C>=0)?1:0;

assign P331C=A231C;

ninexnine_unit ninexnine_unit_2536(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2032C)
);

ninexnine_unit ninexnine_unit_2537(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2132C)
);

ninexnine_unit ninexnine_unit_2538(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2232C)
);

ninexnine_unit ninexnine_unit_2539(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2332C)
);

ninexnine_unit ninexnine_unit_2540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2432C)
);

ninexnine_unit ninexnine_unit_2541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2532C)
);

ninexnine_unit ninexnine_unit_2542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2632C)
);

ninexnine_unit ninexnine_unit_2543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2732C)
);

assign C232C=c2032C+c2132C+c2232C+c2332C+c2432C+c2532C+c2632C+c2732C;
assign A232C=(C232C>=0)?1:0;

assign P332C=A232C;

ninexnine_unit ninexnine_unit_2544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2033C)
);

ninexnine_unit ninexnine_unit_2545(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2133C)
);

ninexnine_unit ninexnine_unit_2546(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2233C)
);

ninexnine_unit ninexnine_unit_2547(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2333C)
);

ninexnine_unit ninexnine_unit_2548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2433C)
);

ninexnine_unit ninexnine_unit_2549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2533C)
);

ninexnine_unit ninexnine_unit_2550(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2633C)
);

ninexnine_unit ninexnine_unit_2551(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2733C)
);

assign C233C=c2033C+c2133C+c2233C+c2333C+c2433C+c2533C+c2633C+c2733C;
assign A233C=(C233C>=0)?1:0;

assign P333C=A233C;

ninexnine_unit ninexnine_unit_2552(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2034C)
);

ninexnine_unit ninexnine_unit_2553(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2134C)
);

ninexnine_unit ninexnine_unit_2554(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2234C)
);

ninexnine_unit ninexnine_unit_2555(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2334C)
);

ninexnine_unit ninexnine_unit_2556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2434C)
);

ninexnine_unit ninexnine_unit_2557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2534C)
);

ninexnine_unit ninexnine_unit_2558(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2634C)
);

ninexnine_unit ninexnine_unit_2559(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2734C)
);

assign C234C=c2034C+c2134C+c2234C+c2334C+c2434C+c2534C+c2634C+c2734C;
assign A234C=(C234C>=0)?1:0;

assign P334C=A234C;

ninexnine_unit ninexnine_unit_2560(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2040C)
);

ninexnine_unit ninexnine_unit_2561(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2140C)
);

ninexnine_unit ninexnine_unit_2562(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2240C)
);

ninexnine_unit ninexnine_unit_2563(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2340C)
);

ninexnine_unit ninexnine_unit_2564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2440C)
);

ninexnine_unit ninexnine_unit_2565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2540C)
);

ninexnine_unit ninexnine_unit_2566(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2640C)
);

ninexnine_unit ninexnine_unit_2567(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2740C)
);

assign C240C=c2040C+c2140C+c2240C+c2340C+c2440C+c2540C+c2640C+c2740C;
assign A240C=(C240C>=0)?1:0;

assign P340C=A240C;

ninexnine_unit ninexnine_unit_2568(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2041C)
);

ninexnine_unit ninexnine_unit_2569(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2141C)
);

ninexnine_unit ninexnine_unit_2570(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2241C)
);

ninexnine_unit ninexnine_unit_2571(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2341C)
);

ninexnine_unit ninexnine_unit_2572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2441C)
);

ninexnine_unit ninexnine_unit_2573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2541C)
);

ninexnine_unit ninexnine_unit_2574(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2641C)
);

ninexnine_unit ninexnine_unit_2575(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2741C)
);

assign C241C=c2041C+c2141C+c2241C+c2341C+c2441C+c2541C+c2641C+c2741C;
assign A241C=(C241C>=0)?1:0;

assign P341C=A241C;

ninexnine_unit ninexnine_unit_2576(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2042C)
);

ninexnine_unit ninexnine_unit_2577(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2142C)
);

ninexnine_unit ninexnine_unit_2578(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2242C)
);

ninexnine_unit ninexnine_unit_2579(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2342C)
);

ninexnine_unit ninexnine_unit_2580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2442C)
);

ninexnine_unit ninexnine_unit_2581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2542C)
);

ninexnine_unit ninexnine_unit_2582(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2642C)
);

ninexnine_unit ninexnine_unit_2583(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2742C)
);

assign C242C=c2042C+c2142C+c2242C+c2342C+c2442C+c2542C+c2642C+c2742C;
assign A242C=(C242C>=0)?1:0;

assign P342C=A242C;

ninexnine_unit ninexnine_unit_2584(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2043C)
);

ninexnine_unit ninexnine_unit_2585(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2143C)
);

ninexnine_unit ninexnine_unit_2586(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2243C)
);

ninexnine_unit ninexnine_unit_2587(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2343C)
);

ninexnine_unit ninexnine_unit_2588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2443C)
);

ninexnine_unit ninexnine_unit_2589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2543C)
);

ninexnine_unit ninexnine_unit_2590(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2643C)
);

ninexnine_unit ninexnine_unit_2591(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2743C)
);

assign C243C=c2043C+c2143C+c2243C+c2343C+c2443C+c2543C+c2643C+c2743C;
assign A243C=(C243C>=0)?1:0;

assign P343C=A243C;

ninexnine_unit ninexnine_unit_2592(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2044C)
);

ninexnine_unit ninexnine_unit_2593(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2144C)
);

ninexnine_unit ninexnine_unit_2594(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2244C)
);

ninexnine_unit ninexnine_unit_2595(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2344C)
);

ninexnine_unit ninexnine_unit_2596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2444C)
);

ninexnine_unit ninexnine_unit_2597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2544C)
);

ninexnine_unit ninexnine_unit_2598(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2644C)
);

ninexnine_unit ninexnine_unit_2599(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2744C)
);

assign C244C=c2044C+c2144C+c2244C+c2344C+c2444C+c2544C+c2644C+c2744C;
assign A244C=(C244C>=0)?1:0;

assign P344C=A244C;

ninexnine_unit ninexnine_unit_2600(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2000D)
);

ninexnine_unit ninexnine_unit_2601(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2100D)
);

ninexnine_unit ninexnine_unit_2602(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2200D)
);

ninexnine_unit ninexnine_unit_2603(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2300D)
);

ninexnine_unit ninexnine_unit_2604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2400D)
);

ninexnine_unit ninexnine_unit_2605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2500D)
);

ninexnine_unit ninexnine_unit_2606(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2600D)
);

ninexnine_unit ninexnine_unit_2607(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2700D)
);

assign C200D=c2000D+c2100D+c2200D+c2300D+c2400D+c2500D+c2600D+c2700D;
assign A200D=(C200D>=0)?1:0;

assign P300D=A200D;

ninexnine_unit ninexnine_unit_2608(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2001D)
);

ninexnine_unit ninexnine_unit_2609(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2101D)
);

ninexnine_unit ninexnine_unit_2610(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2201D)
);

ninexnine_unit ninexnine_unit_2611(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2301D)
);

ninexnine_unit ninexnine_unit_2612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2401D)
);

ninexnine_unit ninexnine_unit_2613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2501D)
);

ninexnine_unit ninexnine_unit_2614(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2601D)
);

ninexnine_unit ninexnine_unit_2615(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2701D)
);

assign C201D=c2001D+c2101D+c2201D+c2301D+c2401D+c2501D+c2601D+c2701D;
assign A201D=(C201D>=0)?1:0;

assign P301D=A201D;

ninexnine_unit ninexnine_unit_2616(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2002D)
);

ninexnine_unit ninexnine_unit_2617(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2102D)
);

ninexnine_unit ninexnine_unit_2618(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2202D)
);

ninexnine_unit ninexnine_unit_2619(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2302D)
);

ninexnine_unit ninexnine_unit_2620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2402D)
);

ninexnine_unit ninexnine_unit_2621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2502D)
);

ninexnine_unit ninexnine_unit_2622(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2602D)
);

ninexnine_unit ninexnine_unit_2623(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2702D)
);

assign C202D=c2002D+c2102D+c2202D+c2302D+c2402D+c2502D+c2602D+c2702D;
assign A202D=(C202D>=0)?1:0;

assign P302D=A202D;

ninexnine_unit ninexnine_unit_2624(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2003D)
);

ninexnine_unit ninexnine_unit_2625(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2103D)
);

ninexnine_unit ninexnine_unit_2626(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2203D)
);

ninexnine_unit ninexnine_unit_2627(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2303D)
);

ninexnine_unit ninexnine_unit_2628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2403D)
);

ninexnine_unit ninexnine_unit_2629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2503D)
);

ninexnine_unit ninexnine_unit_2630(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2603D)
);

ninexnine_unit ninexnine_unit_2631(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2703D)
);

assign C203D=c2003D+c2103D+c2203D+c2303D+c2403D+c2503D+c2603D+c2703D;
assign A203D=(C203D>=0)?1:0;

assign P303D=A203D;

ninexnine_unit ninexnine_unit_2632(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2004D)
);

ninexnine_unit ninexnine_unit_2633(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2104D)
);

ninexnine_unit ninexnine_unit_2634(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2204D)
);

ninexnine_unit ninexnine_unit_2635(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2304D)
);

ninexnine_unit ninexnine_unit_2636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2404D)
);

ninexnine_unit ninexnine_unit_2637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2504D)
);

ninexnine_unit ninexnine_unit_2638(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2604D)
);

ninexnine_unit ninexnine_unit_2639(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2704D)
);

assign C204D=c2004D+c2104D+c2204D+c2304D+c2404D+c2504D+c2604D+c2704D;
assign A204D=(C204D>=0)?1:0;

assign P304D=A204D;

ninexnine_unit ninexnine_unit_2640(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2010D)
);

ninexnine_unit ninexnine_unit_2641(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2110D)
);

ninexnine_unit ninexnine_unit_2642(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2210D)
);

ninexnine_unit ninexnine_unit_2643(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2310D)
);

ninexnine_unit ninexnine_unit_2644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2410D)
);

ninexnine_unit ninexnine_unit_2645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2510D)
);

ninexnine_unit ninexnine_unit_2646(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2610D)
);

ninexnine_unit ninexnine_unit_2647(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2710D)
);

assign C210D=c2010D+c2110D+c2210D+c2310D+c2410D+c2510D+c2610D+c2710D;
assign A210D=(C210D>=0)?1:0;

assign P310D=A210D;

ninexnine_unit ninexnine_unit_2648(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2011D)
);

ninexnine_unit ninexnine_unit_2649(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2111D)
);

ninexnine_unit ninexnine_unit_2650(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2211D)
);

ninexnine_unit ninexnine_unit_2651(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2311D)
);

ninexnine_unit ninexnine_unit_2652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2411D)
);

ninexnine_unit ninexnine_unit_2653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2511D)
);

ninexnine_unit ninexnine_unit_2654(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2611D)
);

ninexnine_unit ninexnine_unit_2655(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2711D)
);

assign C211D=c2011D+c2111D+c2211D+c2311D+c2411D+c2511D+c2611D+c2711D;
assign A211D=(C211D>=0)?1:0;

assign P311D=A211D;

ninexnine_unit ninexnine_unit_2656(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2012D)
);

ninexnine_unit ninexnine_unit_2657(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2112D)
);

ninexnine_unit ninexnine_unit_2658(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2212D)
);

ninexnine_unit ninexnine_unit_2659(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2312D)
);

ninexnine_unit ninexnine_unit_2660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2412D)
);

ninexnine_unit ninexnine_unit_2661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2512D)
);

ninexnine_unit ninexnine_unit_2662(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2612D)
);

ninexnine_unit ninexnine_unit_2663(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2712D)
);

assign C212D=c2012D+c2112D+c2212D+c2312D+c2412D+c2512D+c2612D+c2712D;
assign A212D=(C212D>=0)?1:0;

assign P312D=A212D;

ninexnine_unit ninexnine_unit_2664(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2013D)
);

ninexnine_unit ninexnine_unit_2665(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2113D)
);

ninexnine_unit ninexnine_unit_2666(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2213D)
);

ninexnine_unit ninexnine_unit_2667(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2313D)
);

ninexnine_unit ninexnine_unit_2668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2413D)
);

ninexnine_unit ninexnine_unit_2669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2513D)
);

ninexnine_unit ninexnine_unit_2670(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2613D)
);

ninexnine_unit ninexnine_unit_2671(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2713D)
);

assign C213D=c2013D+c2113D+c2213D+c2313D+c2413D+c2513D+c2613D+c2713D;
assign A213D=(C213D>=0)?1:0;

assign P313D=A213D;

ninexnine_unit ninexnine_unit_2672(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2014D)
);

ninexnine_unit ninexnine_unit_2673(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2114D)
);

ninexnine_unit ninexnine_unit_2674(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2214D)
);

ninexnine_unit ninexnine_unit_2675(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2314D)
);

ninexnine_unit ninexnine_unit_2676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2414D)
);

ninexnine_unit ninexnine_unit_2677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2514D)
);

ninexnine_unit ninexnine_unit_2678(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2614D)
);

ninexnine_unit ninexnine_unit_2679(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2714D)
);

assign C214D=c2014D+c2114D+c2214D+c2314D+c2414D+c2514D+c2614D+c2714D;
assign A214D=(C214D>=0)?1:0;

assign P314D=A214D;

ninexnine_unit ninexnine_unit_2680(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2020D)
);

ninexnine_unit ninexnine_unit_2681(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2120D)
);

ninexnine_unit ninexnine_unit_2682(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2220D)
);

ninexnine_unit ninexnine_unit_2683(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2320D)
);

ninexnine_unit ninexnine_unit_2684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2420D)
);

ninexnine_unit ninexnine_unit_2685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2520D)
);

ninexnine_unit ninexnine_unit_2686(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2620D)
);

ninexnine_unit ninexnine_unit_2687(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2720D)
);

assign C220D=c2020D+c2120D+c2220D+c2320D+c2420D+c2520D+c2620D+c2720D;
assign A220D=(C220D>=0)?1:0;

assign P320D=A220D;

ninexnine_unit ninexnine_unit_2688(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2021D)
);

ninexnine_unit ninexnine_unit_2689(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2121D)
);

ninexnine_unit ninexnine_unit_2690(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2221D)
);

ninexnine_unit ninexnine_unit_2691(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2321D)
);

ninexnine_unit ninexnine_unit_2692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2421D)
);

ninexnine_unit ninexnine_unit_2693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2521D)
);

ninexnine_unit ninexnine_unit_2694(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2621D)
);

ninexnine_unit ninexnine_unit_2695(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2721D)
);

assign C221D=c2021D+c2121D+c2221D+c2321D+c2421D+c2521D+c2621D+c2721D;
assign A221D=(C221D>=0)?1:0;

assign P321D=A221D;

ninexnine_unit ninexnine_unit_2696(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2022D)
);

ninexnine_unit ninexnine_unit_2697(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2122D)
);

ninexnine_unit ninexnine_unit_2698(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2222D)
);

ninexnine_unit ninexnine_unit_2699(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2322D)
);

ninexnine_unit ninexnine_unit_2700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2422D)
);

ninexnine_unit ninexnine_unit_2701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2522D)
);

ninexnine_unit ninexnine_unit_2702(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2622D)
);

ninexnine_unit ninexnine_unit_2703(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2722D)
);

assign C222D=c2022D+c2122D+c2222D+c2322D+c2422D+c2522D+c2622D+c2722D;
assign A222D=(C222D>=0)?1:0;

assign P322D=A222D;

ninexnine_unit ninexnine_unit_2704(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2023D)
);

ninexnine_unit ninexnine_unit_2705(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2123D)
);

ninexnine_unit ninexnine_unit_2706(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2223D)
);

ninexnine_unit ninexnine_unit_2707(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2323D)
);

ninexnine_unit ninexnine_unit_2708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2423D)
);

ninexnine_unit ninexnine_unit_2709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2523D)
);

ninexnine_unit ninexnine_unit_2710(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2623D)
);

ninexnine_unit ninexnine_unit_2711(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2723D)
);

assign C223D=c2023D+c2123D+c2223D+c2323D+c2423D+c2523D+c2623D+c2723D;
assign A223D=(C223D>=0)?1:0;

assign P323D=A223D;

ninexnine_unit ninexnine_unit_2712(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2024D)
);

ninexnine_unit ninexnine_unit_2713(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2124D)
);

ninexnine_unit ninexnine_unit_2714(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2224D)
);

ninexnine_unit ninexnine_unit_2715(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2324D)
);

ninexnine_unit ninexnine_unit_2716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2424D)
);

ninexnine_unit ninexnine_unit_2717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2524D)
);

ninexnine_unit ninexnine_unit_2718(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2624D)
);

ninexnine_unit ninexnine_unit_2719(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2724D)
);

assign C224D=c2024D+c2124D+c2224D+c2324D+c2424D+c2524D+c2624D+c2724D;
assign A224D=(C224D>=0)?1:0;

assign P324D=A224D;

ninexnine_unit ninexnine_unit_2720(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2030D)
);

ninexnine_unit ninexnine_unit_2721(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2130D)
);

ninexnine_unit ninexnine_unit_2722(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2230D)
);

ninexnine_unit ninexnine_unit_2723(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2330D)
);

ninexnine_unit ninexnine_unit_2724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2430D)
);

ninexnine_unit ninexnine_unit_2725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2530D)
);

ninexnine_unit ninexnine_unit_2726(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2630D)
);

ninexnine_unit ninexnine_unit_2727(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2730D)
);

assign C230D=c2030D+c2130D+c2230D+c2330D+c2430D+c2530D+c2630D+c2730D;
assign A230D=(C230D>=0)?1:0;

assign P330D=A230D;

ninexnine_unit ninexnine_unit_2728(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2031D)
);

ninexnine_unit ninexnine_unit_2729(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2131D)
);

ninexnine_unit ninexnine_unit_2730(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2231D)
);

ninexnine_unit ninexnine_unit_2731(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2331D)
);

ninexnine_unit ninexnine_unit_2732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2431D)
);

ninexnine_unit ninexnine_unit_2733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2531D)
);

ninexnine_unit ninexnine_unit_2734(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2631D)
);

ninexnine_unit ninexnine_unit_2735(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2731D)
);

assign C231D=c2031D+c2131D+c2231D+c2331D+c2431D+c2531D+c2631D+c2731D;
assign A231D=(C231D>=0)?1:0;

assign P331D=A231D;

ninexnine_unit ninexnine_unit_2736(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2032D)
);

ninexnine_unit ninexnine_unit_2737(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2132D)
);

ninexnine_unit ninexnine_unit_2738(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2232D)
);

ninexnine_unit ninexnine_unit_2739(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2332D)
);

ninexnine_unit ninexnine_unit_2740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2432D)
);

ninexnine_unit ninexnine_unit_2741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2532D)
);

ninexnine_unit ninexnine_unit_2742(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2632D)
);

ninexnine_unit ninexnine_unit_2743(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2732D)
);

assign C232D=c2032D+c2132D+c2232D+c2332D+c2432D+c2532D+c2632D+c2732D;
assign A232D=(C232D>=0)?1:0;

assign P332D=A232D;

ninexnine_unit ninexnine_unit_2744(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2033D)
);

ninexnine_unit ninexnine_unit_2745(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2133D)
);

ninexnine_unit ninexnine_unit_2746(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2233D)
);

ninexnine_unit ninexnine_unit_2747(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2333D)
);

ninexnine_unit ninexnine_unit_2748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2433D)
);

ninexnine_unit ninexnine_unit_2749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2533D)
);

ninexnine_unit ninexnine_unit_2750(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2633D)
);

ninexnine_unit ninexnine_unit_2751(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2733D)
);

assign C233D=c2033D+c2133D+c2233D+c2333D+c2433D+c2533D+c2633D+c2733D;
assign A233D=(C233D>=0)?1:0;

assign P333D=A233D;

ninexnine_unit ninexnine_unit_2752(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2034D)
);

ninexnine_unit ninexnine_unit_2753(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2134D)
);

ninexnine_unit ninexnine_unit_2754(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2234D)
);

ninexnine_unit ninexnine_unit_2755(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2334D)
);

ninexnine_unit ninexnine_unit_2756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2434D)
);

ninexnine_unit ninexnine_unit_2757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2534D)
);

ninexnine_unit ninexnine_unit_2758(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2634D)
);

ninexnine_unit ninexnine_unit_2759(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2734D)
);

assign C234D=c2034D+c2134D+c2234D+c2334D+c2434D+c2534D+c2634D+c2734D;
assign A234D=(C234D>=0)?1:0;

assign P334D=A234D;

ninexnine_unit ninexnine_unit_2760(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2040D)
);

ninexnine_unit ninexnine_unit_2761(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2140D)
);

ninexnine_unit ninexnine_unit_2762(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2240D)
);

ninexnine_unit ninexnine_unit_2763(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2340D)
);

ninexnine_unit ninexnine_unit_2764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2440D)
);

ninexnine_unit ninexnine_unit_2765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2540D)
);

ninexnine_unit ninexnine_unit_2766(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2640D)
);

ninexnine_unit ninexnine_unit_2767(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2740D)
);

assign C240D=c2040D+c2140D+c2240D+c2340D+c2440D+c2540D+c2640D+c2740D;
assign A240D=(C240D>=0)?1:0;

assign P340D=A240D;

ninexnine_unit ninexnine_unit_2768(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2041D)
);

ninexnine_unit ninexnine_unit_2769(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2141D)
);

ninexnine_unit ninexnine_unit_2770(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2241D)
);

ninexnine_unit ninexnine_unit_2771(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2341D)
);

ninexnine_unit ninexnine_unit_2772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2441D)
);

ninexnine_unit ninexnine_unit_2773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2541D)
);

ninexnine_unit ninexnine_unit_2774(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2641D)
);

ninexnine_unit ninexnine_unit_2775(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2741D)
);

assign C241D=c2041D+c2141D+c2241D+c2341D+c2441D+c2541D+c2641D+c2741D;
assign A241D=(C241D>=0)?1:0;

assign P341D=A241D;

ninexnine_unit ninexnine_unit_2776(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2042D)
);

ninexnine_unit ninexnine_unit_2777(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2142D)
);

ninexnine_unit ninexnine_unit_2778(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2242D)
);

ninexnine_unit ninexnine_unit_2779(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2342D)
);

ninexnine_unit ninexnine_unit_2780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2442D)
);

ninexnine_unit ninexnine_unit_2781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2542D)
);

ninexnine_unit ninexnine_unit_2782(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2642D)
);

ninexnine_unit ninexnine_unit_2783(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2742D)
);

assign C242D=c2042D+c2142D+c2242D+c2342D+c2442D+c2542D+c2642D+c2742D;
assign A242D=(C242D>=0)?1:0;

assign P342D=A242D;

ninexnine_unit ninexnine_unit_2784(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2043D)
);

ninexnine_unit ninexnine_unit_2785(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2143D)
);

ninexnine_unit ninexnine_unit_2786(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2243D)
);

ninexnine_unit ninexnine_unit_2787(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2343D)
);

ninexnine_unit ninexnine_unit_2788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2443D)
);

ninexnine_unit ninexnine_unit_2789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2543D)
);

ninexnine_unit ninexnine_unit_2790(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2643D)
);

ninexnine_unit ninexnine_unit_2791(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2743D)
);

assign C243D=c2043D+c2143D+c2243D+c2343D+c2443D+c2543D+c2643D+c2743D;
assign A243D=(C243D>=0)?1:0;

assign P343D=A243D;

ninexnine_unit ninexnine_unit_2792(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2044D)
);

ninexnine_unit ninexnine_unit_2793(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2144D)
);

ninexnine_unit ninexnine_unit_2794(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2244D)
);

ninexnine_unit ninexnine_unit_2795(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2344D)
);

ninexnine_unit ninexnine_unit_2796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2444D)
);

ninexnine_unit ninexnine_unit_2797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2544D)
);

ninexnine_unit ninexnine_unit_2798(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2644D)
);

ninexnine_unit ninexnine_unit_2799(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2744D)
);

assign C244D=c2044D+c2144D+c2244D+c2344D+c2444D+c2544D+c2644D+c2744D;
assign A244D=(C244D>=0)?1:0;

assign P344D=A244D;

ninexnine_unit ninexnine_unit_2800(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2000E)
);

ninexnine_unit ninexnine_unit_2801(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2100E)
);

ninexnine_unit ninexnine_unit_2802(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2200E)
);

ninexnine_unit ninexnine_unit_2803(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2300E)
);

ninexnine_unit ninexnine_unit_2804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2400E)
);

ninexnine_unit ninexnine_unit_2805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2500E)
);

ninexnine_unit ninexnine_unit_2806(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2600E)
);

ninexnine_unit ninexnine_unit_2807(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2700E)
);

assign C200E=c2000E+c2100E+c2200E+c2300E+c2400E+c2500E+c2600E+c2700E;
assign A200E=(C200E>=0)?1:0;

assign P300E=A200E;

ninexnine_unit ninexnine_unit_2808(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2001E)
);

ninexnine_unit ninexnine_unit_2809(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2101E)
);

ninexnine_unit ninexnine_unit_2810(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2201E)
);

ninexnine_unit ninexnine_unit_2811(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2301E)
);

ninexnine_unit ninexnine_unit_2812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2401E)
);

ninexnine_unit ninexnine_unit_2813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2501E)
);

ninexnine_unit ninexnine_unit_2814(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2601E)
);

ninexnine_unit ninexnine_unit_2815(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2701E)
);

assign C201E=c2001E+c2101E+c2201E+c2301E+c2401E+c2501E+c2601E+c2701E;
assign A201E=(C201E>=0)?1:0;

assign P301E=A201E;

ninexnine_unit ninexnine_unit_2816(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2002E)
);

ninexnine_unit ninexnine_unit_2817(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2102E)
);

ninexnine_unit ninexnine_unit_2818(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2202E)
);

ninexnine_unit ninexnine_unit_2819(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2302E)
);

ninexnine_unit ninexnine_unit_2820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2402E)
);

ninexnine_unit ninexnine_unit_2821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2502E)
);

ninexnine_unit ninexnine_unit_2822(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2602E)
);

ninexnine_unit ninexnine_unit_2823(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2702E)
);

assign C202E=c2002E+c2102E+c2202E+c2302E+c2402E+c2502E+c2602E+c2702E;
assign A202E=(C202E>=0)?1:0;

assign P302E=A202E;

ninexnine_unit ninexnine_unit_2824(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2003E)
);

ninexnine_unit ninexnine_unit_2825(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2103E)
);

ninexnine_unit ninexnine_unit_2826(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2203E)
);

ninexnine_unit ninexnine_unit_2827(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2303E)
);

ninexnine_unit ninexnine_unit_2828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2403E)
);

ninexnine_unit ninexnine_unit_2829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2503E)
);

ninexnine_unit ninexnine_unit_2830(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2603E)
);

ninexnine_unit ninexnine_unit_2831(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2703E)
);

assign C203E=c2003E+c2103E+c2203E+c2303E+c2403E+c2503E+c2603E+c2703E;
assign A203E=(C203E>=0)?1:0;

assign P303E=A203E;

ninexnine_unit ninexnine_unit_2832(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2004E)
);

ninexnine_unit ninexnine_unit_2833(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2104E)
);

ninexnine_unit ninexnine_unit_2834(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2204E)
);

ninexnine_unit ninexnine_unit_2835(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2304E)
);

ninexnine_unit ninexnine_unit_2836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2404E)
);

ninexnine_unit ninexnine_unit_2837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2504E)
);

ninexnine_unit ninexnine_unit_2838(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2604E)
);

ninexnine_unit ninexnine_unit_2839(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2704E)
);

assign C204E=c2004E+c2104E+c2204E+c2304E+c2404E+c2504E+c2604E+c2704E;
assign A204E=(C204E>=0)?1:0;

assign P304E=A204E;

ninexnine_unit ninexnine_unit_2840(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2010E)
);

ninexnine_unit ninexnine_unit_2841(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2110E)
);

ninexnine_unit ninexnine_unit_2842(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2210E)
);

ninexnine_unit ninexnine_unit_2843(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2310E)
);

ninexnine_unit ninexnine_unit_2844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2410E)
);

ninexnine_unit ninexnine_unit_2845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2510E)
);

ninexnine_unit ninexnine_unit_2846(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2610E)
);

ninexnine_unit ninexnine_unit_2847(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2710E)
);

assign C210E=c2010E+c2110E+c2210E+c2310E+c2410E+c2510E+c2610E+c2710E;
assign A210E=(C210E>=0)?1:0;

assign P310E=A210E;

ninexnine_unit ninexnine_unit_2848(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2011E)
);

ninexnine_unit ninexnine_unit_2849(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2111E)
);

ninexnine_unit ninexnine_unit_2850(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2211E)
);

ninexnine_unit ninexnine_unit_2851(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2311E)
);

ninexnine_unit ninexnine_unit_2852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2411E)
);

ninexnine_unit ninexnine_unit_2853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2511E)
);

ninexnine_unit ninexnine_unit_2854(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2611E)
);

ninexnine_unit ninexnine_unit_2855(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2711E)
);

assign C211E=c2011E+c2111E+c2211E+c2311E+c2411E+c2511E+c2611E+c2711E;
assign A211E=(C211E>=0)?1:0;

assign P311E=A211E;

ninexnine_unit ninexnine_unit_2856(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2012E)
);

ninexnine_unit ninexnine_unit_2857(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2112E)
);

ninexnine_unit ninexnine_unit_2858(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2212E)
);

ninexnine_unit ninexnine_unit_2859(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2312E)
);

ninexnine_unit ninexnine_unit_2860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2412E)
);

ninexnine_unit ninexnine_unit_2861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2512E)
);

ninexnine_unit ninexnine_unit_2862(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2612E)
);

ninexnine_unit ninexnine_unit_2863(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2712E)
);

assign C212E=c2012E+c2112E+c2212E+c2312E+c2412E+c2512E+c2612E+c2712E;
assign A212E=(C212E>=0)?1:0;

assign P312E=A212E;

ninexnine_unit ninexnine_unit_2864(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2013E)
);

ninexnine_unit ninexnine_unit_2865(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2113E)
);

ninexnine_unit ninexnine_unit_2866(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2213E)
);

ninexnine_unit ninexnine_unit_2867(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2313E)
);

ninexnine_unit ninexnine_unit_2868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2413E)
);

ninexnine_unit ninexnine_unit_2869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2513E)
);

ninexnine_unit ninexnine_unit_2870(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2613E)
);

ninexnine_unit ninexnine_unit_2871(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2713E)
);

assign C213E=c2013E+c2113E+c2213E+c2313E+c2413E+c2513E+c2613E+c2713E;
assign A213E=(C213E>=0)?1:0;

assign P313E=A213E;

ninexnine_unit ninexnine_unit_2872(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2014E)
);

ninexnine_unit ninexnine_unit_2873(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2114E)
);

ninexnine_unit ninexnine_unit_2874(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2214E)
);

ninexnine_unit ninexnine_unit_2875(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2314E)
);

ninexnine_unit ninexnine_unit_2876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2414E)
);

ninexnine_unit ninexnine_unit_2877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2514E)
);

ninexnine_unit ninexnine_unit_2878(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2614E)
);

ninexnine_unit ninexnine_unit_2879(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2714E)
);

assign C214E=c2014E+c2114E+c2214E+c2314E+c2414E+c2514E+c2614E+c2714E;
assign A214E=(C214E>=0)?1:0;

assign P314E=A214E;

ninexnine_unit ninexnine_unit_2880(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2020E)
);

ninexnine_unit ninexnine_unit_2881(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2120E)
);

ninexnine_unit ninexnine_unit_2882(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2220E)
);

ninexnine_unit ninexnine_unit_2883(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2320E)
);

ninexnine_unit ninexnine_unit_2884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2420E)
);

ninexnine_unit ninexnine_unit_2885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2520E)
);

ninexnine_unit ninexnine_unit_2886(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2620E)
);

ninexnine_unit ninexnine_unit_2887(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2720E)
);

assign C220E=c2020E+c2120E+c2220E+c2320E+c2420E+c2520E+c2620E+c2720E;
assign A220E=(C220E>=0)?1:0;

assign P320E=A220E;

ninexnine_unit ninexnine_unit_2888(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2021E)
);

ninexnine_unit ninexnine_unit_2889(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2121E)
);

ninexnine_unit ninexnine_unit_2890(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2221E)
);

ninexnine_unit ninexnine_unit_2891(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2321E)
);

ninexnine_unit ninexnine_unit_2892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2421E)
);

ninexnine_unit ninexnine_unit_2893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2521E)
);

ninexnine_unit ninexnine_unit_2894(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2621E)
);

ninexnine_unit ninexnine_unit_2895(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2721E)
);

assign C221E=c2021E+c2121E+c2221E+c2321E+c2421E+c2521E+c2621E+c2721E;
assign A221E=(C221E>=0)?1:0;

assign P321E=A221E;

ninexnine_unit ninexnine_unit_2896(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2022E)
);

ninexnine_unit ninexnine_unit_2897(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2122E)
);

ninexnine_unit ninexnine_unit_2898(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2222E)
);

ninexnine_unit ninexnine_unit_2899(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2322E)
);

ninexnine_unit ninexnine_unit_2900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2422E)
);

ninexnine_unit ninexnine_unit_2901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2522E)
);

ninexnine_unit ninexnine_unit_2902(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2622E)
);

ninexnine_unit ninexnine_unit_2903(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2722E)
);

assign C222E=c2022E+c2122E+c2222E+c2322E+c2422E+c2522E+c2622E+c2722E;
assign A222E=(C222E>=0)?1:0;

assign P322E=A222E;

ninexnine_unit ninexnine_unit_2904(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2023E)
);

ninexnine_unit ninexnine_unit_2905(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2123E)
);

ninexnine_unit ninexnine_unit_2906(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2223E)
);

ninexnine_unit ninexnine_unit_2907(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2323E)
);

ninexnine_unit ninexnine_unit_2908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2423E)
);

ninexnine_unit ninexnine_unit_2909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2523E)
);

ninexnine_unit ninexnine_unit_2910(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2623E)
);

ninexnine_unit ninexnine_unit_2911(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2723E)
);

assign C223E=c2023E+c2123E+c2223E+c2323E+c2423E+c2523E+c2623E+c2723E;
assign A223E=(C223E>=0)?1:0;

assign P323E=A223E;

ninexnine_unit ninexnine_unit_2912(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2024E)
);

ninexnine_unit ninexnine_unit_2913(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2124E)
);

ninexnine_unit ninexnine_unit_2914(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2224E)
);

ninexnine_unit ninexnine_unit_2915(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2324E)
);

ninexnine_unit ninexnine_unit_2916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2424E)
);

ninexnine_unit ninexnine_unit_2917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2524E)
);

ninexnine_unit ninexnine_unit_2918(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2624E)
);

ninexnine_unit ninexnine_unit_2919(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2724E)
);

assign C224E=c2024E+c2124E+c2224E+c2324E+c2424E+c2524E+c2624E+c2724E;
assign A224E=(C224E>=0)?1:0;

assign P324E=A224E;

ninexnine_unit ninexnine_unit_2920(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2030E)
);

ninexnine_unit ninexnine_unit_2921(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2130E)
);

ninexnine_unit ninexnine_unit_2922(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2230E)
);

ninexnine_unit ninexnine_unit_2923(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2330E)
);

ninexnine_unit ninexnine_unit_2924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2430E)
);

ninexnine_unit ninexnine_unit_2925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2530E)
);

ninexnine_unit ninexnine_unit_2926(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2630E)
);

ninexnine_unit ninexnine_unit_2927(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2730E)
);

assign C230E=c2030E+c2130E+c2230E+c2330E+c2430E+c2530E+c2630E+c2730E;
assign A230E=(C230E>=0)?1:0;

assign P330E=A230E;

ninexnine_unit ninexnine_unit_2928(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2031E)
);

ninexnine_unit ninexnine_unit_2929(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2131E)
);

ninexnine_unit ninexnine_unit_2930(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2231E)
);

ninexnine_unit ninexnine_unit_2931(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2331E)
);

ninexnine_unit ninexnine_unit_2932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2431E)
);

ninexnine_unit ninexnine_unit_2933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2531E)
);

ninexnine_unit ninexnine_unit_2934(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2631E)
);

ninexnine_unit ninexnine_unit_2935(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2731E)
);

assign C231E=c2031E+c2131E+c2231E+c2331E+c2431E+c2531E+c2631E+c2731E;
assign A231E=(C231E>=0)?1:0;

assign P331E=A231E;

ninexnine_unit ninexnine_unit_2936(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2032E)
);

ninexnine_unit ninexnine_unit_2937(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2132E)
);

ninexnine_unit ninexnine_unit_2938(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2232E)
);

ninexnine_unit ninexnine_unit_2939(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2332E)
);

ninexnine_unit ninexnine_unit_2940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2432E)
);

ninexnine_unit ninexnine_unit_2941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2532E)
);

ninexnine_unit ninexnine_unit_2942(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2632E)
);

ninexnine_unit ninexnine_unit_2943(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2732E)
);

assign C232E=c2032E+c2132E+c2232E+c2332E+c2432E+c2532E+c2632E+c2732E;
assign A232E=(C232E>=0)?1:0;

assign P332E=A232E;

ninexnine_unit ninexnine_unit_2944(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2033E)
);

ninexnine_unit ninexnine_unit_2945(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2133E)
);

ninexnine_unit ninexnine_unit_2946(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2233E)
);

ninexnine_unit ninexnine_unit_2947(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2333E)
);

ninexnine_unit ninexnine_unit_2948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2433E)
);

ninexnine_unit ninexnine_unit_2949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2533E)
);

ninexnine_unit ninexnine_unit_2950(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2633E)
);

ninexnine_unit ninexnine_unit_2951(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2733E)
);

assign C233E=c2033E+c2133E+c2233E+c2333E+c2433E+c2533E+c2633E+c2733E;
assign A233E=(C233E>=0)?1:0;

assign P333E=A233E;

ninexnine_unit ninexnine_unit_2952(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2034E)
);

ninexnine_unit ninexnine_unit_2953(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2134E)
);

ninexnine_unit ninexnine_unit_2954(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2234E)
);

ninexnine_unit ninexnine_unit_2955(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2334E)
);

ninexnine_unit ninexnine_unit_2956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2434E)
);

ninexnine_unit ninexnine_unit_2957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2534E)
);

ninexnine_unit ninexnine_unit_2958(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2634E)
);

ninexnine_unit ninexnine_unit_2959(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2734E)
);

assign C234E=c2034E+c2134E+c2234E+c2334E+c2434E+c2534E+c2634E+c2734E;
assign A234E=(C234E>=0)?1:0;

assign P334E=A234E;

ninexnine_unit ninexnine_unit_2960(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2040E)
);

ninexnine_unit ninexnine_unit_2961(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2140E)
);

ninexnine_unit ninexnine_unit_2962(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2240E)
);

ninexnine_unit ninexnine_unit_2963(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2340E)
);

ninexnine_unit ninexnine_unit_2964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2440E)
);

ninexnine_unit ninexnine_unit_2965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2540E)
);

ninexnine_unit ninexnine_unit_2966(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2640E)
);

ninexnine_unit ninexnine_unit_2967(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2740E)
);

assign C240E=c2040E+c2140E+c2240E+c2340E+c2440E+c2540E+c2640E+c2740E;
assign A240E=(C240E>=0)?1:0;

assign P340E=A240E;

ninexnine_unit ninexnine_unit_2968(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2041E)
);

ninexnine_unit ninexnine_unit_2969(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2141E)
);

ninexnine_unit ninexnine_unit_2970(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2241E)
);

ninexnine_unit ninexnine_unit_2971(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2341E)
);

ninexnine_unit ninexnine_unit_2972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2441E)
);

ninexnine_unit ninexnine_unit_2973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2541E)
);

ninexnine_unit ninexnine_unit_2974(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2641E)
);

ninexnine_unit ninexnine_unit_2975(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2741E)
);

assign C241E=c2041E+c2141E+c2241E+c2341E+c2441E+c2541E+c2641E+c2741E;
assign A241E=(C241E>=0)?1:0;

assign P341E=A241E;

ninexnine_unit ninexnine_unit_2976(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2042E)
);

ninexnine_unit ninexnine_unit_2977(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2142E)
);

ninexnine_unit ninexnine_unit_2978(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2242E)
);

ninexnine_unit ninexnine_unit_2979(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2342E)
);

ninexnine_unit ninexnine_unit_2980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2442E)
);

ninexnine_unit ninexnine_unit_2981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2542E)
);

ninexnine_unit ninexnine_unit_2982(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2642E)
);

ninexnine_unit ninexnine_unit_2983(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2742E)
);

assign C242E=c2042E+c2142E+c2242E+c2342E+c2442E+c2542E+c2642E+c2742E;
assign A242E=(C242E>=0)?1:0;

assign P342E=A242E;

ninexnine_unit ninexnine_unit_2984(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2043E)
);

ninexnine_unit ninexnine_unit_2985(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2143E)
);

ninexnine_unit ninexnine_unit_2986(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2243E)
);

ninexnine_unit ninexnine_unit_2987(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2343E)
);

ninexnine_unit ninexnine_unit_2988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2443E)
);

ninexnine_unit ninexnine_unit_2989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2543E)
);

ninexnine_unit ninexnine_unit_2990(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2643E)
);

ninexnine_unit ninexnine_unit_2991(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2743E)
);

assign C243E=c2043E+c2143E+c2243E+c2343E+c2443E+c2543E+c2643E+c2743E;
assign A243E=(C243E>=0)?1:0;

assign P343E=A243E;

ninexnine_unit ninexnine_unit_2992(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2044E)
);

ninexnine_unit ninexnine_unit_2993(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2144E)
);

ninexnine_unit ninexnine_unit_2994(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2244E)
);

ninexnine_unit ninexnine_unit_2995(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2344E)
);

ninexnine_unit ninexnine_unit_2996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2444E)
);

ninexnine_unit ninexnine_unit_2997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2544E)
);

ninexnine_unit ninexnine_unit_2998(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2644E)
);

ninexnine_unit ninexnine_unit_2999(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2744E)
);

assign C244E=c2044E+c2144E+c2244E+c2344E+c2444E+c2544E+c2644E+c2744E;
assign A244E=(C244E>=0)?1:0;

assign P344E=A244E;

ninexnine_unit ninexnine_unit_3000(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2000F)
);

ninexnine_unit ninexnine_unit_3001(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2100F)
);

ninexnine_unit ninexnine_unit_3002(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2200F)
);

ninexnine_unit ninexnine_unit_3003(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2300F)
);

ninexnine_unit ninexnine_unit_3004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2400F)
);

ninexnine_unit ninexnine_unit_3005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2500F)
);

ninexnine_unit ninexnine_unit_3006(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2600F)
);

ninexnine_unit ninexnine_unit_3007(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2700F)
);

assign C200F=c2000F+c2100F+c2200F+c2300F+c2400F+c2500F+c2600F+c2700F;
assign A200F=(C200F>=0)?1:0;

assign P300F=A200F;

ninexnine_unit ninexnine_unit_3008(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2001F)
);

ninexnine_unit ninexnine_unit_3009(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2101F)
);

ninexnine_unit ninexnine_unit_3010(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2201F)
);

ninexnine_unit ninexnine_unit_3011(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2301F)
);

ninexnine_unit ninexnine_unit_3012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2401F)
);

ninexnine_unit ninexnine_unit_3013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2501F)
);

ninexnine_unit ninexnine_unit_3014(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2601F)
);

ninexnine_unit ninexnine_unit_3015(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2701F)
);

assign C201F=c2001F+c2101F+c2201F+c2301F+c2401F+c2501F+c2601F+c2701F;
assign A201F=(C201F>=0)?1:0;

assign P301F=A201F;

ninexnine_unit ninexnine_unit_3016(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2002F)
);

ninexnine_unit ninexnine_unit_3017(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2102F)
);

ninexnine_unit ninexnine_unit_3018(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2202F)
);

ninexnine_unit ninexnine_unit_3019(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2302F)
);

ninexnine_unit ninexnine_unit_3020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2402F)
);

ninexnine_unit ninexnine_unit_3021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2502F)
);

ninexnine_unit ninexnine_unit_3022(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2602F)
);

ninexnine_unit ninexnine_unit_3023(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2702F)
);

assign C202F=c2002F+c2102F+c2202F+c2302F+c2402F+c2502F+c2602F+c2702F;
assign A202F=(C202F>=0)?1:0;

assign P302F=A202F;

ninexnine_unit ninexnine_unit_3024(
				.clk(clk),
				.rstn(rstn),
				.a0(P2030),
				.a1(P2040),
				.a2(P2050),
				.a3(P2130),
				.a4(P2140),
				.a5(P2150),
				.a6(P2230),
				.a7(P2240),
				.a8(P2250),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2003F)
);

ninexnine_unit ninexnine_unit_3025(
				.clk(clk),
				.rstn(rstn),
				.a0(P2031),
				.a1(P2041),
				.a2(P2051),
				.a3(P2131),
				.a4(P2141),
				.a5(P2151),
				.a6(P2231),
				.a7(P2241),
				.a8(P2251),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2103F)
);

ninexnine_unit ninexnine_unit_3026(
				.clk(clk),
				.rstn(rstn),
				.a0(P2032),
				.a1(P2042),
				.a2(P2052),
				.a3(P2132),
				.a4(P2142),
				.a5(P2152),
				.a6(P2232),
				.a7(P2242),
				.a8(P2252),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2203F)
);

ninexnine_unit ninexnine_unit_3027(
				.clk(clk),
				.rstn(rstn),
				.a0(P2033),
				.a1(P2043),
				.a2(P2053),
				.a3(P2133),
				.a4(P2143),
				.a5(P2153),
				.a6(P2233),
				.a7(P2243),
				.a8(P2253),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2303F)
);

ninexnine_unit ninexnine_unit_3028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2034),
				.a1(P2044),
				.a2(P2054),
				.a3(P2134),
				.a4(P2144),
				.a5(P2154),
				.a6(P2234),
				.a7(P2244),
				.a8(P2254),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2403F)
);

ninexnine_unit ninexnine_unit_3029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2035),
				.a1(P2045),
				.a2(P2055),
				.a3(P2135),
				.a4(P2145),
				.a5(P2155),
				.a6(P2235),
				.a7(P2245),
				.a8(P2255),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2503F)
);

ninexnine_unit ninexnine_unit_3030(
				.clk(clk),
				.rstn(rstn),
				.a0(P2036),
				.a1(P2046),
				.a2(P2056),
				.a3(P2136),
				.a4(P2146),
				.a5(P2156),
				.a6(P2236),
				.a7(P2246),
				.a8(P2256),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2603F)
);

ninexnine_unit ninexnine_unit_3031(
				.clk(clk),
				.rstn(rstn),
				.a0(P2037),
				.a1(P2047),
				.a2(P2057),
				.a3(P2137),
				.a4(P2147),
				.a5(P2157),
				.a6(P2237),
				.a7(P2247),
				.a8(P2257),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2703F)
);

assign C203F=c2003F+c2103F+c2203F+c2303F+c2403F+c2503F+c2603F+c2703F;
assign A203F=(C203F>=0)?1:0;

assign P303F=A203F;

ninexnine_unit ninexnine_unit_3032(
				.clk(clk),
				.rstn(rstn),
				.a0(P2040),
				.a1(P2050),
				.a2(P2060),
				.a3(P2140),
				.a4(P2150),
				.a5(P2160),
				.a6(P2240),
				.a7(P2250),
				.a8(P2260),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2004F)
);

ninexnine_unit ninexnine_unit_3033(
				.clk(clk),
				.rstn(rstn),
				.a0(P2041),
				.a1(P2051),
				.a2(P2061),
				.a3(P2141),
				.a4(P2151),
				.a5(P2161),
				.a6(P2241),
				.a7(P2251),
				.a8(P2261),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2104F)
);

ninexnine_unit ninexnine_unit_3034(
				.clk(clk),
				.rstn(rstn),
				.a0(P2042),
				.a1(P2052),
				.a2(P2062),
				.a3(P2142),
				.a4(P2152),
				.a5(P2162),
				.a6(P2242),
				.a7(P2252),
				.a8(P2262),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2204F)
);

ninexnine_unit ninexnine_unit_3035(
				.clk(clk),
				.rstn(rstn),
				.a0(P2043),
				.a1(P2053),
				.a2(P2063),
				.a3(P2143),
				.a4(P2153),
				.a5(P2163),
				.a6(P2243),
				.a7(P2253),
				.a8(P2263),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2304F)
);

ninexnine_unit ninexnine_unit_3036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2044),
				.a1(P2054),
				.a2(P2064),
				.a3(P2144),
				.a4(P2154),
				.a5(P2164),
				.a6(P2244),
				.a7(P2254),
				.a8(P2264),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2404F)
);

ninexnine_unit ninexnine_unit_3037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2045),
				.a1(P2055),
				.a2(P2065),
				.a3(P2145),
				.a4(P2155),
				.a5(P2165),
				.a6(P2245),
				.a7(P2255),
				.a8(P2265),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2504F)
);

ninexnine_unit ninexnine_unit_3038(
				.clk(clk),
				.rstn(rstn),
				.a0(P2046),
				.a1(P2056),
				.a2(P2066),
				.a3(P2146),
				.a4(P2156),
				.a5(P2166),
				.a6(P2246),
				.a7(P2256),
				.a8(P2266),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2604F)
);

ninexnine_unit ninexnine_unit_3039(
				.clk(clk),
				.rstn(rstn),
				.a0(P2047),
				.a1(P2057),
				.a2(P2067),
				.a3(P2147),
				.a4(P2157),
				.a5(P2167),
				.a6(P2247),
				.a7(P2257),
				.a8(P2267),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2704F)
);

assign C204F=c2004F+c2104F+c2204F+c2304F+c2404F+c2504F+c2604F+c2704F;
assign A204F=(C204F>=0)?1:0;

assign P304F=A204F;

ninexnine_unit ninexnine_unit_3040(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2010F)
);

ninexnine_unit ninexnine_unit_3041(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2110F)
);

ninexnine_unit ninexnine_unit_3042(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2210F)
);

ninexnine_unit ninexnine_unit_3043(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2310F)
);

ninexnine_unit ninexnine_unit_3044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2410F)
);

ninexnine_unit ninexnine_unit_3045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2510F)
);

ninexnine_unit ninexnine_unit_3046(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2610F)
);

ninexnine_unit ninexnine_unit_3047(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2710F)
);

assign C210F=c2010F+c2110F+c2210F+c2310F+c2410F+c2510F+c2610F+c2710F;
assign A210F=(C210F>=0)?1:0;

assign P310F=A210F;

ninexnine_unit ninexnine_unit_3048(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2011F)
);

ninexnine_unit ninexnine_unit_3049(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2111F)
);

ninexnine_unit ninexnine_unit_3050(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2211F)
);

ninexnine_unit ninexnine_unit_3051(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2311F)
);

ninexnine_unit ninexnine_unit_3052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2411F)
);

ninexnine_unit ninexnine_unit_3053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2511F)
);

ninexnine_unit ninexnine_unit_3054(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2611F)
);

ninexnine_unit ninexnine_unit_3055(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2711F)
);

assign C211F=c2011F+c2111F+c2211F+c2311F+c2411F+c2511F+c2611F+c2711F;
assign A211F=(C211F>=0)?1:0;

assign P311F=A211F;

ninexnine_unit ninexnine_unit_3056(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2012F)
);

ninexnine_unit ninexnine_unit_3057(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2112F)
);

ninexnine_unit ninexnine_unit_3058(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2212F)
);

ninexnine_unit ninexnine_unit_3059(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2312F)
);

ninexnine_unit ninexnine_unit_3060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2412F)
);

ninexnine_unit ninexnine_unit_3061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2512F)
);

ninexnine_unit ninexnine_unit_3062(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2612F)
);

ninexnine_unit ninexnine_unit_3063(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2712F)
);

assign C212F=c2012F+c2112F+c2212F+c2312F+c2412F+c2512F+c2612F+c2712F;
assign A212F=(C212F>=0)?1:0;

assign P312F=A212F;

ninexnine_unit ninexnine_unit_3064(
				.clk(clk),
				.rstn(rstn),
				.a0(P2130),
				.a1(P2140),
				.a2(P2150),
				.a3(P2230),
				.a4(P2240),
				.a5(P2250),
				.a6(P2330),
				.a7(P2340),
				.a8(P2350),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2013F)
);

ninexnine_unit ninexnine_unit_3065(
				.clk(clk),
				.rstn(rstn),
				.a0(P2131),
				.a1(P2141),
				.a2(P2151),
				.a3(P2231),
				.a4(P2241),
				.a5(P2251),
				.a6(P2331),
				.a7(P2341),
				.a8(P2351),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2113F)
);

ninexnine_unit ninexnine_unit_3066(
				.clk(clk),
				.rstn(rstn),
				.a0(P2132),
				.a1(P2142),
				.a2(P2152),
				.a3(P2232),
				.a4(P2242),
				.a5(P2252),
				.a6(P2332),
				.a7(P2342),
				.a8(P2352),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2213F)
);

ninexnine_unit ninexnine_unit_3067(
				.clk(clk),
				.rstn(rstn),
				.a0(P2133),
				.a1(P2143),
				.a2(P2153),
				.a3(P2233),
				.a4(P2243),
				.a5(P2253),
				.a6(P2333),
				.a7(P2343),
				.a8(P2353),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2313F)
);

ninexnine_unit ninexnine_unit_3068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2134),
				.a1(P2144),
				.a2(P2154),
				.a3(P2234),
				.a4(P2244),
				.a5(P2254),
				.a6(P2334),
				.a7(P2344),
				.a8(P2354),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2413F)
);

ninexnine_unit ninexnine_unit_3069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2135),
				.a1(P2145),
				.a2(P2155),
				.a3(P2235),
				.a4(P2245),
				.a5(P2255),
				.a6(P2335),
				.a7(P2345),
				.a8(P2355),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2513F)
);

ninexnine_unit ninexnine_unit_3070(
				.clk(clk),
				.rstn(rstn),
				.a0(P2136),
				.a1(P2146),
				.a2(P2156),
				.a3(P2236),
				.a4(P2246),
				.a5(P2256),
				.a6(P2336),
				.a7(P2346),
				.a8(P2356),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2613F)
);

ninexnine_unit ninexnine_unit_3071(
				.clk(clk),
				.rstn(rstn),
				.a0(P2137),
				.a1(P2147),
				.a2(P2157),
				.a3(P2237),
				.a4(P2247),
				.a5(P2257),
				.a6(P2337),
				.a7(P2347),
				.a8(P2357),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2713F)
);

assign C213F=c2013F+c2113F+c2213F+c2313F+c2413F+c2513F+c2613F+c2713F;
assign A213F=(C213F>=0)?1:0;

assign P313F=A213F;

ninexnine_unit ninexnine_unit_3072(
				.clk(clk),
				.rstn(rstn),
				.a0(P2140),
				.a1(P2150),
				.a2(P2160),
				.a3(P2240),
				.a4(P2250),
				.a5(P2260),
				.a6(P2340),
				.a7(P2350),
				.a8(P2360),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2014F)
);

ninexnine_unit ninexnine_unit_3073(
				.clk(clk),
				.rstn(rstn),
				.a0(P2141),
				.a1(P2151),
				.a2(P2161),
				.a3(P2241),
				.a4(P2251),
				.a5(P2261),
				.a6(P2341),
				.a7(P2351),
				.a8(P2361),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2114F)
);

ninexnine_unit ninexnine_unit_3074(
				.clk(clk),
				.rstn(rstn),
				.a0(P2142),
				.a1(P2152),
				.a2(P2162),
				.a3(P2242),
				.a4(P2252),
				.a5(P2262),
				.a6(P2342),
				.a7(P2352),
				.a8(P2362),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2214F)
);

ninexnine_unit ninexnine_unit_3075(
				.clk(clk),
				.rstn(rstn),
				.a0(P2143),
				.a1(P2153),
				.a2(P2163),
				.a3(P2243),
				.a4(P2253),
				.a5(P2263),
				.a6(P2343),
				.a7(P2353),
				.a8(P2363),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2314F)
);

ninexnine_unit ninexnine_unit_3076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2144),
				.a1(P2154),
				.a2(P2164),
				.a3(P2244),
				.a4(P2254),
				.a5(P2264),
				.a6(P2344),
				.a7(P2354),
				.a8(P2364),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2414F)
);

ninexnine_unit ninexnine_unit_3077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2145),
				.a1(P2155),
				.a2(P2165),
				.a3(P2245),
				.a4(P2255),
				.a5(P2265),
				.a6(P2345),
				.a7(P2355),
				.a8(P2365),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2514F)
);

ninexnine_unit ninexnine_unit_3078(
				.clk(clk),
				.rstn(rstn),
				.a0(P2146),
				.a1(P2156),
				.a2(P2166),
				.a3(P2246),
				.a4(P2256),
				.a5(P2266),
				.a6(P2346),
				.a7(P2356),
				.a8(P2366),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2614F)
);

ninexnine_unit ninexnine_unit_3079(
				.clk(clk),
				.rstn(rstn),
				.a0(P2147),
				.a1(P2157),
				.a2(P2167),
				.a3(P2247),
				.a4(P2257),
				.a5(P2267),
				.a6(P2347),
				.a7(P2357),
				.a8(P2367),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2714F)
);

assign C214F=c2014F+c2114F+c2214F+c2314F+c2414F+c2514F+c2614F+c2714F;
assign A214F=(C214F>=0)?1:0;

assign P314F=A214F;

ninexnine_unit ninexnine_unit_3080(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2020F)
);

ninexnine_unit ninexnine_unit_3081(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2120F)
);

ninexnine_unit ninexnine_unit_3082(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2220F)
);

ninexnine_unit ninexnine_unit_3083(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2320F)
);

ninexnine_unit ninexnine_unit_3084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2420F)
);

ninexnine_unit ninexnine_unit_3085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2520F)
);

ninexnine_unit ninexnine_unit_3086(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2620F)
);

ninexnine_unit ninexnine_unit_3087(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2720F)
);

assign C220F=c2020F+c2120F+c2220F+c2320F+c2420F+c2520F+c2620F+c2720F;
assign A220F=(C220F>=0)?1:0;

assign P320F=A220F;

ninexnine_unit ninexnine_unit_3088(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2021F)
);

ninexnine_unit ninexnine_unit_3089(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2121F)
);

ninexnine_unit ninexnine_unit_3090(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2221F)
);

ninexnine_unit ninexnine_unit_3091(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2321F)
);

ninexnine_unit ninexnine_unit_3092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2421F)
);

ninexnine_unit ninexnine_unit_3093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2521F)
);

ninexnine_unit ninexnine_unit_3094(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2621F)
);

ninexnine_unit ninexnine_unit_3095(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2721F)
);

assign C221F=c2021F+c2121F+c2221F+c2321F+c2421F+c2521F+c2621F+c2721F;
assign A221F=(C221F>=0)?1:0;

assign P321F=A221F;

ninexnine_unit ninexnine_unit_3096(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2022F)
);

ninexnine_unit ninexnine_unit_3097(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2122F)
);

ninexnine_unit ninexnine_unit_3098(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2222F)
);

ninexnine_unit ninexnine_unit_3099(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2322F)
);

ninexnine_unit ninexnine_unit_3100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2422F)
);

ninexnine_unit ninexnine_unit_3101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2522F)
);

ninexnine_unit ninexnine_unit_3102(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2622F)
);

ninexnine_unit ninexnine_unit_3103(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2722F)
);

assign C222F=c2022F+c2122F+c2222F+c2322F+c2422F+c2522F+c2622F+c2722F;
assign A222F=(C222F>=0)?1:0;

assign P322F=A222F;

ninexnine_unit ninexnine_unit_3104(
				.clk(clk),
				.rstn(rstn),
				.a0(P2230),
				.a1(P2240),
				.a2(P2250),
				.a3(P2330),
				.a4(P2340),
				.a5(P2350),
				.a6(P2430),
				.a7(P2440),
				.a8(P2450),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2023F)
);

ninexnine_unit ninexnine_unit_3105(
				.clk(clk),
				.rstn(rstn),
				.a0(P2231),
				.a1(P2241),
				.a2(P2251),
				.a3(P2331),
				.a4(P2341),
				.a5(P2351),
				.a6(P2431),
				.a7(P2441),
				.a8(P2451),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2123F)
);

ninexnine_unit ninexnine_unit_3106(
				.clk(clk),
				.rstn(rstn),
				.a0(P2232),
				.a1(P2242),
				.a2(P2252),
				.a3(P2332),
				.a4(P2342),
				.a5(P2352),
				.a6(P2432),
				.a7(P2442),
				.a8(P2452),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2223F)
);

ninexnine_unit ninexnine_unit_3107(
				.clk(clk),
				.rstn(rstn),
				.a0(P2233),
				.a1(P2243),
				.a2(P2253),
				.a3(P2333),
				.a4(P2343),
				.a5(P2353),
				.a6(P2433),
				.a7(P2443),
				.a8(P2453),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2323F)
);

ninexnine_unit ninexnine_unit_3108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2234),
				.a1(P2244),
				.a2(P2254),
				.a3(P2334),
				.a4(P2344),
				.a5(P2354),
				.a6(P2434),
				.a7(P2444),
				.a8(P2454),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2423F)
);

ninexnine_unit ninexnine_unit_3109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2235),
				.a1(P2245),
				.a2(P2255),
				.a3(P2335),
				.a4(P2345),
				.a5(P2355),
				.a6(P2435),
				.a7(P2445),
				.a8(P2455),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2523F)
);

ninexnine_unit ninexnine_unit_3110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2236),
				.a1(P2246),
				.a2(P2256),
				.a3(P2336),
				.a4(P2346),
				.a5(P2356),
				.a6(P2436),
				.a7(P2446),
				.a8(P2456),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2623F)
);

ninexnine_unit ninexnine_unit_3111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2237),
				.a1(P2247),
				.a2(P2257),
				.a3(P2337),
				.a4(P2347),
				.a5(P2357),
				.a6(P2437),
				.a7(P2447),
				.a8(P2457),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2723F)
);

assign C223F=c2023F+c2123F+c2223F+c2323F+c2423F+c2523F+c2623F+c2723F;
assign A223F=(C223F>=0)?1:0;

assign P323F=A223F;

ninexnine_unit ninexnine_unit_3112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2240),
				.a1(P2250),
				.a2(P2260),
				.a3(P2340),
				.a4(P2350),
				.a5(P2360),
				.a6(P2440),
				.a7(P2450),
				.a8(P2460),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2024F)
);

ninexnine_unit ninexnine_unit_3113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2241),
				.a1(P2251),
				.a2(P2261),
				.a3(P2341),
				.a4(P2351),
				.a5(P2361),
				.a6(P2441),
				.a7(P2451),
				.a8(P2461),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2124F)
);

ninexnine_unit ninexnine_unit_3114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2242),
				.a1(P2252),
				.a2(P2262),
				.a3(P2342),
				.a4(P2352),
				.a5(P2362),
				.a6(P2442),
				.a7(P2452),
				.a8(P2462),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2224F)
);

ninexnine_unit ninexnine_unit_3115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2243),
				.a1(P2253),
				.a2(P2263),
				.a3(P2343),
				.a4(P2353),
				.a5(P2363),
				.a6(P2443),
				.a7(P2453),
				.a8(P2463),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2324F)
);

ninexnine_unit ninexnine_unit_3116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2244),
				.a1(P2254),
				.a2(P2264),
				.a3(P2344),
				.a4(P2354),
				.a5(P2364),
				.a6(P2444),
				.a7(P2454),
				.a8(P2464),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2424F)
);

ninexnine_unit ninexnine_unit_3117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2245),
				.a1(P2255),
				.a2(P2265),
				.a3(P2345),
				.a4(P2355),
				.a5(P2365),
				.a6(P2445),
				.a7(P2455),
				.a8(P2465),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2524F)
);

ninexnine_unit ninexnine_unit_3118(
				.clk(clk),
				.rstn(rstn),
				.a0(P2246),
				.a1(P2256),
				.a2(P2266),
				.a3(P2346),
				.a4(P2356),
				.a5(P2366),
				.a6(P2446),
				.a7(P2456),
				.a8(P2466),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2624F)
);

ninexnine_unit ninexnine_unit_3119(
				.clk(clk),
				.rstn(rstn),
				.a0(P2247),
				.a1(P2257),
				.a2(P2267),
				.a3(P2347),
				.a4(P2357),
				.a5(P2367),
				.a6(P2447),
				.a7(P2457),
				.a8(P2467),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2724F)
);

assign C224F=c2024F+c2124F+c2224F+c2324F+c2424F+c2524F+c2624F+c2724F;
assign A224F=(C224F>=0)?1:0;

assign P324F=A224F;

ninexnine_unit ninexnine_unit_3120(
				.clk(clk),
				.rstn(rstn),
				.a0(P2300),
				.a1(P2310),
				.a2(P2320),
				.a3(P2400),
				.a4(P2410),
				.a5(P2420),
				.a6(P2500),
				.a7(P2510),
				.a8(P2520),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2030F)
);

ninexnine_unit ninexnine_unit_3121(
				.clk(clk),
				.rstn(rstn),
				.a0(P2301),
				.a1(P2311),
				.a2(P2321),
				.a3(P2401),
				.a4(P2411),
				.a5(P2421),
				.a6(P2501),
				.a7(P2511),
				.a8(P2521),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2130F)
);

ninexnine_unit ninexnine_unit_3122(
				.clk(clk),
				.rstn(rstn),
				.a0(P2302),
				.a1(P2312),
				.a2(P2322),
				.a3(P2402),
				.a4(P2412),
				.a5(P2422),
				.a6(P2502),
				.a7(P2512),
				.a8(P2522),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2230F)
);

ninexnine_unit ninexnine_unit_3123(
				.clk(clk),
				.rstn(rstn),
				.a0(P2303),
				.a1(P2313),
				.a2(P2323),
				.a3(P2403),
				.a4(P2413),
				.a5(P2423),
				.a6(P2503),
				.a7(P2513),
				.a8(P2523),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2330F)
);

ninexnine_unit ninexnine_unit_3124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2304),
				.a1(P2314),
				.a2(P2324),
				.a3(P2404),
				.a4(P2414),
				.a5(P2424),
				.a6(P2504),
				.a7(P2514),
				.a8(P2524),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2430F)
);

ninexnine_unit ninexnine_unit_3125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2305),
				.a1(P2315),
				.a2(P2325),
				.a3(P2405),
				.a4(P2415),
				.a5(P2425),
				.a6(P2505),
				.a7(P2515),
				.a8(P2525),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2530F)
);

ninexnine_unit ninexnine_unit_3126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2306),
				.a1(P2316),
				.a2(P2326),
				.a3(P2406),
				.a4(P2416),
				.a5(P2426),
				.a6(P2506),
				.a7(P2516),
				.a8(P2526),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2630F)
);

ninexnine_unit ninexnine_unit_3127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2307),
				.a1(P2317),
				.a2(P2327),
				.a3(P2407),
				.a4(P2417),
				.a5(P2427),
				.a6(P2507),
				.a7(P2517),
				.a8(P2527),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2730F)
);

assign C230F=c2030F+c2130F+c2230F+c2330F+c2430F+c2530F+c2630F+c2730F;
assign A230F=(C230F>=0)?1:0;

assign P330F=A230F;

ninexnine_unit ninexnine_unit_3128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2310),
				.a1(P2320),
				.a2(P2330),
				.a3(P2410),
				.a4(P2420),
				.a5(P2430),
				.a6(P2510),
				.a7(P2520),
				.a8(P2530),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2031F)
);

ninexnine_unit ninexnine_unit_3129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2311),
				.a1(P2321),
				.a2(P2331),
				.a3(P2411),
				.a4(P2421),
				.a5(P2431),
				.a6(P2511),
				.a7(P2521),
				.a8(P2531),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2131F)
);

ninexnine_unit ninexnine_unit_3130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2312),
				.a1(P2322),
				.a2(P2332),
				.a3(P2412),
				.a4(P2422),
				.a5(P2432),
				.a6(P2512),
				.a7(P2522),
				.a8(P2532),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2231F)
);

ninexnine_unit ninexnine_unit_3131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2313),
				.a1(P2323),
				.a2(P2333),
				.a3(P2413),
				.a4(P2423),
				.a5(P2433),
				.a6(P2513),
				.a7(P2523),
				.a8(P2533),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2331F)
);

ninexnine_unit ninexnine_unit_3132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2314),
				.a1(P2324),
				.a2(P2334),
				.a3(P2414),
				.a4(P2424),
				.a5(P2434),
				.a6(P2514),
				.a7(P2524),
				.a8(P2534),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2431F)
);

ninexnine_unit ninexnine_unit_3133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2315),
				.a1(P2325),
				.a2(P2335),
				.a3(P2415),
				.a4(P2425),
				.a5(P2435),
				.a6(P2515),
				.a7(P2525),
				.a8(P2535),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2531F)
);

ninexnine_unit ninexnine_unit_3134(
				.clk(clk),
				.rstn(rstn),
				.a0(P2316),
				.a1(P2326),
				.a2(P2336),
				.a3(P2416),
				.a4(P2426),
				.a5(P2436),
				.a6(P2516),
				.a7(P2526),
				.a8(P2536),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2631F)
);

ninexnine_unit ninexnine_unit_3135(
				.clk(clk),
				.rstn(rstn),
				.a0(P2317),
				.a1(P2327),
				.a2(P2337),
				.a3(P2417),
				.a4(P2427),
				.a5(P2437),
				.a6(P2517),
				.a7(P2527),
				.a8(P2537),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2731F)
);

assign C231F=c2031F+c2131F+c2231F+c2331F+c2431F+c2531F+c2631F+c2731F;
assign A231F=(C231F>=0)?1:0;

assign P331F=A231F;

ninexnine_unit ninexnine_unit_3136(
				.clk(clk),
				.rstn(rstn),
				.a0(P2320),
				.a1(P2330),
				.a2(P2340),
				.a3(P2420),
				.a4(P2430),
				.a5(P2440),
				.a6(P2520),
				.a7(P2530),
				.a8(P2540),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2032F)
);

ninexnine_unit ninexnine_unit_3137(
				.clk(clk),
				.rstn(rstn),
				.a0(P2321),
				.a1(P2331),
				.a2(P2341),
				.a3(P2421),
				.a4(P2431),
				.a5(P2441),
				.a6(P2521),
				.a7(P2531),
				.a8(P2541),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2132F)
);

ninexnine_unit ninexnine_unit_3138(
				.clk(clk),
				.rstn(rstn),
				.a0(P2322),
				.a1(P2332),
				.a2(P2342),
				.a3(P2422),
				.a4(P2432),
				.a5(P2442),
				.a6(P2522),
				.a7(P2532),
				.a8(P2542),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2232F)
);

ninexnine_unit ninexnine_unit_3139(
				.clk(clk),
				.rstn(rstn),
				.a0(P2323),
				.a1(P2333),
				.a2(P2343),
				.a3(P2423),
				.a4(P2433),
				.a5(P2443),
				.a6(P2523),
				.a7(P2533),
				.a8(P2543),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2332F)
);

ninexnine_unit ninexnine_unit_3140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2324),
				.a1(P2334),
				.a2(P2344),
				.a3(P2424),
				.a4(P2434),
				.a5(P2444),
				.a6(P2524),
				.a7(P2534),
				.a8(P2544),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2432F)
);

ninexnine_unit ninexnine_unit_3141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2325),
				.a1(P2335),
				.a2(P2345),
				.a3(P2425),
				.a4(P2435),
				.a5(P2445),
				.a6(P2525),
				.a7(P2535),
				.a8(P2545),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2532F)
);

ninexnine_unit ninexnine_unit_3142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2326),
				.a1(P2336),
				.a2(P2346),
				.a3(P2426),
				.a4(P2436),
				.a5(P2446),
				.a6(P2526),
				.a7(P2536),
				.a8(P2546),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2632F)
);

ninexnine_unit ninexnine_unit_3143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2327),
				.a1(P2337),
				.a2(P2347),
				.a3(P2427),
				.a4(P2437),
				.a5(P2447),
				.a6(P2527),
				.a7(P2537),
				.a8(P2547),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2732F)
);

assign C232F=c2032F+c2132F+c2232F+c2332F+c2432F+c2532F+c2632F+c2732F;
assign A232F=(C232F>=0)?1:0;

assign P332F=A232F;

ninexnine_unit ninexnine_unit_3144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2330),
				.a1(P2340),
				.a2(P2350),
				.a3(P2430),
				.a4(P2440),
				.a5(P2450),
				.a6(P2530),
				.a7(P2540),
				.a8(P2550),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2033F)
);

ninexnine_unit ninexnine_unit_3145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2331),
				.a1(P2341),
				.a2(P2351),
				.a3(P2431),
				.a4(P2441),
				.a5(P2451),
				.a6(P2531),
				.a7(P2541),
				.a8(P2551),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2133F)
);

ninexnine_unit ninexnine_unit_3146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2332),
				.a1(P2342),
				.a2(P2352),
				.a3(P2432),
				.a4(P2442),
				.a5(P2452),
				.a6(P2532),
				.a7(P2542),
				.a8(P2552),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2233F)
);

ninexnine_unit ninexnine_unit_3147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2333),
				.a1(P2343),
				.a2(P2353),
				.a3(P2433),
				.a4(P2443),
				.a5(P2453),
				.a6(P2533),
				.a7(P2543),
				.a8(P2553),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2333F)
);

ninexnine_unit ninexnine_unit_3148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2334),
				.a1(P2344),
				.a2(P2354),
				.a3(P2434),
				.a4(P2444),
				.a5(P2454),
				.a6(P2534),
				.a7(P2544),
				.a8(P2554),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2433F)
);

ninexnine_unit ninexnine_unit_3149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2335),
				.a1(P2345),
				.a2(P2355),
				.a3(P2435),
				.a4(P2445),
				.a5(P2455),
				.a6(P2535),
				.a7(P2545),
				.a8(P2555),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2533F)
);

ninexnine_unit ninexnine_unit_3150(
				.clk(clk),
				.rstn(rstn),
				.a0(P2336),
				.a1(P2346),
				.a2(P2356),
				.a3(P2436),
				.a4(P2446),
				.a5(P2456),
				.a6(P2536),
				.a7(P2546),
				.a8(P2556),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2633F)
);

ninexnine_unit ninexnine_unit_3151(
				.clk(clk),
				.rstn(rstn),
				.a0(P2337),
				.a1(P2347),
				.a2(P2357),
				.a3(P2437),
				.a4(P2447),
				.a5(P2457),
				.a6(P2537),
				.a7(P2547),
				.a8(P2557),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2733F)
);

assign C233F=c2033F+c2133F+c2233F+c2333F+c2433F+c2533F+c2633F+c2733F;
assign A233F=(C233F>=0)?1:0;

assign P333F=A233F;

ninexnine_unit ninexnine_unit_3152(
				.clk(clk),
				.rstn(rstn),
				.a0(P2340),
				.a1(P2350),
				.a2(P2360),
				.a3(P2440),
				.a4(P2450),
				.a5(P2460),
				.a6(P2540),
				.a7(P2550),
				.a8(P2560),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2034F)
);

ninexnine_unit ninexnine_unit_3153(
				.clk(clk),
				.rstn(rstn),
				.a0(P2341),
				.a1(P2351),
				.a2(P2361),
				.a3(P2441),
				.a4(P2451),
				.a5(P2461),
				.a6(P2541),
				.a7(P2551),
				.a8(P2561),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2134F)
);

ninexnine_unit ninexnine_unit_3154(
				.clk(clk),
				.rstn(rstn),
				.a0(P2342),
				.a1(P2352),
				.a2(P2362),
				.a3(P2442),
				.a4(P2452),
				.a5(P2462),
				.a6(P2542),
				.a7(P2552),
				.a8(P2562),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2234F)
);

ninexnine_unit ninexnine_unit_3155(
				.clk(clk),
				.rstn(rstn),
				.a0(P2343),
				.a1(P2353),
				.a2(P2363),
				.a3(P2443),
				.a4(P2453),
				.a5(P2463),
				.a6(P2543),
				.a7(P2553),
				.a8(P2563),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2334F)
);

ninexnine_unit ninexnine_unit_3156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2344),
				.a1(P2354),
				.a2(P2364),
				.a3(P2444),
				.a4(P2454),
				.a5(P2464),
				.a6(P2544),
				.a7(P2554),
				.a8(P2564),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2434F)
);

ninexnine_unit ninexnine_unit_3157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2345),
				.a1(P2355),
				.a2(P2365),
				.a3(P2445),
				.a4(P2455),
				.a5(P2465),
				.a6(P2545),
				.a7(P2555),
				.a8(P2565),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2534F)
);

ninexnine_unit ninexnine_unit_3158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2346),
				.a1(P2356),
				.a2(P2366),
				.a3(P2446),
				.a4(P2456),
				.a5(P2466),
				.a6(P2546),
				.a7(P2556),
				.a8(P2566),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2634F)
);

ninexnine_unit ninexnine_unit_3159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2347),
				.a1(P2357),
				.a2(P2367),
				.a3(P2447),
				.a4(P2457),
				.a5(P2467),
				.a6(P2547),
				.a7(P2557),
				.a8(P2567),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2734F)
);

assign C234F=c2034F+c2134F+c2234F+c2334F+c2434F+c2534F+c2634F+c2734F;
assign A234F=(C234F>=0)?1:0;

assign P334F=A234F;

ninexnine_unit ninexnine_unit_3160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2400),
				.a1(P2410),
				.a2(P2420),
				.a3(P2500),
				.a4(P2510),
				.a5(P2520),
				.a6(P2600),
				.a7(P2610),
				.a8(P2620),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2040F)
);

ninexnine_unit ninexnine_unit_3161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2401),
				.a1(P2411),
				.a2(P2421),
				.a3(P2501),
				.a4(P2511),
				.a5(P2521),
				.a6(P2601),
				.a7(P2611),
				.a8(P2621),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2140F)
);

ninexnine_unit ninexnine_unit_3162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2402),
				.a1(P2412),
				.a2(P2422),
				.a3(P2502),
				.a4(P2512),
				.a5(P2522),
				.a6(P2602),
				.a7(P2612),
				.a8(P2622),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2240F)
);

ninexnine_unit ninexnine_unit_3163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2403),
				.a1(P2413),
				.a2(P2423),
				.a3(P2503),
				.a4(P2513),
				.a5(P2523),
				.a6(P2603),
				.a7(P2613),
				.a8(P2623),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2340F)
);

ninexnine_unit ninexnine_unit_3164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2404),
				.a1(P2414),
				.a2(P2424),
				.a3(P2504),
				.a4(P2514),
				.a5(P2524),
				.a6(P2604),
				.a7(P2614),
				.a8(P2624),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2440F)
);

ninexnine_unit ninexnine_unit_3165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2405),
				.a1(P2415),
				.a2(P2425),
				.a3(P2505),
				.a4(P2515),
				.a5(P2525),
				.a6(P2605),
				.a7(P2615),
				.a8(P2625),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2540F)
);

ninexnine_unit ninexnine_unit_3166(
				.clk(clk),
				.rstn(rstn),
				.a0(P2406),
				.a1(P2416),
				.a2(P2426),
				.a3(P2506),
				.a4(P2516),
				.a5(P2526),
				.a6(P2606),
				.a7(P2616),
				.a8(P2626),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2640F)
);

ninexnine_unit ninexnine_unit_3167(
				.clk(clk),
				.rstn(rstn),
				.a0(P2407),
				.a1(P2417),
				.a2(P2427),
				.a3(P2507),
				.a4(P2517),
				.a5(P2527),
				.a6(P2607),
				.a7(P2617),
				.a8(P2627),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2740F)
);

assign C240F=c2040F+c2140F+c2240F+c2340F+c2440F+c2540F+c2640F+c2740F;
assign A240F=(C240F>=0)?1:0;

assign P340F=A240F;

ninexnine_unit ninexnine_unit_3168(
				.clk(clk),
				.rstn(rstn),
				.a0(P2410),
				.a1(P2420),
				.a2(P2430),
				.a3(P2510),
				.a4(P2520),
				.a5(P2530),
				.a6(P2610),
				.a7(P2620),
				.a8(P2630),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2041F)
);

ninexnine_unit ninexnine_unit_3169(
				.clk(clk),
				.rstn(rstn),
				.a0(P2411),
				.a1(P2421),
				.a2(P2431),
				.a3(P2511),
				.a4(P2521),
				.a5(P2531),
				.a6(P2611),
				.a7(P2621),
				.a8(P2631),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2141F)
);

ninexnine_unit ninexnine_unit_3170(
				.clk(clk),
				.rstn(rstn),
				.a0(P2412),
				.a1(P2422),
				.a2(P2432),
				.a3(P2512),
				.a4(P2522),
				.a5(P2532),
				.a6(P2612),
				.a7(P2622),
				.a8(P2632),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2241F)
);

ninexnine_unit ninexnine_unit_3171(
				.clk(clk),
				.rstn(rstn),
				.a0(P2413),
				.a1(P2423),
				.a2(P2433),
				.a3(P2513),
				.a4(P2523),
				.a5(P2533),
				.a6(P2613),
				.a7(P2623),
				.a8(P2633),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2341F)
);

ninexnine_unit ninexnine_unit_3172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2414),
				.a1(P2424),
				.a2(P2434),
				.a3(P2514),
				.a4(P2524),
				.a5(P2534),
				.a6(P2614),
				.a7(P2624),
				.a8(P2634),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2441F)
);

ninexnine_unit ninexnine_unit_3173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2415),
				.a1(P2425),
				.a2(P2435),
				.a3(P2515),
				.a4(P2525),
				.a5(P2535),
				.a6(P2615),
				.a7(P2625),
				.a8(P2635),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2541F)
);

ninexnine_unit ninexnine_unit_3174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2416),
				.a1(P2426),
				.a2(P2436),
				.a3(P2516),
				.a4(P2526),
				.a5(P2536),
				.a6(P2616),
				.a7(P2626),
				.a8(P2636),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2641F)
);

ninexnine_unit ninexnine_unit_3175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2417),
				.a1(P2427),
				.a2(P2437),
				.a3(P2517),
				.a4(P2527),
				.a5(P2537),
				.a6(P2617),
				.a7(P2627),
				.a8(P2637),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2741F)
);

assign C241F=c2041F+c2141F+c2241F+c2341F+c2441F+c2541F+c2641F+c2741F;
assign A241F=(C241F>=0)?1:0;

assign P341F=A241F;

ninexnine_unit ninexnine_unit_3176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2420),
				.a1(P2430),
				.a2(P2440),
				.a3(P2520),
				.a4(P2530),
				.a5(P2540),
				.a6(P2620),
				.a7(P2630),
				.a8(P2640),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2042F)
);

ninexnine_unit ninexnine_unit_3177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2421),
				.a1(P2431),
				.a2(P2441),
				.a3(P2521),
				.a4(P2531),
				.a5(P2541),
				.a6(P2621),
				.a7(P2631),
				.a8(P2641),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2142F)
);

ninexnine_unit ninexnine_unit_3178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2422),
				.a1(P2432),
				.a2(P2442),
				.a3(P2522),
				.a4(P2532),
				.a5(P2542),
				.a6(P2622),
				.a7(P2632),
				.a8(P2642),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2242F)
);

ninexnine_unit ninexnine_unit_3179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2423),
				.a1(P2433),
				.a2(P2443),
				.a3(P2523),
				.a4(P2533),
				.a5(P2543),
				.a6(P2623),
				.a7(P2633),
				.a8(P2643),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2342F)
);

ninexnine_unit ninexnine_unit_3180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2424),
				.a1(P2434),
				.a2(P2444),
				.a3(P2524),
				.a4(P2534),
				.a5(P2544),
				.a6(P2624),
				.a7(P2634),
				.a8(P2644),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2442F)
);

ninexnine_unit ninexnine_unit_3181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2425),
				.a1(P2435),
				.a2(P2445),
				.a3(P2525),
				.a4(P2535),
				.a5(P2545),
				.a6(P2625),
				.a7(P2635),
				.a8(P2645),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2542F)
);

ninexnine_unit ninexnine_unit_3182(
				.clk(clk),
				.rstn(rstn),
				.a0(P2426),
				.a1(P2436),
				.a2(P2446),
				.a3(P2526),
				.a4(P2536),
				.a5(P2546),
				.a6(P2626),
				.a7(P2636),
				.a8(P2646),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2642F)
);

ninexnine_unit ninexnine_unit_3183(
				.clk(clk),
				.rstn(rstn),
				.a0(P2427),
				.a1(P2437),
				.a2(P2447),
				.a3(P2527),
				.a4(P2537),
				.a5(P2547),
				.a6(P2627),
				.a7(P2637),
				.a8(P2647),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2742F)
);

assign C242F=c2042F+c2142F+c2242F+c2342F+c2442F+c2542F+c2642F+c2742F;
assign A242F=(C242F>=0)?1:0;

assign P342F=A242F;

ninexnine_unit ninexnine_unit_3184(
				.clk(clk),
				.rstn(rstn),
				.a0(P2430),
				.a1(P2440),
				.a2(P2450),
				.a3(P2530),
				.a4(P2540),
				.a5(P2550),
				.a6(P2630),
				.a7(P2640),
				.a8(P2650),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2043F)
);

ninexnine_unit ninexnine_unit_3185(
				.clk(clk),
				.rstn(rstn),
				.a0(P2431),
				.a1(P2441),
				.a2(P2451),
				.a3(P2531),
				.a4(P2541),
				.a5(P2551),
				.a6(P2631),
				.a7(P2641),
				.a8(P2651),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2143F)
);

ninexnine_unit ninexnine_unit_3186(
				.clk(clk),
				.rstn(rstn),
				.a0(P2432),
				.a1(P2442),
				.a2(P2452),
				.a3(P2532),
				.a4(P2542),
				.a5(P2552),
				.a6(P2632),
				.a7(P2642),
				.a8(P2652),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2243F)
);

ninexnine_unit ninexnine_unit_3187(
				.clk(clk),
				.rstn(rstn),
				.a0(P2433),
				.a1(P2443),
				.a2(P2453),
				.a3(P2533),
				.a4(P2543),
				.a5(P2553),
				.a6(P2633),
				.a7(P2643),
				.a8(P2653),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2343F)
);

ninexnine_unit ninexnine_unit_3188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2434),
				.a1(P2444),
				.a2(P2454),
				.a3(P2534),
				.a4(P2544),
				.a5(P2554),
				.a6(P2634),
				.a7(P2644),
				.a8(P2654),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2443F)
);

ninexnine_unit ninexnine_unit_3189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2435),
				.a1(P2445),
				.a2(P2455),
				.a3(P2535),
				.a4(P2545),
				.a5(P2555),
				.a6(P2635),
				.a7(P2645),
				.a8(P2655),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2543F)
);

ninexnine_unit ninexnine_unit_3190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2436),
				.a1(P2446),
				.a2(P2456),
				.a3(P2536),
				.a4(P2546),
				.a5(P2556),
				.a6(P2636),
				.a7(P2646),
				.a8(P2656),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2643F)
);

ninexnine_unit ninexnine_unit_3191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2437),
				.a1(P2447),
				.a2(P2457),
				.a3(P2537),
				.a4(P2547),
				.a5(P2557),
				.a6(P2637),
				.a7(P2647),
				.a8(P2657),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2743F)
);

assign C243F=c2043F+c2143F+c2243F+c2343F+c2443F+c2543F+c2643F+c2743F;
assign A243F=(C243F>=0)?1:0;

assign P343F=A243F;

ninexnine_unit ninexnine_unit_3192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2440),
				.a1(P2450),
				.a2(P2460),
				.a3(P2540),
				.a4(P2550),
				.a5(P2560),
				.a6(P2640),
				.a7(P2650),
				.a8(P2660),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2044F)
);

ninexnine_unit ninexnine_unit_3193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2441),
				.a1(P2451),
				.a2(P2461),
				.a3(P2541),
				.a4(P2551),
				.a5(P2561),
				.a6(P2641),
				.a7(P2651),
				.a8(P2661),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2144F)
);

ninexnine_unit ninexnine_unit_3194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2442),
				.a1(P2452),
				.a2(P2462),
				.a3(P2542),
				.a4(P2552),
				.a5(P2562),
				.a6(P2642),
				.a7(P2652),
				.a8(P2662),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2244F)
);

ninexnine_unit ninexnine_unit_3195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2443),
				.a1(P2453),
				.a2(P2463),
				.a3(P2543),
				.a4(P2553),
				.a5(P2563),
				.a6(P2643),
				.a7(P2653),
				.a8(P2663),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2344F)
);

ninexnine_unit ninexnine_unit_3196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2444),
				.a1(P2454),
				.a2(P2464),
				.a3(P2544),
				.a4(P2554),
				.a5(P2564),
				.a6(P2644),
				.a7(P2654),
				.a8(P2664),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2444F)
);

ninexnine_unit ninexnine_unit_3197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2445),
				.a1(P2455),
				.a2(P2465),
				.a3(P2545),
				.a4(P2555),
				.a5(P2565),
				.a6(P2645),
				.a7(P2655),
				.a8(P2665),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2544F)
);

ninexnine_unit ninexnine_unit_3198(
				.clk(clk),
				.rstn(rstn),
				.a0(P2446),
				.a1(P2456),
				.a2(P2466),
				.a3(P2546),
				.a4(P2556),
				.a5(P2566),
				.a6(P2646),
				.a7(P2656),
				.a8(P2666),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2644F)
);

ninexnine_unit ninexnine_unit_3199(
				.clk(clk),
				.rstn(rstn),
				.a0(P2447),
				.a1(P2457),
				.a2(P2467),
				.a3(P2547),
				.a4(P2557),
				.a5(P2567),
				.a6(P2647),
				.a7(P2657),
				.a8(P2667),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2744F)
);

assign C244F=c2044F+c2144F+c2244F+c2344F+c2444F+c2544F+c2644F+c2744F;
assign A244F=(C244F>=0)?1:0;

assign P344F=A244F;

//layer2 done, begain next layer
(*DONT_TOUCH="true"*) wire P4000;
(*DONT_TOUCH="true"*) wire P4010;
(*DONT_TOUCH="true"*) wire P4020;
(*DONT_TOUCH="true"*) wire P4100;
(*DONT_TOUCH="true"*) wire P4110;
(*DONT_TOUCH="true"*) wire P4120;
(*DONT_TOUCH="true"*) wire P4200;
(*DONT_TOUCH="true"*) wire P4210;
(*DONT_TOUCH="true"*) wire P4220;
(*DONT_TOUCH="true"*) wire P4001;
(*DONT_TOUCH="true"*) wire P4011;
(*DONT_TOUCH="true"*) wire P4021;
(*DONT_TOUCH="true"*) wire P4101;
(*DONT_TOUCH="true"*) wire P4111;
(*DONT_TOUCH="true"*) wire P4121;
(*DONT_TOUCH="true"*) wire P4201;
(*DONT_TOUCH="true"*) wire P4211;
(*DONT_TOUCH="true"*) wire P4221;
(*DONT_TOUCH="true"*) wire P4002;
(*DONT_TOUCH="true"*) wire P4012;
(*DONT_TOUCH="true"*) wire P4022;
(*DONT_TOUCH="true"*) wire P4102;
(*DONT_TOUCH="true"*) wire P4112;
(*DONT_TOUCH="true"*) wire P4122;
(*DONT_TOUCH="true"*) wire P4202;
(*DONT_TOUCH="true"*) wire P4212;
(*DONT_TOUCH="true"*) wire P4222;
(*DONT_TOUCH="true"*) wire P4003;
(*DONT_TOUCH="true"*) wire P4013;
(*DONT_TOUCH="true"*) wire P4023;
(*DONT_TOUCH="true"*) wire P4103;
(*DONT_TOUCH="true"*) wire P4113;
(*DONT_TOUCH="true"*) wire P4123;
(*DONT_TOUCH="true"*) wire P4203;
(*DONT_TOUCH="true"*) wire P4213;
(*DONT_TOUCH="true"*) wire P4223;
(*DONT_TOUCH="true"*) wire P4004;
(*DONT_TOUCH="true"*) wire P4014;
(*DONT_TOUCH="true"*) wire P4024;
(*DONT_TOUCH="true"*) wire P4104;
(*DONT_TOUCH="true"*) wire P4114;
(*DONT_TOUCH="true"*) wire P4124;
(*DONT_TOUCH="true"*) wire P4204;
(*DONT_TOUCH="true"*) wire P4214;
(*DONT_TOUCH="true"*) wire P4224;
(*DONT_TOUCH="true"*) wire P4005;
(*DONT_TOUCH="true"*) wire P4015;
(*DONT_TOUCH="true"*) wire P4025;
(*DONT_TOUCH="true"*) wire P4105;
(*DONT_TOUCH="true"*) wire P4115;
(*DONT_TOUCH="true"*) wire P4125;
(*DONT_TOUCH="true"*) wire P4205;
(*DONT_TOUCH="true"*) wire P4215;
(*DONT_TOUCH="true"*) wire P4225;
(*DONT_TOUCH="true"*) wire P4006;
(*DONT_TOUCH="true"*) wire P4016;
(*DONT_TOUCH="true"*) wire P4026;
(*DONT_TOUCH="true"*) wire P4106;
(*DONT_TOUCH="true"*) wire P4116;
(*DONT_TOUCH="true"*) wire P4126;
(*DONT_TOUCH="true"*) wire P4206;
(*DONT_TOUCH="true"*) wire P4216;
(*DONT_TOUCH="true"*) wire P4226;
(*DONT_TOUCH="true"*) wire P4007;
(*DONT_TOUCH="true"*) wire P4017;
(*DONT_TOUCH="true"*) wire P4027;
(*DONT_TOUCH="true"*) wire P4107;
(*DONT_TOUCH="true"*) wire P4117;
(*DONT_TOUCH="true"*) wire P4127;
(*DONT_TOUCH="true"*) wire P4207;
(*DONT_TOUCH="true"*) wire P4217;
(*DONT_TOUCH="true"*) wire P4227;
(*DONT_TOUCH="true"*) wire P4008;
(*DONT_TOUCH="true"*) wire P4018;
(*DONT_TOUCH="true"*) wire P4028;
(*DONT_TOUCH="true"*) wire P4108;
(*DONT_TOUCH="true"*) wire P4118;
(*DONT_TOUCH="true"*) wire P4128;
(*DONT_TOUCH="true"*) wire P4208;
(*DONT_TOUCH="true"*) wire P4218;
(*DONT_TOUCH="true"*) wire P4228;
(*DONT_TOUCH="true"*) wire P4009;
(*DONT_TOUCH="true"*) wire P4019;
(*DONT_TOUCH="true"*) wire P4029;
(*DONT_TOUCH="true"*) wire P4109;
(*DONT_TOUCH="true"*) wire P4119;
(*DONT_TOUCH="true"*) wire P4129;
(*DONT_TOUCH="true"*) wire P4209;
(*DONT_TOUCH="true"*) wire P4219;
(*DONT_TOUCH="true"*) wire P4229;
(*DONT_TOUCH="true"*) wire P400A;
(*DONT_TOUCH="true"*) wire P401A;
(*DONT_TOUCH="true"*) wire P402A;
(*DONT_TOUCH="true"*) wire P410A;
(*DONT_TOUCH="true"*) wire P411A;
(*DONT_TOUCH="true"*) wire P412A;
(*DONT_TOUCH="true"*) wire P420A;
(*DONT_TOUCH="true"*) wire P421A;
(*DONT_TOUCH="true"*) wire P422A;
(*DONT_TOUCH="true"*) wire P400B;
(*DONT_TOUCH="true"*) wire P401B;
(*DONT_TOUCH="true"*) wire P402B;
(*DONT_TOUCH="true"*) wire P410B;
(*DONT_TOUCH="true"*) wire P411B;
(*DONT_TOUCH="true"*) wire P412B;
(*DONT_TOUCH="true"*) wire P420B;
(*DONT_TOUCH="true"*) wire P421B;
(*DONT_TOUCH="true"*) wire P422B;
(*DONT_TOUCH="true"*) wire P400C;
(*DONT_TOUCH="true"*) wire P401C;
(*DONT_TOUCH="true"*) wire P402C;
(*DONT_TOUCH="true"*) wire P410C;
(*DONT_TOUCH="true"*) wire P411C;
(*DONT_TOUCH="true"*) wire P412C;
(*DONT_TOUCH="true"*) wire P420C;
(*DONT_TOUCH="true"*) wire P421C;
(*DONT_TOUCH="true"*) wire P422C;
(*DONT_TOUCH="true"*) wire P400D;
(*DONT_TOUCH="true"*) wire P401D;
(*DONT_TOUCH="true"*) wire P402D;
(*DONT_TOUCH="true"*) wire P410D;
(*DONT_TOUCH="true"*) wire P411D;
(*DONT_TOUCH="true"*) wire P412D;
(*DONT_TOUCH="true"*) wire P420D;
(*DONT_TOUCH="true"*) wire P421D;
(*DONT_TOUCH="true"*) wire P422D;
(*DONT_TOUCH="true"*) wire P400E;
(*DONT_TOUCH="true"*) wire P401E;
(*DONT_TOUCH="true"*) wire P402E;
(*DONT_TOUCH="true"*) wire P410E;
(*DONT_TOUCH="true"*) wire P411E;
(*DONT_TOUCH="true"*) wire P412E;
(*DONT_TOUCH="true"*) wire P420E;
(*DONT_TOUCH="true"*) wire P421E;
(*DONT_TOUCH="true"*) wire P422E;
(*DONT_TOUCH="true"*) wire P400F;
(*DONT_TOUCH="true"*) wire P401F;
(*DONT_TOUCH="true"*) wire P402F;
(*DONT_TOUCH="true"*) wire P410F;
(*DONT_TOUCH="true"*) wire P411F;
(*DONT_TOUCH="true"*) wire P412F;
(*DONT_TOUCH="true"*) wire P420F;
(*DONT_TOUCH="true"*) wire P421F;
(*DONT_TOUCH="true"*) wire P422F;
(*DONT_TOUCH="true"*) wire P400G;
(*DONT_TOUCH="true"*) wire P401G;
(*DONT_TOUCH="true"*) wire P402G;
(*DONT_TOUCH="true"*) wire P410G;
(*DONT_TOUCH="true"*) wire P411G;
(*DONT_TOUCH="true"*) wire P412G;
(*DONT_TOUCH="true"*) wire P420G;
(*DONT_TOUCH="true"*) wire P421G;
(*DONT_TOUCH="true"*) wire P422G;
(*DONT_TOUCH="true"*) wire P400H;
(*DONT_TOUCH="true"*) wire P401H;
(*DONT_TOUCH="true"*) wire P402H;
(*DONT_TOUCH="true"*) wire P410H;
(*DONT_TOUCH="true"*) wire P411H;
(*DONT_TOUCH="true"*) wire P412H;
(*DONT_TOUCH="true"*) wire P420H;
(*DONT_TOUCH="true"*) wire P421H;
(*DONT_TOUCH="true"*) wire P422H;
(*DONT_TOUCH="true"*) wire P400I;
(*DONT_TOUCH="true"*) wire P401I;
(*DONT_TOUCH="true"*) wire P402I;
(*DONT_TOUCH="true"*) wire P410I;
(*DONT_TOUCH="true"*) wire P411I;
(*DONT_TOUCH="true"*) wire P412I;
(*DONT_TOUCH="true"*) wire P420I;
(*DONT_TOUCH="true"*) wire P421I;
(*DONT_TOUCH="true"*) wire P422I;
(*DONT_TOUCH="true"*) wire P400J;
(*DONT_TOUCH="true"*) wire P401J;
(*DONT_TOUCH="true"*) wire P402J;
(*DONT_TOUCH="true"*) wire P410J;
(*DONT_TOUCH="true"*) wire P411J;
(*DONT_TOUCH="true"*) wire P412J;
(*DONT_TOUCH="true"*) wire P420J;
(*DONT_TOUCH="true"*) wire P421J;
(*DONT_TOUCH="true"*) wire P422J;
(*DONT_TOUCH="true"*) wire P400K;
(*DONT_TOUCH="true"*) wire P401K;
(*DONT_TOUCH="true"*) wire P402K;
(*DONT_TOUCH="true"*) wire P410K;
(*DONT_TOUCH="true"*) wire P411K;
(*DONT_TOUCH="true"*) wire P412K;
(*DONT_TOUCH="true"*) wire P420K;
(*DONT_TOUCH="true"*) wire P421K;
(*DONT_TOUCH="true"*) wire P422K;
(*DONT_TOUCH="true"*) wire P400L;
(*DONT_TOUCH="true"*) wire P401L;
(*DONT_TOUCH="true"*) wire P402L;
(*DONT_TOUCH="true"*) wire P410L;
(*DONT_TOUCH="true"*) wire P411L;
(*DONT_TOUCH="true"*) wire P412L;
(*DONT_TOUCH="true"*) wire P420L;
(*DONT_TOUCH="true"*) wire P421L;
(*DONT_TOUCH="true"*) wire P422L;
(*DONT_TOUCH="true"*) wire P400M;
(*DONT_TOUCH="true"*) wire P401M;
(*DONT_TOUCH="true"*) wire P402M;
(*DONT_TOUCH="true"*) wire P410M;
(*DONT_TOUCH="true"*) wire P411M;
(*DONT_TOUCH="true"*) wire P412M;
(*DONT_TOUCH="true"*) wire P420M;
(*DONT_TOUCH="true"*) wire P421M;
(*DONT_TOUCH="true"*) wire P422M;
(*DONT_TOUCH="true"*) wire P400N;
(*DONT_TOUCH="true"*) wire P401N;
(*DONT_TOUCH="true"*) wire P402N;
(*DONT_TOUCH="true"*) wire P410N;
(*DONT_TOUCH="true"*) wire P411N;
(*DONT_TOUCH="true"*) wire P412N;
(*DONT_TOUCH="true"*) wire P420N;
(*DONT_TOUCH="true"*) wire P421N;
(*DONT_TOUCH="true"*) wire P422N;
(*DONT_TOUCH="true"*) wire P400O;
(*DONT_TOUCH="true"*) wire P401O;
(*DONT_TOUCH="true"*) wire P402O;
(*DONT_TOUCH="true"*) wire P410O;
(*DONT_TOUCH="true"*) wire P411O;
(*DONT_TOUCH="true"*) wire P412O;
(*DONT_TOUCH="true"*) wire P420O;
(*DONT_TOUCH="true"*) wire P421O;
(*DONT_TOUCH="true"*) wire P422O;
(*DONT_TOUCH="true"*) wire P400P;
(*DONT_TOUCH="true"*) wire P401P;
(*DONT_TOUCH="true"*) wire P402P;
(*DONT_TOUCH="true"*) wire P410P;
(*DONT_TOUCH="true"*) wire P411P;
(*DONT_TOUCH="true"*) wire P412P;
(*DONT_TOUCH="true"*) wire P420P;
(*DONT_TOUCH="true"*) wire P421P;
(*DONT_TOUCH="true"*) wire P422P;
(*DONT_TOUCH="true"*) wire P400Q;
(*DONT_TOUCH="true"*) wire P401Q;
(*DONT_TOUCH="true"*) wire P402Q;
(*DONT_TOUCH="true"*) wire P410Q;
(*DONT_TOUCH="true"*) wire P411Q;
(*DONT_TOUCH="true"*) wire P412Q;
(*DONT_TOUCH="true"*) wire P420Q;
(*DONT_TOUCH="true"*) wire P421Q;
(*DONT_TOUCH="true"*) wire P422Q;
(*DONT_TOUCH="true"*) wire P400R;
(*DONT_TOUCH="true"*) wire P401R;
(*DONT_TOUCH="true"*) wire P402R;
(*DONT_TOUCH="true"*) wire P410R;
(*DONT_TOUCH="true"*) wire P411R;
(*DONT_TOUCH="true"*) wire P412R;
(*DONT_TOUCH="true"*) wire P420R;
(*DONT_TOUCH="true"*) wire P421R;
(*DONT_TOUCH="true"*) wire P422R;
(*DONT_TOUCH="true"*) wire P400S;
(*DONT_TOUCH="true"*) wire P401S;
(*DONT_TOUCH="true"*) wire P402S;
(*DONT_TOUCH="true"*) wire P410S;
(*DONT_TOUCH="true"*) wire P411S;
(*DONT_TOUCH="true"*) wire P412S;
(*DONT_TOUCH="true"*) wire P420S;
(*DONT_TOUCH="true"*) wire P421S;
(*DONT_TOUCH="true"*) wire P422S;
(*DONT_TOUCH="true"*) wire P400T;
(*DONT_TOUCH="true"*) wire P401T;
(*DONT_TOUCH="true"*) wire P402T;
(*DONT_TOUCH="true"*) wire P410T;
(*DONT_TOUCH="true"*) wire P411T;
(*DONT_TOUCH="true"*) wire P412T;
(*DONT_TOUCH="true"*) wire P420T;
(*DONT_TOUCH="true"*) wire P421T;
(*DONT_TOUCH="true"*) wire P422T;
(*DONT_TOUCH="true"*) wire P400U;
(*DONT_TOUCH="true"*) wire P401U;
(*DONT_TOUCH="true"*) wire P402U;
(*DONT_TOUCH="true"*) wire P410U;
(*DONT_TOUCH="true"*) wire P411U;
(*DONT_TOUCH="true"*) wire P412U;
(*DONT_TOUCH="true"*) wire P420U;
(*DONT_TOUCH="true"*) wire P421U;
(*DONT_TOUCH="true"*) wire P422U;
(*DONT_TOUCH="true"*) wire P400V;
(*DONT_TOUCH="true"*) wire P401V;
(*DONT_TOUCH="true"*) wire P402V;
(*DONT_TOUCH="true"*) wire P410V;
(*DONT_TOUCH="true"*) wire P411V;
(*DONT_TOUCH="true"*) wire P412V;
(*DONT_TOUCH="true"*) wire P420V;
(*DONT_TOUCH="true"*) wire P421V;
(*DONT_TOUCH="true"*) wire P422V;
(*DONT_TOUCH="true"*) wire W30000,W30010,W30020,W30100,W30110,W30120,W30200,W30210,W30220;
(*DONT_TOUCH="true"*) wire W30001,W30011,W30021,W30101,W30111,W30121,W30201,W30211,W30221;
(*DONT_TOUCH="true"*) wire W30002,W30012,W30022,W30102,W30112,W30122,W30202,W30212,W30222;
(*DONT_TOUCH="true"*) wire W30003,W30013,W30023,W30103,W30113,W30123,W30203,W30213,W30223;
(*DONT_TOUCH="true"*) wire W30004,W30014,W30024,W30104,W30114,W30124,W30204,W30214,W30224;
(*DONT_TOUCH="true"*) wire W30005,W30015,W30025,W30105,W30115,W30125,W30205,W30215,W30225;
(*DONT_TOUCH="true"*) wire W30006,W30016,W30026,W30106,W30116,W30126,W30206,W30216,W30226;
(*DONT_TOUCH="true"*) wire W30007,W30017,W30027,W30107,W30117,W30127,W30207,W30217,W30227;
(*DONT_TOUCH="true"*) wire W30008,W30018,W30028,W30108,W30118,W30128,W30208,W30218,W30228;
(*DONT_TOUCH="true"*) wire W30009,W30019,W30029,W30109,W30119,W30129,W30209,W30219,W30229;
(*DONT_TOUCH="true"*) wire W3000A,W3001A,W3002A,W3010A,W3011A,W3012A,W3020A,W3021A,W3022A;
(*DONT_TOUCH="true"*) wire W3000B,W3001B,W3002B,W3010B,W3011B,W3012B,W3020B,W3021B,W3022B;
(*DONT_TOUCH="true"*) wire W3000C,W3001C,W3002C,W3010C,W3011C,W3012C,W3020C,W3021C,W3022C;
(*DONT_TOUCH="true"*) wire W3000D,W3001D,W3002D,W3010D,W3011D,W3012D,W3020D,W3021D,W3022D;
(*DONT_TOUCH="true"*) wire W3000E,W3001E,W3002E,W3010E,W3011E,W3012E,W3020E,W3021E,W3022E;
(*DONT_TOUCH="true"*) wire W3000F,W3001F,W3002F,W3010F,W3011F,W3012F,W3020F,W3021F,W3022F;
(*DONT_TOUCH="true"*) wire W31000,W31010,W31020,W31100,W31110,W31120,W31200,W31210,W31220;
(*DONT_TOUCH="true"*) wire W31001,W31011,W31021,W31101,W31111,W31121,W31201,W31211,W31221;
(*DONT_TOUCH="true"*) wire W31002,W31012,W31022,W31102,W31112,W31122,W31202,W31212,W31222;
(*DONT_TOUCH="true"*) wire W31003,W31013,W31023,W31103,W31113,W31123,W31203,W31213,W31223;
(*DONT_TOUCH="true"*) wire W31004,W31014,W31024,W31104,W31114,W31124,W31204,W31214,W31224;
(*DONT_TOUCH="true"*) wire W31005,W31015,W31025,W31105,W31115,W31125,W31205,W31215,W31225;
(*DONT_TOUCH="true"*) wire W31006,W31016,W31026,W31106,W31116,W31126,W31206,W31216,W31226;
(*DONT_TOUCH="true"*) wire W31007,W31017,W31027,W31107,W31117,W31127,W31207,W31217,W31227;
(*DONT_TOUCH="true"*) wire W31008,W31018,W31028,W31108,W31118,W31128,W31208,W31218,W31228;
(*DONT_TOUCH="true"*) wire W31009,W31019,W31029,W31109,W31119,W31129,W31209,W31219,W31229;
(*DONT_TOUCH="true"*) wire W3100A,W3101A,W3102A,W3110A,W3111A,W3112A,W3120A,W3121A,W3122A;
(*DONT_TOUCH="true"*) wire W3100B,W3101B,W3102B,W3110B,W3111B,W3112B,W3120B,W3121B,W3122B;
(*DONT_TOUCH="true"*) wire W3100C,W3101C,W3102C,W3110C,W3111C,W3112C,W3120C,W3121C,W3122C;
(*DONT_TOUCH="true"*) wire W3100D,W3101D,W3102D,W3110D,W3111D,W3112D,W3120D,W3121D,W3122D;
(*DONT_TOUCH="true"*) wire W3100E,W3101E,W3102E,W3110E,W3111E,W3112E,W3120E,W3121E,W3122E;
(*DONT_TOUCH="true"*) wire W3100F,W3101F,W3102F,W3110F,W3111F,W3112F,W3120F,W3121F,W3122F;
(*DONT_TOUCH="true"*) wire W32000,W32010,W32020,W32100,W32110,W32120,W32200,W32210,W32220;
(*DONT_TOUCH="true"*) wire W32001,W32011,W32021,W32101,W32111,W32121,W32201,W32211,W32221;
(*DONT_TOUCH="true"*) wire W32002,W32012,W32022,W32102,W32112,W32122,W32202,W32212,W32222;
(*DONT_TOUCH="true"*) wire W32003,W32013,W32023,W32103,W32113,W32123,W32203,W32213,W32223;
(*DONT_TOUCH="true"*) wire W32004,W32014,W32024,W32104,W32114,W32124,W32204,W32214,W32224;
(*DONT_TOUCH="true"*) wire W32005,W32015,W32025,W32105,W32115,W32125,W32205,W32215,W32225;
(*DONT_TOUCH="true"*) wire W32006,W32016,W32026,W32106,W32116,W32126,W32206,W32216,W32226;
(*DONT_TOUCH="true"*) wire W32007,W32017,W32027,W32107,W32117,W32127,W32207,W32217,W32227;
(*DONT_TOUCH="true"*) wire W32008,W32018,W32028,W32108,W32118,W32128,W32208,W32218,W32228;
(*DONT_TOUCH="true"*) wire W32009,W32019,W32029,W32109,W32119,W32129,W32209,W32219,W32229;
(*DONT_TOUCH="true"*) wire W3200A,W3201A,W3202A,W3210A,W3211A,W3212A,W3220A,W3221A,W3222A;
(*DONT_TOUCH="true"*) wire W3200B,W3201B,W3202B,W3210B,W3211B,W3212B,W3220B,W3221B,W3222B;
(*DONT_TOUCH="true"*) wire W3200C,W3201C,W3202C,W3210C,W3211C,W3212C,W3220C,W3221C,W3222C;
(*DONT_TOUCH="true"*) wire W3200D,W3201D,W3202D,W3210D,W3211D,W3212D,W3220D,W3221D,W3222D;
(*DONT_TOUCH="true"*) wire W3200E,W3201E,W3202E,W3210E,W3211E,W3212E,W3220E,W3221E,W3222E;
(*DONT_TOUCH="true"*) wire W3200F,W3201F,W3202F,W3210F,W3211F,W3212F,W3220F,W3221F,W3222F;
(*DONT_TOUCH="true"*) wire W33000,W33010,W33020,W33100,W33110,W33120,W33200,W33210,W33220;
(*DONT_TOUCH="true"*) wire W33001,W33011,W33021,W33101,W33111,W33121,W33201,W33211,W33221;
(*DONT_TOUCH="true"*) wire W33002,W33012,W33022,W33102,W33112,W33122,W33202,W33212,W33222;
(*DONT_TOUCH="true"*) wire W33003,W33013,W33023,W33103,W33113,W33123,W33203,W33213,W33223;
(*DONT_TOUCH="true"*) wire W33004,W33014,W33024,W33104,W33114,W33124,W33204,W33214,W33224;
(*DONT_TOUCH="true"*) wire W33005,W33015,W33025,W33105,W33115,W33125,W33205,W33215,W33225;
(*DONT_TOUCH="true"*) wire W33006,W33016,W33026,W33106,W33116,W33126,W33206,W33216,W33226;
(*DONT_TOUCH="true"*) wire W33007,W33017,W33027,W33107,W33117,W33127,W33207,W33217,W33227;
(*DONT_TOUCH="true"*) wire W33008,W33018,W33028,W33108,W33118,W33128,W33208,W33218,W33228;
(*DONT_TOUCH="true"*) wire W33009,W33019,W33029,W33109,W33119,W33129,W33209,W33219,W33229;
(*DONT_TOUCH="true"*) wire W3300A,W3301A,W3302A,W3310A,W3311A,W3312A,W3320A,W3321A,W3322A;
(*DONT_TOUCH="true"*) wire W3300B,W3301B,W3302B,W3310B,W3311B,W3312B,W3320B,W3321B,W3322B;
(*DONT_TOUCH="true"*) wire W3300C,W3301C,W3302C,W3310C,W3311C,W3312C,W3320C,W3321C,W3322C;
(*DONT_TOUCH="true"*) wire W3300D,W3301D,W3302D,W3310D,W3311D,W3312D,W3320D,W3321D,W3322D;
(*DONT_TOUCH="true"*) wire W3300E,W3301E,W3302E,W3310E,W3311E,W3312E,W3320E,W3321E,W3322E;
(*DONT_TOUCH="true"*) wire W3300F,W3301F,W3302F,W3310F,W3311F,W3312F,W3320F,W3321F,W3322F;
(*DONT_TOUCH="true"*) wire W34000,W34010,W34020,W34100,W34110,W34120,W34200,W34210,W34220;
(*DONT_TOUCH="true"*) wire W34001,W34011,W34021,W34101,W34111,W34121,W34201,W34211,W34221;
(*DONT_TOUCH="true"*) wire W34002,W34012,W34022,W34102,W34112,W34122,W34202,W34212,W34222;
(*DONT_TOUCH="true"*) wire W34003,W34013,W34023,W34103,W34113,W34123,W34203,W34213,W34223;
(*DONT_TOUCH="true"*) wire W34004,W34014,W34024,W34104,W34114,W34124,W34204,W34214,W34224;
(*DONT_TOUCH="true"*) wire W34005,W34015,W34025,W34105,W34115,W34125,W34205,W34215,W34225;
(*DONT_TOUCH="true"*) wire W34006,W34016,W34026,W34106,W34116,W34126,W34206,W34216,W34226;
(*DONT_TOUCH="true"*) wire W34007,W34017,W34027,W34107,W34117,W34127,W34207,W34217,W34227;
(*DONT_TOUCH="true"*) wire W34008,W34018,W34028,W34108,W34118,W34128,W34208,W34218,W34228;
(*DONT_TOUCH="true"*) wire W34009,W34019,W34029,W34109,W34119,W34129,W34209,W34219,W34229;
(*DONT_TOUCH="true"*) wire W3400A,W3401A,W3402A,W3410A,W3411A,W3412A,W3420A,W3421A,W3422A;
(*DONT_TOUCH="true"*) wire W3400B,W3401B,W3402B,W3410B,W3411B,W3412B,W3420B,W3421B,W3422B;
(*DONT_TOUCH="true"*) wire W3400C,W3401C,W3402C,W3410C,W3411C,W3412C,W3420C,W3421C,W3422C;
(*DONT_TOUCH="true"*) wire W3400D,W3401D,W3402D,W3410D,W3411D,W3412D,W3420D,W3421D,W3422D;
(*DONT_TOUCH="true"*) wire W3400E,W3401E,W3402E,W3410E,W3411E,W3412E,W3420E,W3421E,W3422E;
(*DONT_TOUCH="true"*) wire W3400F,W3401F,W3402F,W3410F,W3411F,W3412F,W3420F,W3421F,W3422F;
(*DONT_TOUCH="true"*) wire W35000,W35010,W35020,W35100,W35110,W35120,W35200,W35210,W35220;
(*DONT_TOUCH="true"*) wire W35001,W35011,W35021,W35101,W35111,W35121,W35201,W35211,W35221;
(*DONT_TOUCH="true"*) wire W35002,W35012,W35022,W35102,W35112,W35122,W35202,W35212,W35222;
(*DONT_TOUCH="true"*) wire W35003,W35013,W35023,W35103,W35113,W35123,W35203,W35213,W35223;
(*DONT_TOUCH="true"*) wire W35004,W35014,W35024,W35104,W35114,W35124,W35204,W35214,W35224;
(*DONT_TOUCH="true"*) wire W35005,W35015,W35025,W35105,W35115,W35125,W35205,W35215,W35225;
(*DONT_TOUCH="true"*) wire W35006,W35016,W35026,W35106,W35116,W35126,W35206,W35216,W35226;
(*DONT_TOUCH="true"*) wire W35007,W35017,W35027,W35107,W35117,W35127,W35207,W35217,W35227;
(*DONT_TOUCH="true"*) wire W35008,W35018,W35028,W35108,W35118,W35128,W35208,W35218,W35228;
(*DONT_TOUCH="true"*) wire W35009,W35019,W35029,W35109,W35119,W35129,W35209,W35219,W35229;
(*DONT_TOUCH="true"*) wire W3500A,W3501A,W3502A,W3510A,W3511A,W3512A,W3520A,W3521A,W3522A;
(*DONT_TOUCH="true"*) wire W3500B,W3501B,W3502B,W3510B,W3511B,W3512B,W3520B,W3521B,W3522B;
(*DONT_TOUCH="true"*) wire W3500C,W3501C,W3502C,W3510C,W3511C,W3512C,W3520C,W3521C,W3522C;
(*DONT_TOUCH="true"*) wire W3500D,W3501D,W3502D,W3510D,W3511D,W3512D,W3520D,W3521D,W3522D;
(*DONT_TOUCH="true"*) wire W3500E,W3501E,W3502E,W3510E,W3511E,W3512E,W3520E,W3521E,W3522E;
(*DONT_TOUCH="true"*) wire W3500F,W3501F,W3502F,W3510F,W3511F,W3512F,W3520F,W3521F,W3522F;
(*DONT_TOUCH="true"*) wire W36000,W36010,W36020,W36100,W36110,W36120,W36200,W36210,W36220;
(*DONT_TOUCH="true"*) wire W36001,W36011,W36021,W36101,W36111,W36121,W36201,W36211,W36221;
(*DONT_TOUCH="true"*) wire W36002,W36012,W36022,W36102,W36112,W36122,W36202,W36212,W36222;
(*DONT_TOUCH="true"*) wire W36003,W36013,W36023,W36103,W36113,W36123,W36203,W36213,W36223;
(*DONT_TOUCH="true"*) wire W36004,W36014,W36024,W36104,W36114,W36124,W36204,W36214,W36224;
(*DONT_TOUCH="true"*) wire W36005,W36015,W36025,W36105,W36115,W36125,W36205,W36215,W36225;
(*DONT_TOUCH="true"*) wire W36006,W36016,W36026,W36106,W36116,W36126,W36206,W36216,W36226;
(*DONT_TOUCH="true"*) wire W36007,W36017,W36027,W36107,W36117,W36127,W36207,W36217,W36227;
(*DONT_TOUCH="true"*) wire W36008,W36018,W36028,W36108,W36118,W36128,W36208,W36218,W36228;
(*DONT_TOUCH="true"*) wire W36009,W36019,W36029,W36109,W36119,W36129,W36209,W36219,W36229;
(*DONT_TOUCH="true"*) wire W3600A,W3601A,W3602A,W3610A,W3611A,W3612A,W3620A,W3621A,W3622A;
(*DONT_TOUCH="true"*) wire W3600B,W3601B,W3602B,W3610B,W3611B,W3612B,W3620B,W3621B,W3622B;
(*DONT_TOUCH="true"*) wire W3600C,W3601C,W3602C,W3610C,W3611C,W3612C,W3620C,W3621C,W3622C;
(*DONT_TOUCH="true"*) wire W3600D,W3601D,W3602D,W3610D,W3611D,W3612D,W3620D,W3621D,W3622D;
(*DONT_TOUCH="true"*) wire W3600E,W3601E,W3602E,W3610E,W3611E,W3612E,W3620E,W3621E,W3622E;
(*DONT_TOUCH="true"*) wire W3600F,W3601F,W3602F,W3610F,W3611F,W3612F,W3620F,W3621F,W3622F;
(*DONT_TOUCH="true"*) wire W37000,W37010,W37020,W37100,W37110,W37120,W37200,W37210,W37220;
(*DONT_TOUCH="true"*) wire W37001,W37011,W37021,W37101,W37111,W37121,W37201,W37211,W37221;
(*DONT_TOUCH="true"*) wire W37002,W37012,W37022,W37102,W37112,W37122,W37202,W37212,W37222;
(*DONT_TOUCH="true"*) wire W37003,W37013,W37023,W37103,W37113,W37123,W37203,W37213,W37223;
(*DONT_TOUCH="true"*) wire W37004,W37014,W37024,W37104,W37114,W37124,W37204,W37214,W37224;
(*DONT_TOUCH="true"*) wire W37005,W37015,W37025,W37105,W37115,W37125,W37205,W37215,W37225;
(*DONT_TOUCH="true"*) wire W37006,W37016,W37026,W37106,W37116,W37126,W37206,W37216,W37226;
(*DONT_TOUCH="true"*) wire W37007,W37017,W37027,W37107,W37117,W37127,W37207,W37217,W37227;
(*DONT_TOUCH="true"*) wire W37008,W37018,W37028,W37108,W37118,W37128,W37208,W37218,W37228;
(*DONT_TOUCH="true"*) wire W37009,W37019,W37029,W37109,W37119,W37129,W37209,W37219,W37229;
(*DONT_TOUCH="true"*) wire W3700A,W3701A,W3702A,W3710A,W3711A,W3712A,W3720A,W3721A,W3722A;
(*DONT_TOUCH="true"*) wire W3700B,W3701B,W3702B,W3710B,W3711B,W3712B,W3720B,W3721B,W3722B;
(*DONT_TOUCH="true"*) wire W3700C,W3701C,W3702C,W3710C,W3711C,W3712C,W3720C,W3721C,W3722C;
(*DONT_TOUCH="true"*) wire W3700D,W3701D,W3702D,W3710D,W3711D,W3712D,W3720D,W3721D,W3722D;
(*DONT_TOUCH="true"*) wire W3700E,W3701E,W3702E,W3710E,W3711E,W3712E,W3720E,W3721E,W3722E;
(*DONT_TOUCH="true"*) wire W3700F,W3701F,W3702F,W3710F,W3711F,W3712F,W3720F,W3721F,W3722F;
(*DONT_TOUCH="true"*) wire W38000,W38010,W38020,W38100,W38110,W38120,W38200,W38210,W38220;
(*DONT_TOUCH="true"*) wire W38001,W38011,W38021,W38101,W38111,W38121,W38201,W38211,W38221;
(*DONT_TOUCH="true"*) wire W38002,W38012,W38022,W38102,W38112,W38122,W38202,W38212,W38222;
(*DONT_TOUCH="true"*) wire W38003,W38013,W38023,W38103,W38113,W38123,W38203,W38213,W38223;
(*DONT_TOUCH="true"*) wire W38004,W38014,W38024,W38104,W38114,W38124,W38204,W38214,W38224;
(*DONT_TOUCH="true"*) wire W38005,W38015,W38025,W38105,W38115,W38125,W38205,W38215,W38225;
(*DONT_TOUCH="true"*) wire W38006,W38016,W38026,W38106,W38116,W38126,W38206,W38216,W38226;
(*DONT_TOUCH="true"*) wire W38007,W38017,W38027,W38107,W38117,W38127,W38207,W38217,W38227;
(*DONT_TOUCH="true"*) wire W38008,W38018,W38028,W38108,W38118,W38128,W38208,W38218,W38228;
(*DONT_TOUCH="true"*) wire W38009,W38019,W38029,W38109,W38119,W38129,W38209,W38219,W38229;
(*DONT_TOUCH="true"*) wire W3800A,W3801A,W3802A,W3810A,W3811A,W3812A,W3820A,W3821A,W3822A;
(*DONT_TOUCH="true"*) wire W3800B,W3801B,W3802B,W3810B,W3811B,W3812B,W3820B,W3821B,W3822B;
(*DONT_TOUCH="true"*) wire W3800C,W3801C,W3802C,W3810C,W3811C,W3812C,W3820C,W3821C,W3822C;
(*DONT_TOUCH="true"*) wire W3800D,W3801D,W3802D,W3810D,W3811D,W3812D,W3820D,W3821D,W3822D;
(*DONT_TOUCH="true"*) wire W3800E,W3801E,W3802E,W3810E,W3811E,W3812E,W3820E,W3821E,W3822E;
(*DONT_TOUCH="true"*) wire W3800F,W3801F,W3802F,W3810F,W3811F,W3812F,W3820F,W3821F,W3822F;
(*DONT_TOUCH="true"*) wire W39000,W39010,W39020,W39100,W39110,W39120,W39200,W39210,W39220;
(*DONT_TOUCH="true"*) wire W39001,W39011,W39021,W39101,W39111,W39121,W39201,W39211,W39221;
(*DONT_TOUCH="true"*) wire W39002,W39012,W39022,W39102,W39112,W39122,W39202,W39212,W39222;
(*DONT_TOUCH="true"*) wire W39003,W39013,W39023,W39103,W39113,W39123,W39203,W39213,W39223;
(*DONT_TOUCH="true"*) wire W39004,W39014,W39024,W39104,W39114,W39124,W39204,W39214,W39224;
(*DONT_TOUCH="true"*) wire W39005,W39015,W39025,W39105,W39115,W39125,W39205,W39215,W39225;
(*DONT_TOUCH="true"*) wire W39006,W39016,W39026,W39106,W39116,W39126,W39206,W39216,W39226;
(*DONT_TOUCH="true"*) wire W39007,W39017,W39027,W39107,W39117,W39127,W39207,W39217,W39227;
(*DONT_TOUCH="true"*) wire W39008,W39018,W39028,W39108,W39118,W39128,W39208,W39218,W39228;
(*DONT_TOUCH="true"*) wire W39009,W39019,W39029,W39109,W39119,W39129,W39209,W39219,W39229;
(*DONT_TOUCH="true"*) wire W3900A,W3901A,W3902A,W3910A,W3911A,W3912A,W3920A,W3921A,W3922A;
(*DONT_TOUCH="true"*) wire W3900B,W3901B,W3902B,W3910B,W3911B,W3912B,W3920B,W3921B,W3922B;
(*DONT_TOUCH="true"*) wire W3900C,W3901C,W3902C,W3910C,W3911C,W3912C,W3920C,W3921C,W3922C;
(*DONT_TOUCH="true"*) wire W3900D,W3901D,W3902D,W3910D,W3911D,W3912D,W3920D,W3921D,W3922D;
(*DONT_TOUCH="true"*) wire W3900E,W3901E,W3902E,W3910E,W3911E,W3912E,W3920E,W3921E,W3922E;
(*DONT_TOUCH="true"*) wire W3900F,W3901F,W3902F,W3910F,W3911F,W3912F,W3920F,W3921F,W3922F;
(*DONT_TOUCH="true"*) wire W3A000,W3A010,W3A020,W3A100,W3A110,W3A120,W3A200,W3A210,W3A220;
(*DONT_TOUCH="true"*) wire W3A001,W3A011,W3A021,W3A101,W3A111,W3A121,W3A201,W3A211,W3A221;
(*DONT_TOUCH="true"*) wire W3A002,W3A012,W3A022,W3A102,W3A112,W3A122,W3A202,W3A212,W3A222;
(*DONT_TOUCH="true"*) wire W3A003,W3A013,W3A023,W3A103,W3A113,W3A123,W3A203,W3A213,W3A223;
(*DONT_TOUCH="true"*) wire W3A004,W3A014,W3A024,W3A104,W3A114,W3A124,W3A204,W3A214,W3A224;
(*DONT_TOUCH="true"*) wire W3A005,W3A015,W3A025,W3A105,W3A115,W3A125,W3A205,W3A215,W3A225;
(*DONT_TOUCH="true"*) wire W3A006,W3A016,W3A026,W3A106,W3A116,W3A126,W3A206,W3A216,W3A226;
(*DONT_TOUCH="true"*) wire W3A007,W3A017,W3A027,W3A107,W3A117,W3A127,W3A207,W3A217,W3A227;
(*DONT_TOUCH="true"*) wire W3A008,W3A018,W3A028,W3A108,W3A118,W3A128,W3A208,W3A218,W3A228;
(*DONT_TOUCH="true"*) wire W3A009,W3A019,W3A029,W3A109,W3A119,W3A129,W3A209,W3A219,W3A229;
(*DONT_TOUCH="true"*) wire W3A00A,W3A01A,W3A02A,W3A10A,W3A11A,W3A12A,W3A20A,W3A21A,W3A22A;
(*DONT_TOUCH="true"*) wire W3A00B,W3A01B,W3A02B,W3A10B,W3A11B,W3A12B,W3A20B,W3A21B,W3A22B;
(*DONT_TOUCH="true"*) wire W3A00C,W3A01C,W3A02C,W3A10C,W3A11C,W3A12C,W3A20C,W3A21C,W3A22C;
(*DONT_TOUCH="true"*) wire W3A00D,W3A01D,W3A02D,W3A10D,W3A11D,W3A12D,W3A20D,W3A21D,W3A22D;
(*DONT_TOUCH="true"*) wire W3A00E,W3A01E,W3A02E,W3A10E,W3A11E,W3A12E,W3A20E,W3A21E,W3A22E;
(*DONT_TOUCH="true"*) wire W3A00F,W3A01F,W3A02F,W3A10F,W3A11F,W3A12F,W3A20F,W3A21F,W3A22F;
(*DONT_TOUCH="true"*) wire W3B000,W3B010,W3B020,W3B100,W3B110,W3B120,W3B200,W3B210,W3B220;
(*DONT_TOUCH="true"*) wire W3B001,W3B011,W3B021,W3B101,W3B111,W3B121,W3B201,W3B211,W3B221;
(*DONT_TOUCH="true"*) wire W3B002,W3B012,W3B022,W3B102,W3B112,W3B122,W3B202,W3B212,W3B222;
(*DONT_TOUCH="true"*) wire W3B003,W3B013,W3B023,W3B103,W3B113,W3B123,W3B203,W3B213,W3B223;
(*DONT_TOUCH="true"*) wire W3B004,W3B014,W3B024,W3B104,W3B114,W3B124,W3B204,W3B214,W3B224;
(*DONT_TOUCH="true"*) wire W3B005,W3B015,W3B025,W3B105,W3B115,W3B125,W3B205,W3B215,W3B225;
(*DONT_TOUCH="true"*) wire W3B006,W3B016,W3B026,W3B106,W3B116,W3B126,W3B206,W3B216,W3B226;
(*DONT_TOUCH="true"*) wire W3B007,W3B017,W3B027,W3B107,W3B117,W3B127,W3B207,W3B217,W3B227;
(*DONT_TOUCH="true"*) wire W3B008,W3B018,W3B028,W3B108,W3B118,W3B128,W3B208,W3B218,W3B228;
(*DONT_TOUCH="true"*) wire W3B009,W3B019,W3B029,W3B109,W3B119,W3B129,W3B209,W3B219,W3B229;
(*DONT_TOUCH="true"*) wire W3B00A,W3B01A,W3B02A,W3B10A,W3B11A,W3B12A,W3B20A,W3B21A,W3B22A;
(*DONT_TOUCH="true"*) wire W3B00B,W3B01B,W3B02B,W3B10B,W3B11B,W3B12B,W3B20B,W3B21B,W3B22B;
(*DONT_TOUCH="true"*) wire W3B00C,W3B01C,W3B02C,W3B10C,W3B11C,W3B12C,W3B20C,W3B21C,W3B22C;
(*DONT_TOUCH="true"*) wire W3B00D,W3B01D,W3B02D,W3B10D,W3B11D,W3B12D,W3B20D,W3B21D,W3B22D;
(*DONT_TOUCH="true"*) wire W3B00E,W3B01E,W3B02E,W3B10E,W3B11E,W3B12E,W3B20E,W3B21E,W3B22E;
(*DONT_TOUCH="true"*) wire W3B00F,W3B01F,W3B02F,W3B10F,W3B11F,W3B12F,W3B20F,W3B21F,W3B22F;
(*DONT_TOUCH="true"*) wire W3C000,W3C010,W3C020,W3C100,W3C110,W3C120,W3C200,W3C210,W3C220;
(*DONT_TOUCH="true"*) wire W3C001,W3C011,W3C021,W3C101,W3C111,W3C121,W3C201,W3C211,W3C221;
(*DONT_TOUCH="true"*) wire W3C002,W3C012,W3C022,W3C102,W3C112,W3C122,W3C202,W3C212,W3C222;
(*DONT_TOUCH="true"*) wire W3C003,W3C013,W3C023,W3C103,W3C113,W3C123,W3C203,W3C213,W3C223;
(*DONT_TOUCH="true"*) wire W3C004,W3C014,W3C024,W3C104,W3C114,W3C124,W3C204,W3C214,W3C224;
(*DONT_TOUCH="true"*) wire W3C005,W3C015,W3C025,W3C105,W3C115,W3C125,W3C205,W3C215,W3C225;
(*DONT_TOUCH="true"*) wire W3C006,W3C016,W3C026,W3C106,W3C116,W3C126,W3C206,W3C216,W3C226;
(*DONT_TOUCH="true"*) wire W3C007,W3C017,W3C027,W3C107,W3C117,W3C127,W3C207,W3C217,W3C227;
(*DONT_TOUCH="true"*) wire W3C008,W3C018,W3C028,W3C108,W3C118,W3C128,W3C208,W3C218,W3C228;
(*DONT_TOUCH="true"*) wire W3C009,W3C019,W3C029,W3C109,W3C119,W3C129,W3C209,W3C219,W3C229;
(*DONT_TOUCH="true"*) wire W3C00A,W3C01A,W3C02A,W3C10A,W3C11A,W3C12A,W3C20A,W3C21A,W3C22A;
(*DONT_TOUCH="true"*) wire W3C00B,W3C01B,W3C02B,W3C10B,W3C11B,W3C12B,W3C20B,W3C21B,W3C22B;
(*DONT_TOUCH="true"*) wire W3C00C,W3C01C,W3C02C,W3C10C,W3C11C,W3C12C,W3C20C,W3C21C,W3C22C;
(*DONT_TOUCH="true"*) wire W3C00D,W3C01D,W3C02D,W3C10D,W3C11D,W3C12D,W3C20D,W3C21D,W3C22D;
(*DONT_TOUCH="true"*) wire W3C00E,W3C01E,W3C02E,W3C10E,W3C11E,W3C12E,W3C20E,W3C21E,W3C22E;
(*DONT_TOUCH="true"*) wire W3C00F,W3C01F,W3C02F,W3C10F,W3C11F,W3C12F,W3C20F,W3C21F,W3C22F;
(*DONT_TOUCH="true"*) wire W3D000,W3D010,W3D020,W3D100,W3D110,W3D120,W3D200,W3D210,W3D220;
(*DONT_TOUCH="true"*) wire W3D001,W3D011,W3D021,W3D101,W3D111,W3D121,W3D201,W3D211,W3D221;
(*DONT_TOUCH="true"*) wire W3D002,W3D012,W3D022,W3D102,W3D112,W3D122,W3D202,W3D212,W3D222;
(*DONT_TOUCH="true"*) wire W3D003,W3D013,W3D023,W3D103,W3D113,W3D123,W3D203,W3D213,W3D223;
(*DONT_TOUCH="true"*) wire W3D004,W3D014,W3D024,W3D104,W3D114,W3D124,W3D204,W3D214,W3D224;
(*DONT_TOUCH="true"*) wire W3D005,W3D015,W3D025,W3D105,W3D115,W3D125,W3D205,W3D215,W3D225;
(*DONT_TOUCH="true"*) wire W3D006,W3D016,W3D026,W3D106,W3D116,W3D126,W3D206,W3D216,W3D226;
(*DONT_TOUCH="true"*) wire W3D007,W3D017,W3D027,W3D107,W3D117,W3D127,W3D207,W3D217,W3D227;
(*DONT_TOUCH="true"*) wire W3D008,W3D018,W3D028,W3D108,W3D118,W3D128,W3D208,W3D218,W3D228;
(*DONT_TOUCH="true"*) wire W3D009,W3D019,W3D029,W3D109,W3D119,W3D129,W3D209,W3D219,W3D229;
(*DONT_TOUCH="true"*) wire W3D00A,W3D01A,W3D02A,W3D10A,W3D11A,W3D12A,W3D20A,W3D21A,W3D22A;
(*DONT_TOUCH="true"*) wire W3D00B,W3D01B,W3D02B,W3D10B,W3D11B,W3D12B,W3D20B,W3D21B,W3D22B;
(*DONT_TOUCH="true"*) wire W3D00C,W3D01C,W3D02C,W3D10C,W3D11C,W3D12C,W3D20C,W3D21C,W3D22C;
(*DONT_TOUCH="true"*) wire W3D00D,W3D01D,W3D02D,W3D10D,W3D11D,W3D12D,W3D20D,W3D21D,W3D22D;
(*DONT_TOUCH="true"*) wire W3D00E,W3D01E,W3D02E,W3D10E,W3D11E,W3D12E,W3D20E,W3D21E,W3D22E;
(*DONT_TOUCH="true"*) wire W3D00F,W3D01F,W3D02F,W3D10F,W3D11F,W3D12F,W3D20F,W3D21F,W3D22F;
(*DONT_TOUCH="true"*) wire W3E000,W3E010,W3E020,W3E100,W3E110,W3E120,W3E200,W3E210,W3E220;
(*DONT_TOUCH="true"*) wire W3E001,W3E011,W3E021,W3E101,W3E111,W3E121,W3E201,W3E211,W3E221;
(*DONT_TOUCH="true"*) wire W3E002,W3E012,W3E022,W3E102,W3E112,W3E122,W3E202,W3E212,W3E222;
(*DONT_TOUCH="true"*) wire W3E003,W3E013,W3E023,W3E103,W3E113,W3E123,W3E203,W3E213,W3E223;
(*DONT_TOUCH="true"*) wire W3E004,W3E014,W3E024,W3E104,W3E114,W3E124,W3E204,W3E214,W3E224;
(*DONT_TOUCH="true"*) wire W3E005,W3E015,W3E025,W3E105,W3E115,W3E125,W3E205,W3E215,W3E225;
(*DONT_TOUCH="true"*) wire W3E006,W3E016,W3E026,W3E106,W3E116,W3E126,W3E206,W3E216,W3E226;
(*DONT_TOUCH="true"*) wire W3E007,W3E017,W3E027,W3E107,W3E117,W3E127,W3E207,W3E217,W3E227;
(*DONT_TOUCH="true"*) wire W3E008,W3E018,W3E028,W3E108,W3E118,W3E128,W3E208,W3E218,W3E228;
(*DONT_TOUCH="true"*) wire W3E009,W3E019,W3E029,W3E109,W3E119,W3E129,W3E209,W3E219,W3E229;
(*DONT_TOUCH="true"*) wire W3E00A,W3E01A,W3E02A,W3E10A,W3E11A,W3E12A,W3E20A,W3E21A,W3E22A;
(*DONT_TOUCH="true"*) wire W3E00B,W3E01B,W3E02B,W3E10B,W3E11B,W3E12B,W3E20B,W3E21B,W3E22B;
(*DONT_TOUCH="true"*) wire W3E00C,W3E01C,W3E02C,W3E10C,W3E11C,W3E12C,W3E20C,W3E21C,W3E22C;
(*DONT_TOUCH="true"*) wire W3E00D,W3E01D,W3E02D,W3E10D,W3E11D,W3E12D,W3E20D,W3E21D,W3E22D;
(*DONT_TOUCH="true"*) wire W3E00E,W3E01E,W3E02E,W3E10E,W3E11E,W3E12E,W3E20E,W3E21E,W3E22E;
(*DONT_TOUCH="true"*) wire W3E00F,W3E01F,W3E02F,W3E10F,W3E11F,W3E12F,W3E20F,W3E21F,W3E22F;
(*DONT_TOUCH="true"*) wire W3F000,W3F010,W3F020,W3F100,W3F110,W3F120,W3F200,W3F210,W3F220;
(*DONT_TOUCH="true"*) wire W3F001,W3F011,W3F021,W3F101,W3F111,W3F121,W3F201,W3F211,W3F221;
(*DONT_TOUCH="true"*) wire W3F002,W3F012,W3F022,W3F102,W3F112,W3F122,W3F202,W3F212,W3F222;
(*DONT_TOUCH="true"*) wire W3F003,W3F013,W3F023,W3F103,W3F113,W3F123,W3F203,W3F213,W3F223;
(*DONT_TOUCH="true"*) wire W3F004,W3F014,W3F024,W3F104,W3F114,W3F124,W3F204,W3F214,W3F224;
(*DONT_TOUCH="true"*) wire W3F005,W3F015,W3F025,W3F105,W3F115,W3F125,W3F205,W3F215,W3F225;
(*DONT_TOUCH="true"*) wire W3F006,W3F016,W3F026,W3F106,W3F116,W3F126,W3F206,W3F216,W3F226;
(*DONT_TOUCH="true"*) wire W3F007,W3F017,W3F027,W3F107,W3F117,W3F127,W3F207,W3F217,W3F227;
(*DONT_TOUCH="true"*) wire W3F008,W3F018,W3F028,W3F108,W3F118,W3F128,W3F208,W3F218,W3F228;
(*DONT_TOUCH="true"*) wire W3F009,W3F019,W3F029,W3F109,W3F119,W3F129,W3F209,W3F219,W3F229;
(*DONT_TOUCH="true"*) wire W3F00A,W3F01A,W3F02A,W3F10A,W3F11A,W3F12A,W3F20A,W3F21A,W3F22A;
(*DONT_TOUCH="true"*) wire W3F00B,W3F01B,W3F02B,W3F10B,W3F11B,W3F12B,W3F20B,W3F21B,W3F22B;
(*DONT_TOUCH="true"*) wire W3F00C,W3F01C,W3F02C,W3F10C,W3F11C,W3F12C,W3F20C,W3F21C,W3F22C;
(*DONT_TOUCH="true"*) wire W3F00D,W3F01D,W3F02D,W3F10D,W3F11D,W3F12D,W3F20D,W3F21D,W3F22D;
(*DONT_TOUCH="true"*) wire W3F00E,W3F01E,W3F02E,W3F10E,W3F11E,W3F12E,W3F20E,W3F21E,W3F22E;
(*DONT_TOUCH="true"*) wire W3F00F,W3F01F,W3F02F,W3F10F,W3F11F,W3F12F,W3F20F,W3F21F,W3F22F;
(*DONT_TOUCH="true"*) wire W3G000,W3G010,W3G020,W3G100,W3G110,W3G120,W3G200,W3G210,W3G220;
(*DONT_TOUCH="true"*) wire W3G001,W3G011,W3G021,W3G101,W3G111,W3G121,W3G201,W3G211,W3G221;
(*DONT_TOUCH="true"*) wire W3G002,W3G012,W3G022,W3G102,W3G112,W3G122,W3G202,W3G212,W3G222;
(*DONT_TOUCH="true"*) wire W3G003,W3G013,W3G023,W3G103,W3G113,W3G123,W3G203,W3G213,W3G223;
(*DONT_TOUCH="true"*) wire W3G004,W3G014,W3G024,W3G104,W3G114,W3G124,W3G204,W3G214,W3G224;
(*DONT_TOUCH="true"*) wire W3G005,W3G015,W3G025,W3G105,W3G115,W3G125,W3G205,W3G215,W3G225;
(*DONT_TOUCH="true"*) wire W3G006,W3G016,W3G026,W3G106,W3G116,W3G126,W3G206,W3G216,W3G226;
(*DONT_TOUCH="true"*) wire W3G007,W3G017,W3G027,W3G107,W3G117,W3G127,W3G207,W3G217,W3G227;
(*DONT_TOUCH="true"*) wire W3G008,W3G018,W3G028,W3G108,W3G118,W3G128,W3G208,W3G218,W3G228;
(*DONT_TOUCH="true"*) wire W3G009,W3G019,W3G029,W3G109,W3G119,W3G129,W3G209,W3G219,W3G229;
(*DONT_TOUCH="true"*) wire W3G00A,W3G01A,W3G02A,W3G10A,W3G11A,W3G12A,W3G20A,W3G21A,W3G22A;
(*DONT_TOUCH="true"*) wire W3G00B,W3G01B,W3G02B,W3G10B,W3G11B,W3G12B,W3G20B,W3G21B,W3G22B;
(*DONT_TOUCH="true"*) wire W3G00C,W3G01C,W3G02C,W3G10C,W3G11C,W3G12C,W3G20C,W3G21C,W3G22C;
(*DONT_TOUCH="true"*) wire W3G00D,W3G01D,W3G02D,W3G10D,W3G11D,W3G12D,W3G20D,W3G21D,W3G22D;
(*DONT_TOUCH="true"*) wire W3G00E,W3G01E,W3G02E,W3G10E,W3G11E,W3G12E,W3G20E,W3G21E,W3G22E;
(*DONT_TOUCH="true"*) wire W3G00F,W3G01F,W3G02F,W3G10F,W3G11F,W3G12F,W3G20F,W3G21F,W3G22F;
(*DONT_TOUCH="true"*) wire W3H000,W3H010,W3H020,W3H100,W3H110,W3H120,W3H200,W3H210,W3H220;
(*DONT_TOUCH="true"*) wire W3H001,W3H011,W3H021,W3H101,W3H111,W3H121,W3H201,W3H211,W3H221;
(*DONT_TOUCH="true"*) wire W3H002,W3H012,W3H022,W3H102,W3H112,W3H122,W3H202,W3H212,W3H222;
(*DONT_TOUCH="true"*) wire W3H003,W3H013,W3H023,W3H103,W3H113,W3H123,W3H203,W3H213,W3H223;
(*DONT_TOUCH="true"*) wire W3H004,W3H014,W3H024,W3H104,W3H114,W3H124,W3H204,W3H214,W3H224;
(*DONT_TOUCH="true"*) wire W3H005,W3H015,W3H025,W3H105,W3H115,W3H125,W3H205,W3H215,W3H225;
(*DONT_TOUCH="true"*) wire W3H006,W3H016,W3H026,W3H106,W3H116,W3H126,W3H206,W3H216,W3H226;
(*DONT_TOUCH="true"*) wire W3H007,W3H017,W3H027,W3H107,W3H117,W3H127,W3H207,W3H217,W3H227;
(*DONT_TOUCH="true"*) wire W3H008,W3H018,W3H028,W3H108,W3H118,W3H128,W3H208,W3H218,W3H228;
(*DONT_TOUCH="true"*) wire W3H009,W3H019,W3H029,W3H109,W3H119,W3H129,W3H209,W3H219,W3H229;
(*DONT_TOUCH="true"*) wire W3H00A,W3H01A,W3H02A,W3H10A,W3H11A,W3H12A,W3H20A,W3H21A,W3H22A;
(*DONT_TOUCH="true"*) wire W3H00B,W3H01B,W3H02B,W3H10B,W3H11B,W3H12B,W3H20B,W3H21B,W3H22B;
(*DONT_TOUCH="true"*) wire W3H00C,W3H01C,W3H02C,W3H10C,W3H11C,W3H12C,W3H20C,W3H21C,W3H22C;
(*DONT_TOUCH="true"*) wire W3H00D,W3H01D,W3H02D,W3H10D,W3H11D,W3H12D,W3H20D,W3H21D,W3H22D;
(*DONT_TOUCH="true"*) wire W3H00E,W3H01E,W3H02E,W3H10E,W3H11E,W3H12E,W3H20E,W3H21E,W3H22E;
(*DONT_TOUCH="true"*) wire W3H00F,W3H01F,W3H02F,W3H10F,W3H11F,W3H12F,W3H20F,W3H21F,W3H22F;
(*DONT_TOUCH="true"*) wire W3I000,W3I010,W3I020,W3I100,W3I110,W3I120,W3I200,W3I210,W3I220;
(*DONT_TOUCH="true"*) wire W3I001,W3I011,W3I021,W3I101,W3I111,W3I121,W3I201,W3I211,W3I221;
(*DONT_TOUCH="true"*) wire W3I002,W3I012,W3I022,W3I102,W3I112,W3I122,W3I202,W3I212,W3I222;
(*DONT_TOUCH="true"*) wire W3I003,W3I013,W3I023,W3I103,W3I113,W3I123,W3I203,W3I213,W3I223;
(*DONT_TOUCH="true"*) wire W3I004,W3I014,W3I024,W3I104,W3I114,W3I124,W3I204,W3I214,W3I224;
(*DONT_TOUCH="true"*) wire W3I005,W3I015,W3I025,W3I105,W3I115,W3I125,W3I205,W3I215,W3I225;
(*DONT_TOUCH="true"*) wire W3I006,W3I016,W3I026,W3I106,W3I116,W3I126,W3I206,W3I216,W3I226;
(*DONT_TOUCH="true"*) wire W3I007,W3I017,W3I027,W3I107,W3I117,W3I127,W3I207,W3I217,W3I227;
(*DONT_TOUCH="true"*) wire W3I008,W3I018,W3I028,W3I108,W3I118,W3I128,W3I208,W3I218,W3I228;
(*DONT_TOUCH="true"*) wire W3I009,W3I019,W3I029,W3I109,W3I119,W3I129,W3I209,W3I219,W3I229;
(*DONT_TOUCH="true"*) wire W3I00A,W3I01A,W3I02A,W3I10A,W3I11A,W3I12A,W3I20A,W3I21A,W3I22A;
(*DONT_TOUCH="true"*) wire W3I00B,W3I01B,W3I02B,W3I10B,W3I11B,W3I12B,W3I20B,W3I21B,W3I22B;
(*DONT_TOUCH="true"*) wire W3I00C,W3I01C,W3I02C,W3I10C,W3I11C,W3I12C,W3I20C,W3I21C,W3I22C;
(*DONT_TOUCH="true"*) wire W3I00D,W3I01D,W3I02D,W3I10D,W3I11D,W3I12D,W3I20D,W3I21D,W3I22D;
(*DONT_TOUCH="true"*) wire W3I00E,W3I01E,W3I02E,W3I10E,W3I11E,W3I12E,W3I20E,W3I21E,W3I22E;
(*DONT_TOUCH="true"*) wire W3I00F,W3I01F,W3I02F,W3I10F,W3I11F,W3I12F,W3I20F,W3I21F,W3I22F;
(*DONT_TOUCH="true"*) wire W3J000,W3J010,W3J020,W3J100,W3J110,W3J120,W3J200,W3J210,W3J220;
(*DONT_TOUCH="true"*) wire W3J001,W3J011,W3J021,W3J101,W3J111,W3J121,W3J201,W3J211,W3J221;
(*DONT_TOUCH="true"*) wire W3J002,W3J012,W3J022,W3J102,W3J112,W3J122,W3J202,W3J212,W3J222;
(*DONT_TOUCH="true"*) wire W3J003,W3J013,W3J023,W3J103,W3J113,W3J123,W3J203,W3J213,W3J223;
(*DONT_TOUCH="true"*) wire W3J004,W3J014,W3J024,W3J104,W3J114,W3J124,W3J204,W3J214,W3J224;
(*DONT_TOUCH="true"*) wire W3J005,W3J015,W3J025,W3J105,W3J115,W3J125,W3J205,W3J215,W3J225;
(*DONT_TOUCH="true"*) wire W3J006,W3J016,W3J026,W3J106,W3J116,W3J126,W3J206,W3J216,W3J226;
(*DONT_TOUCH="true"*) wire W3J007,W3J017,W3J027,W3J107,W3J117,W3J127,W3J207,W3J217,W3J227;
(*DONT_TOUCH="true"*) wire W3J008,W3J018,W3J028,W3J108,W3J118,W3J128,W3J208,W3J218,W3J228;
(*DONT_TOUCH="true"*) wire W3J009,W3J019,W3J029,W3J109,W3J119,W3J129,W3J209,W3J219,W3J229;
(*DONT_TOUCH="true"*) wire W3J00A,W3J01A,W3J02A,W3J10A,W3J11A,W3J12A,W3J20A,W3J21A,W3J22A;
(*DONT_TOUCH="true"*) wire W3J00B,W3J01B,W3J02B,W3J10B,W3J11B,W3J12B,W3J20B,W3J21B,W3J22B;
(*DONT_TOUCH="true"*) wire W3J00C,W3J01C,W3J02C,W3J10C,W3J11C,W3J12C,W3J20C,W3J21C,W3J22C;
(*DONT_TOUCH="true"*) wire W3J00D,W3J01D,W3J02D,W3J10D,W3J11D,W3J12D,W3J20D,W3J21D,W3J22D;
(*DONT_TOUCH="true"*) wire W3J00E,W3J01E,W3J02E,W3J10E,W3J11E,W3J12E,W3J20E,W3J21E,W3J22E;
(*DONT_TOUCH="true"*) wire W3J00F,W3J01F,W3J02F,W3J10F,W3J11F,W3J12F,W3J20F,W3J21F,W3J22F;
(*DONT_TOUCH="true"*) wire W3K000,W3K010,W3K020,W3K100,W3K110,W3K120,W3K200,W3K210,W3K220;
(*DONT_TOUCH="true"*) wire W3K001,W3K011,W3K021,W3K101,W3K111,W3K121,W3K201,W3K211,W3K221;
(*DONT_TOUCH="true"*) wire W3K002,W3K012,W3K022,W3K102,W3K112,W3K122,W3K202,W3K212,W3K222;
(*DONT_TOUCH="true"*) wire W3K003,W3K013,W3K023,W3K103,W3K113,W3K123,W3K203,W3K213,W3K223;
(*DONT_TOUCH="true"*) wire W3K004,W3K014,W3K024,W3K104,W3K114,W3K124,W3K204,W3K214,W3K224;
(*DONT_TOUCH="true"*) wire W3K005,W3K015,W3K025,W3K105,W3K115,W3K125,W3K205,W3K215,W3K225;
(*DONT_TOUCH="true"*) wire W3K006,W3K016,W3K026,W3K106,W3K116,W3K126,W3K206,W3K216,W3K226;
(*DONT_TOUCH="true"*) wire W3K007,W3K017,W3K027,W3K107,W3K117,W3K127,W3K207,W3K217,W3K227;
(*DONT_TOUCH="true"*) wire W3K008,W3K018,W3K028,W3K108,W3K118,W3K128,W3K208,W3K218,W3K228;
(*DONT_TOUCH="true"*) wire W3K009,W3K019,W3K029,W3K109,W3K119,W3K129,W3K209,W3K219,W3K229;
(*DONT_TOUCH="true"*) wire W3K00A,W3K01A,W3K02A,W3K10A,W3K11A,W3K12A,W3K20A,W3K21A,W3K22A;
(*DONT_TOUCH="true"*) wire W3K00B,W3K01B,W3K02B,W3K10B,W3K11B,W3K12B,W3K20B,W3K21B,W3K22B;
(*DONT_TOUCH="true"*) wire W3K00C,W3K01C,W3K02C,W3K10C,W3K11C,W3K12C,W3K20C,W3K21C,W3K22C;
(*DONT_TOUCH="true"*) wire W3K00D,W3K01D,W3K02D,W3K10D,W3K11D,W3K12D,W3K20D,W3K21D,W3K22D;
(*DONT_TOUCH="true"*) wire W3K00E,W3K01E,W3K02E,W3K10E,W3K11E,W3K12E,W3K20E,W3K21E,W3K22E;
(*DONT_TOUCH="true"*) wire W3K00F,W3K01F,W3K02F,W3K10F,W3K11F,W3K12F,W3K20F,W3K21F,W3K22F;
(*DONT_TOUCH="true"*) wire W3L000,W3L010,W3L020,W3L100,W3L110,W3L120,W3L200,W3L210,W3L220;
(*DONT_TOUCH="true"*) wire W3L001,W3L011,W3L021,W3L101,W3L111,W3L121,W3L201,W3L211,W3L221;
(*DONT_TOUCH="true"*) wire W3L002,W3L012,W3L022,W3L102,W3L112,W3L122,W3L202,W3L212,W3L222;
(*DONT_TOUCH="true"*) wire W3L003,W3L013,W3L023,W3L103,W3L113,W3L123,W3L203,W3L213,W3L223;
(*DONT_TOUCH="true"*) wire W3L004,W3L014,W3L024,W3L104,W3L114,W3L124,W3L204,W3L214,W3L224;
(*DONT_TOUCH="true"*) wire W3L005,W3L015,W3L025,W3L105,W3L115,W3L125,W3L205,W3L215,W3L225;
(*DONT_TOUCH="true"*) wire W3L006,W3L016,W3L026,W3L106,W3L116,W3L126,W3L206,W3L216,W3L226;
(*DONT_TOUCH="true"*) wire W3L007,W3L017,W3L027,W3L107,W3L117,W3L127,W3L207,W3L217,W3L227;
(*DONT_TOUCH="true"*) wire W3L008,W3L018,W3L028,W3L108,W3L118,W3L128,W3L208,W3L218,W3L228;
(*DONT_TOUCH="true"*) wire W3L009,W3L019,W3L029,W3L109,W3L119,W3L129,W3L209,W3L219,W3L229;
(*DONT_TOUCH="true"*) wire W3L00A,W3L01A,W3L02A,W3L10A,W3L11A,W3L12A,W3L20A,W3L21A,W3L22A;
(*DONT_TOUCH="true"*) wire W3L00B,W3L01B,W3L02B,W3L10B,W3L11B,W3L12B,W3L20B,W3L21B,W3L22B;
(*DONT_TOUCH="true"*) wire W3L00C,W3L01C,W3L02C,W3L10C,W3L11C,W3L12C,W3L20C,W3L21C,W3L22C;
(*DONT_TOUCH="true"*) wire W3L00D,W3L01D,W3L02D,W3L10D,W3L11D,W3L12D,W3L20D,W3L21D,W3L22D;
(*DONT_TOUCH="true"*) wire W3L00E,W3L01E,W3L02E,W3L10E,W3L11E,W3L12E,W3L20E,W3L21E,W3L22E;
(*DONT_TOUCH="true"*) wire W3L00F,W3L01F,W3L02F,W3L10F,W3L11F,W3L12F,W3L20F,W3L21F,W3L22F;
(*DONT_TOUCH="true"*) wire W3M000,W3M010,W3M020,W3M100,W3M110,W3M120,W3M200,W3M210,W3M220;
(*DONT_TOUCH="true"*) wire W3M001,W3M011,W3M021,W3M101,W3M111,W3M121,W3M201,W3M211,W3M221;
(*DONT_TOUCH="true"*) wire W3M002,W3M012,W3M022,W3M102,W3M112,W3M122,W3M202,W3M212,W3M222;
(*DONT_TOUCH="true"*) wire W3M003,W3M013,W3M023,W3M103,W3M113,W3M123,W3M203,W3M213,W3M223;
(*DONT_TOUCH="true"*) wire W3M004,W3M014,W3M024,W3M104,W3M114,W3M124,W3M204,W3M214,W3M224;
(*DONT_TOUCH="true"*) wire W3M005,W3M015,W3M025,W3M105,W3M115,W3M125,W3M205,W3M215,W3M225;
(*DONT_TOUCH="true"*) wire W3M006,W3M016,W3M026,W3M106,W3M116,W3M126,W3M206,W3M216,W3M226;
(*DONT_TOUCH="true"*) wire W3M007,W3M017,W3M027,W3M107,W3M117,W3M127,W3M207,W3M217,W3M227;
(*DONT_TOUCH="true"*) wire W3M008,W3M018,W3M028,W3M108,W3M118,W3M128,W3M208,W3M218,W3M228;
(*DONT_TOUCH="true"*) wire W3M009,W3M019,W3M029,W3M109,W3M119,W3M129,W3M209,W3M219,W3M229;
(*DONT_TOUCH="true"*) wire W3M00A,W3M01A,W3M02A,W3M10A,W3M11A,W3M12A,W3M20A,W3M21A,W3M22A;
(*DONT_TOUCH="true"*) wire W3M00B,W3M01B,W3M02B,W3M10B,W3M11B,W3M12B,W3M20B,W3M21B,W3M22B;
(*DONT_TOUCH="true"*) wire W3M00C,W3M01C,W3M02C,W3M10C,W3M11C,W3M12C,W3M20C,W3M21C,W3M22C;
(*DONT_TOUCH="true"*) wire W3M00D,W3M01D,W3M02D,W3M10D,W3M11D,W3M12D,W3M20D,W3M21D,W3M22D;
(*DONT_TOUCH="true"*) wire W3M00E,W3M01E,W3M02E,W3M10E,W3M11E,W3M12E,W3M20E,W3M21E,W3M22E;
(*DONT_TOUCH="true"*) wire W3M00F,W3M01F,W3M02F,W3M10F,W3M11F,W3M12F,W3M20F,W3M21F,W3M22F;
(*DONT_TOUCH="true"*) wire W3N000,W3N010,W3N020,W3N100,W3N110,W3N120,W3N200,W3N210,W3N220;
(*DONT_TOUCH="true"*) wire W3N001,W3N011,W3N021,W3N101,W3N111,W3N121,W3N201,W3N211,W3N221;
(*DONT_TOUCH="true"*) wire W3N002,W3N012,W3N022,W3N102,W3N112,W3N122,W3N202,W3N212,W3N222;
(*DONT_TOUCH="true"*) wire W3N003,W3N013,W3N023,W3N103,W3N113,W3N123,W3N203,W3N213,W3N223;
(*DONT_TOUCH="true"*) wire W3N004,W3N014,W3N024,W3N104,W3N114,W3N124,W3N204,W3N214,W3N224;
(*DONT_TOUCH="true"*) wire W3N005,W3N015,W3N025,W3N105,W3N115,W3N125,W3N205,W3N215,W3N225;
(*DONT_TOUCH="true"*) wire W3N006,W3N016,W3N026,W3N106,W3N116,W3N126,W3N206,W3N216,W3N226;
(*DONT_TOUCH="true"*) wire W3N007,W3N017,W3N027,W3N107,W3N117,W3N127,W3N207,W3N217,W3N227;
(*DONT_TOUCH="true"*) wire W3N008,W3N018,W3N028,W3N108,W3N118,W3N128,W3N208,W3N218,W3N228;
(*DONT_TOUCH="true"*) wire W3N009,W3N019,W3N029,W3N109,W3N119,W3N129,W3N209,W3N219,W3N229;
(*DONT_TOUCH="true"*) wire W3N00A,W3N01A,W3N02A,W3N10A,W3N11A,W3N12A,W3N20A,W3N21A,W3N22A;
(*DONT_TOUCH="true"*) wire W3N00B,W3N01B,W3N02B,W3N10B,W3N11B,W3N12B,W3N20B,W3N21B,W3N22B;
(*DONT_TOUCH="true"*) wire W3N00C,W3N01C,W3N02C,W3N10C,W3N11C,W3N12C,W3N20C,W3N21C,W3N22C;
(*DONT_TOUCH="true"*) wire W3N00D,W3N01D,W3N02D,W3N10D,W3N11D,W3N12D,W3N20D,W3N21D,W3N22D;
(*DONT_TOUCH="true"*) wire W3N00E,W3N01E,W3N02E,W3N10E,W3N11E,W3N12E,W3N20E,W3N21E,W3N22E;
(*DONT_TOUCH="true"*) wire W3N00F,W3N01F,W3N02F,W3N10F,W3N11F,W3N12F,W3N20F,W3N21F,W3N22F;
(*DONT_TOUCH="true"*) wire W3O000,W3O010,W3O020,W3O100,W3O110,W3O120,W3O200,W3O210,W3O220;
(*DONT_TOUCH="true"*) wire W3O001,W3O011,W3O021,W3O101,W3O111,W3O121,W3O201,W3O211,W3O221;
(*DONT_TOUCH="true"*) wire W3O002,W3O012,W3O022,W3O102,W3O112,W3O122,W3O202,W3O212,W3O222;
(*DONT_TOUCH="true"*) wire W3O003,W3O013,W3O023,W3O103,W3O113,W3O123,W3O203,W3O213,W3O223;
(*DONT_TOUCH="true"*) wire W3O004,W3O014,W3O024,W3O104,W3O114,W3O124,W3O204,W3O214,W3O224;
(*DONT_TOUCH="true"*) wire W3O005,W3O015,W3O025,W3O105,W3O115,W3O125,W3O205,W3O215,W3O225;
(*DONT_TOUCH="true"*) wire W3O006,W3O016,W3O026,W3O106,W3O116,W3O126,W3O206,W3O216,W3O226;
(*DONT_TOUCH="true"*) wire W3O007,W3O017,W3O027,W3O107,W3O117,W3O127,W3O207,W3O217,W3O227;
(*DONT_TOUCH="true"*) wire W3O008,W3O018,W3O028,W3O108,W3O118,W3O128,W3O208,W3O218,W3O228;
(*DONT_TOUCH="true"*) wire W3O009,W3O019,W3O029,W3O109,W3O119,W3O129,W3O209,W3O219,W3O229;
(*DONT_TOUCH="true"*) wire W3O00A,W3O01A,W3O02A,W3O10A,W3O11A,W3O12A,W3O20A,W3O21A,W3O22A;
(*DONT_TOUCH="true"*) wire W3O00B,W3O01B,W3O02B,W3O10B,W3O11B,W3O12B,W3O20B,W3O21B,W3O22B;
(*DONT_TOUCH="true"*) wire W3O00C,W3O01C,W3O02C,W3O10C,W3O11C,W3O12C,W3O20C,W3O21C,W3O22C;
(*DONT_TOUCH="true"*) wire W3O00D,W3O01D,W3O02D,W3O10D,W3O11D,W3O12D,W3O20D,W3O21D,W3O22D;
(*DONT_TOUCH="true"*) wire W3O00E,W3O01E,W3O02E,W3O10E,W3O11E,W3O12E,W3O20E,W3O21E,W3O22E;
(*DONT_TOUCH="true"*) wire W3O00F,W3O01F,W3O02F,W3O10F,W3O11F,W3O12F,W3O20F,W3O21F,W3O22F;
(*DONT_TOUCH="true"*) wire W3P000,W3P010,W3P020,W3P100,W3P110,W3P120,W3P200,W3P210,W3P220;
(*DONT_TOUCH="true"*) wire W3P001,W3P011,W3P021,W3P101,W3P111,W3P121,W3P201,W3P211,W3P221;
(*DONT_TOUCH="true"*) wire W3P002,W3P012,W3P022,W3P102,W3P112,W3P122,W3P202,W3P212,W3P222;
(*DONT_TOUCH="true"*) wire W3P003,W3P013,W3P023,W3P103,W3P113,W3P123,W3P203,W3P213,W3P223;
(*DONT_TOUCH="true"*) wire W3P004,W3P014,W3P024,W3P104,W3P114,W3P124,W3P204,W3P214,W3P224;
(*DONT_TOUCH="true"*) wire W3P005,W3P015,W3P025,W3P105,W3P115,W3P125,W3P205,W3P215,W3P225;
(*DONT_TOUCH="true"*) wire W3P006,W3P016,W3P026,W3P106,W3P116,W3P126,W3P206,W3P216,W3P226;
(*DONT_TOUCH="true"*) wire W3P007,W3P017,W3P027,W3P107,W3P117,W3P127,W3P207,W3P217,W3P227;
(*DONT_TOUCH="true"*) wire W3P008,W3P018,W3P028,W3P108,W3P118,W3P128,W3P208,W3P218,W3P228;
(*DONT_TOUCH="true"*) wire W3P009,W3P019,W3P029,W3P109,W3P119,W3P129,W3P209,W3P219,W3P229;
(*DONT_TOUCH="true"*) wire W3P00A,W3P01A,W3P02A,W3P10A,W3P11A,W3P12A,W3P20A,W3P21A,W3P22A;
(*DONT_TOUCH="true"*) wire W3P00B,W3P01B,W3P02B,W3P10B,W3P11B,W3P12B,W3P20B,W3P21B,W3P22B;
(*DONT_TOUCH="true"*) wire W3P00C,W3P01C,W3P02C,W3P10C,W3P11C,W3P12C,W3P20C,W3P21C,W3P22C;
(*DONT_TOUCH="true"*) wire W3P00D,W3P01D,W3P02D,W3P10D,W3P11D,W3P12D,W3P20D,W3P21D,W3P22D;
(*DONT_TOUCH="true"*) wire W3P00E,W3P01E,W3P02E,W3P10E,W3P11E,W3P12E,W3P20E,W3P21E,W3P22E;
(*DONT_TOUCH="true"*) wire W3P00F,W3P01F,W3P02F,W3P10F,W3P11F,W3P12F,W3P20F,W3P21F,W3P22F;
(*DONT_TOUCH="true"*) wire W3Q000,W3Q010,W3Q020,W3Q100,W3Q110,W3Q120,W3Q200,W3Q210,W3Q220;
(*DONT_TOUCH="true"*) wire W3Q001,W3Q011,W3Q021,W3Q101,W3Q111,W3Q121,W3Q201,W3Q211,W3Q221;
(*DONT_TOUCH="true"*) wire W3Q002,W3Q012,W3Q022,W3Q102,W3Q112,W3Q122,W3Q202,W3Q212,W3Q222;
(*DONT_TOUCH="true"*) wire W3Q003,W3Q013,W3Q023,W3Q103,W3Q113,W3Q123,W3Q203,W3Q213,W3Q223;
(*DONT_TOUCH="true"*) wire W3Q004,W3Q014,W3Q024,W3Q104,W3Q114,W3Q124,W3Q204,W3Q214,W3Q224;
(*DONT_TOUCH="true"*) wire W3Q005,W3Q015,W3Q025,W3Q105,W3Q115,W3Q125,W3Q205,W3Q215,W3Q225;
(*DONT_TOUCH="true"*) wire W3Q006,W3Q016,W3Q026,W3Q106,W3Q116,W3Q126,W3Q206,W3Q216,W3Q226;
(*DONT_TOUCH="true"*) wire W3Q007,W3Q017,W3Q027,W3Q107,W3Q117,W3Q127,W3Q207,W3Q217,W3Q227;
(*DONT_TOUCH="true"*) wire W3Q008,W3Q018,W3Q028,W3Q108,W3Q118,W3Q128,W3Q208,W3Q218,W3Q228;
(*DONT_TOUCH="true"*) wire W3Q009,W3Q019,W3Q029,W3Q109,W3Q119,W3Q129,W3Q209,W3Q219,W3Q229;
(*DONT_TOUCH="true"*) wire W3Q00A,W3Q01A,W3Q02A,W3Q10A,W3Q11A,W3Q12A,W3Q20A,W3Q21A,W3Q22A;
(*DONT_TOUCH="true"*) wire W3Q00B,W3Q01B,W3Q02B,W3Q10B,W3Q11B,W3Q12B,W3Q20B,W3Q21B,W3Q22B;
(*DONT_TOUCH="true"*) wire W3Q00C,W3Q01C,W3Q02C,W3Q10C,W3Q11C,W3Q12C,W3Q20C,W3Q21C,W3Q22C;
(*DONT_TOUCH="true"*) wire W3Q00D,W3Q01D,W3Q02D,W3Q10D,W3Q11D,W3Q12D,W3Q20D,W3Q21D,W3Q22D;
(*DONT_TOUCH="true"*) wire W3Q00E,W3Q01E,W3Q02E,W3Q10E,W3Q11E,W3Q12E,W3Q20E,W3Q21E,W3Q22E;
(*DONT_TOUCH="true"*) wire W3Q00F,W3Q01F,W3Q02F,W3Q10F,W3Q11F,W3Q12F,W3Q20F,W3Q21F,W3Q22F;
(*DONT_TOUCH="true"*) wire W3R000,W3R010,W3R020,W3R100,W3R110,W3R120,W3R200,W3R210,W3R220;
(*DONT_TOUCH="true"*) wire W3R001,W3R011,W3R021,W3R101,W3R111,W3R121,W3R201,W3R211,W3R221;
(*DONT_TOUCH="true"*) wire W3R002,W3R012,W3R022,W3R102,W3R112,W3R122,W3R202,W3R212,W3R222;
(*DONT_TOUCH="true"*) wire W3R003,W3R013,W3R023,W3R103,W3R113,W3R123,W3R203,W3R213,W3R223;
(*DONT_TOUCH="true"*) wire W3R004,W3R014,W3R024,W3R104,W3R114,W3R124,W3R204,W3R214,W3R224;
(*DONT_TOUCH="true"*) wire W3R005,W3R015,W3R025,W3R105,W3R115,W3R125,W3R205,W3R215,W3R225;
(*DONT_TOUCH="true"*) wire W3R006,W3R016,W3R026,W3R106,W3R116,W3R126,W3R206,W3R216,W3R226;
(*DONT_TOUCH="true"*) wire W3R007,W3R017,W3R027,W3R107,W3R117,W3R127,W3R207,W3R217,W3R227;
(*DONT_TOUCH="true"*) wire W3R008,W3R018,W3R028,W3R108,W3R118,W3R128,W3R208,W3R218,W3R228;
(*DONT_TOUCH="true"*) wire W3R009,W3R019,W3R029,W3R109,W3R119,W3R129,W3R209,W3R219,W3R229;
(*DONT_TOUCH="true"*) wire W3R00A,W3R01A,W3R02A,W3R10A,W3R11A,W3R12A,W3R20A,W3R21A,W3R22A;
(*DONT_TOUCH="true"*) wire W3R00B,W3R01B,W3R02B,W3R10B,W3R11B,W3R12B,W3R20B,W3R21B,W3R22B;
(*DONT_TOUCH="true"*) wire W3R00C,W3R01C,W3R02C,W3R10C,W3R11C,W3R12C,W3R20C,W3R21C,W3R22C;
(*DONT_TOUCH="true"*) wire W3R00D,W3R01D,W3R02D,W3R10D,W3R11D,W3R12D,W3R20D,W3R21D,W3R22D;
(*DONT_TOUCH="true"*) wire W3R00E,W3R01E,W3R02E,W3R10E,W3R11E,W3R12E,W3R20E,W3R21E,W3R22E;
(*DONT_TOUCH="true"*) wire W3R00F,W3R01F,W3R02F,W3R10F,W3R11F,W3R12F,W3R20F,W3R21F,W3R22F;
(*DONT_TOUCH="true"*) wire W3S000,W3S010,W3S020,W3S100,W3S110,W3S120,W3S200,W3S210,W3S220;
(*DONT_TOUCH="true"*) wire W3S001,W3S011,W3S021,W3S101,W3S111,W3S121,W3S201,W3S211,W3S221;
(*DONT_TOUCH="true"*) wire W3S002,W3S012,W3S022,W3S102,W3S112,W3S122,W3S202,W3S212,W3S222;
(*DONT_TOUCH="true"*) wire W3S003,W3S013,W3S023,W3S103,W3S113,W3S123,W3S203,W3S213,W3S223;
(*DONT_TOUCH="true"*) wire W3S004,W3S014,W3S024,W3S104,W3S114,W3S124,W3S204,W3S214,W3S224;
(*DONT_TOUCH="true"*) wire W3S005,W3S015,W3S025,W3S105,W3S115,W3S125,W3S205,W3S215,W3S225;
(*DONT_TOUCH="true"*) wire W3S006,W3S016,W3S026,W3S106,W3S116,W3S126,W3S206,W3S216,W3S226;
(*DONT_TOUCH="true"*) wire W3S007,W3S017,W3S027,W3S107,W3S117,W3S127,W3S207,W3S217,W3S227;
(*DONT_TOUCH="true"*) wire W3S008,W3S018,W3S028,W3S108,W3S118,W3S128,W3S208,W3S218,W3S228;
(*DONT_TOUCH="true"*) wire W3S009,W3S019,W3S029,W3S109,W3S119,W3S129,W3S209,W3S219,W3S229;
(*DONT_TOUCH="true"*) wire W3S00A,W3S01A,W3S02A,W3S10A,W3S11A,W3S12A,W3S20A,W3S21A,W3S22A;
(*DONT_TOUCH="true"*) wire W3S00B,W3S01B,W3S02B,W3S10B,W3S11B,W3S12B,W3S20B,W3S21B,W3S22B;
(*DONT_TOUCH="true"*) wire W3S00C,W3S01C,W3S02C,W3S10C,W3S11C,W3S12C,W3S20C,W3S21C,W3S22C;
(*DONT_TOUCH="true"*) wire W3S00D,W3S01D,W3S02D,W3S10D,W3S11D,W3S12D,W3S20D,W3S21D,W3S22D;
(*DONT_TOUCH="true"*) wire W3S00E,W3S01E,W3S02E,W3S10E,W3S11E,W3S12E,W3S20E,W3S21E,W3S22E;
(*DONT_TOUCH="true"*) wire W3S00F,W3S01F,W3S02F,W3S10F,W3S11F,W3S12F,W3S20F,W3S21F,W3S22F;
(*DONT_TOUCH="true"*) wire W3T000,W3T010,W3T020,W3T100,W3T110,W3T120,W3T200,W3T210,W3T220;
(*DONT_TOUCH="true"*) wire W3T001,W3T011,W3T021,W3T101,W3T111,W3T121,W3T201,W3T211,W3T221;
(*DONT_TOUCH="true"*) wire W3T002,W3T012,W3T022,W3T102,W3T112,W3T122,W3T202,W3T212,W3T222;
(*DONT_TOUCH="true"*) wire W3T003,W3T013,W3T023,W3T103,W3T113,W3T123,W3T203,W3T213,W3T223;
(*DONT_TOUCH="true"*) wire W3T004,W3T014,W3T024,W3T104,W3T114,W3T124,W3T204,W3T214,W3T224;
(*DONT_TOUCH="true"*) wire W3T005,W3T015,W3T025,W3T105,W3T115,W3T125,W3T205,W3T215,W3T225;
(*DONT_TOUCH="true"*) wire W3T006,W3T016,W3T026,W3T106,W3T116,W3T126,W3T206,W3T216,W3T226;
(*DONT_TOUCH="true"*) wire W3T007,W3T017,W3T027,W3T107,W3T117,W3T127,W3T207,W3T217,W3T227;
(*DONT_TOUCH="true"*) wire W3T008,W3T018,W3T028,W3T108,W3T118,W3T128,W3T208,W3T218,W3T228;
(*DONT_TOUCH="true"*) wire W3T009,W3T019,W3T029,W3T109,W3T119,W3T129,W3T209,W3T219,W3T229;
(*DONT_TOUCH="true"*) wire W3T00A,W3T01A,W3T02A,W3T10A,W3T11A,W3T12A,W3T20A,W3T21A,W3T22A;
(*DONT_TOUCH="true"*) wire W3T00B,W3T01B,W3T02B,W3T10B,W3T11B,W3T12B,W3T20B,W3T21B,W3T22B;
(*DONT_TOUCH="true"*) wire W3T00C,W3T01C,W3T02C,W3T10C,W3T11C,W3T12C,W3T20C,W3T21C,W3T22C;
(*DONT_TOUCH="true"*) wire W3T00D,W3T01D,W3T02D,W3T10D,W3T11D,W3T12D,W3T20D,W3T21D,W3T22D;
(*DONT_TOUCH="true"*) wire W3T00E,W3T01E,W3T02E,W3T10E,W3T11E,W3T12E,W3T20E,W3T21E,W3T22E;
(*DONT_TOUCH="true"*) wire W3T00F,W3T01F,W3T02F,W3T10F,W3T11F,W3T12F,W3T20F,W3T21F,W3T22F;
(*DONT_TOUCH="true"*) wire W3U000,W3U010,W3U020,W3U100,W3U110,W3U120,W3U200,W3U210,W3U220;
(*DONT_TOUCH="true"*) wire W3U001,W3U011,W3U021,W3U101,W3U111,W3U121,W3U201,W3U211,W3U221;
(*DONT_TOUCH="true"*) wire W3U002,W3U012,W3U022,W3U102,W3U112,W3U122,W3U202,W3U212,W3U222;
(*DONT_TOUCH="true"*) wire W3U003,W3U013,W3U023,W3U103,W3U113,W3U123,W3U203,W3U213,W3U223;
(*DONT_TOUCH="true"*) wire W3U004,W3U014,W3U024,W3U104,W3U114,W3U124,W3U204,W3U214,W3U224;
(*DONT_TOUCH="true"*) wire W3U005,W3U015,W3U025,W3U105,W3U115,W3U125,W3U205,W3U215,W3U225;
(*DONT_TOUCH="true"*) wire W3U006,W3U016,W3U026,W3U106,W3U116,W3U126,W3U206,W3U216,W3U226;
(*DONT_TOUCH="true"*) wire W3U007,W3U017,W3U027,W3U107,W3U117,W3U127,W3U207,W3U217,W3U227;
(*DONT_TOUCH="true"*) wire W3U008,W3U018,W3U028,W3U108,W3U118,W3U128,W3U208,W3U218,W3U228;
(*DONT_TOUCH="true"*) wire W3U009,W3U019,W3U029,W3U109,W3U119,W3U129,W3U209,W3U219,W3U229;
(*DONT_TOUCH="true"*) wire W3U00A,W3U01A,W3U02A,W3U10A,W3U11A,W3U12A,W3U20A,W3U21A,W3U22A;
(*DONT_TOUCH="true"*) wire W3U00B,W3U01B,W3U02B,W3U10B,W3U11B,W3U12B,W3U20B,W3U21B,W3U22B;
(*DONT_TOUCH="true"*) wire W3U00C,W3U01C,W3U02C,W3U10C,W3U11C,W3U12C,W3U20C,W3U21C,W3U22C;
(*DONT_TOUCH="true"*) wire W3U00D,W3U01D,W3U02D,W3U10D,W3U11D,W3U12D,W3U20D,W3U21D,W3U22D;
(*DONT_TOUCH="true"*) wire W3U00E,W3U01E,W3U02E,W3U10E,W3U11E,W3U12E,W3U20E,W3U21E,W3U22E;
(*DONT_TOUCH="true"*) wire W3U00F,W3U01F,W3U02F,W3U10F,W3U11F,W3U12F,W3U20F,W3U21F,W3U22F;
(*DONT_TOUCH="true"*) wire W3V000,W3V010,W3V020,W3V100,W3V110,W3V120,W3V200,W3V210,W3V220;
(*DONT_TOUCH="true"*) wire W3V001,W3V011,W3V021,W3V101,W3V111,W3V121,W3V201,W3V211,W3V221;
(*DONT_TOUCH="true"*) wire W3V002,W3V012,W3V022,W3V102,W3V112,W3V122,W3V202,W3V212,W3V222;
(*DONT_TOUCH="true"*) wire W3V003,W3V013,W3V023,W3V103,W3V113,W3V123,W3V203,W3V213,W3V223;
(*DONT_TOUCH="true"*) wire W3V004,W3V014,W3V024,W3V104,W3V114,W3V124,W3V204,W3V214,W3V224;
(*DONT_TOUCH="true"*) wire W3V005,W3V015,W3V025,W3V105,W3V115,W3V125,W3V205,W3V215,W3V225;
(*DONT_TOUCH="true"*) wire W3V006,W3V016,W3V026,W3V106,W3V116,W3V126,W3V206,W3V216,W3V226;
(*DONT_TOUCH="true"*) wire W3V007,W3V017,W3V027,W3V107,W3V117,W3V127,W3V207,W3V217,W3V227;
(*DONT_TOUCH="true"*) wire W3V008,W3V018,W3V028,W3V108,W3V118,W3V128,W3V208,W3V218,W3V228;
(*DONT_TOUCH="true"*) wire W3V009,W3V019,W3V029,W3V109,W3V119,W3V129,W3V209,W3V219,W3V229;
(*DONT_TOUCH="true"*) wire W3V00A,W3V01A,W3V02A,W3V10A,W3V11A,W3V12A,W3V20A,W3V21A,W3V22A;
(*DONT_TOUCH="true"*) wire W3V00B,W3V01B,W3V02B,W3V10B,W3V11B,W3V12B,W3V20B,W3V21B,W3V22B;
(*DONT_TOUCH="true"*) wire W3V00C,W3V01C,W3V02C,W3V10C,W3V11C,W3V12C,W3V20C,W3V21C,W3V22C;
(*DONT_TOUCH="true"*) wire W3V00D,W3V01D,W3V02D,W3V10D,W3V11D,W3V12D,W3V20D,W3V21D,W3V22D;
(*DONT_TOUCH="true"*) wire W3V00E,W3V01E,W3V02E,W3V10E,W3V11E,W3V12E,W3V20E,W3V21E,W3V22E;
(*DONT_TOUCH="true"*) wire W3V00F,W3V01F,W3V02F,W3V10F,W3V11F,W3V12F,W3V20F,W3V21F,W3V22F;
(*DONT_TOUCH="true"*) wire signed [4:0] c30000,c31000,c32000,c33000,c34000,c35000,c36000,c37000,c38000,c39000,c3A000,c3B000,c3C000,c3D000,c3E000,c3F000;
(*DONT_TOUCH="true"*) wire signed [4:0] c30010,c31010,c32010,c33010,c34010,c35010,c36010,c37010,c38010,c39010,c3A010,c3B010,c3C010,c3D010,c3E010,c3F010;
(*DONT_TOUCH="true"*) wire signed [4:0] c30020,c31020,c32020,c33020,c34020,c35020,c36020,c37020,c38020,c39020,c3A020,c3B020,c3C020,c3D020,c3E020,c3F020;
(*DONT_TOUCH="true"*) wire signed [4:0] c30100,c31100,c32100,c33100,c34100,c35100,c36100,c37100,c38100,c39100,c3A100,c3B100,c3C100,c3D100,c3E100,c3F100;
(*DONT_TOUCH="true"*) wire signed [4:0] c30110,c31110,c32110,c33110,c34110,c35110,c36110,c37110,c38110,c39110,c3A110,c3B110,c3C110,c3D110,c3E110,c3F110;
(*DONT_TOUCH="true"*) wire signed [4:0] c30120,c31120,c32120,c33120,c34120,c35120,c36120,c37120,c38120,c39120,c3A120,c3B120,c3C120,c3D120,c3E120,c3F120;
(*DONT_TOUCH="true"*) wire signed [4:0] c30200,c31200,c32200,c33200,c34200,c35200,c36200,c37200,c38200,c39200,c3A200,c3B200,c3C200,c3D200,c3E200,c3F200;
(*DONT_TOUCH="true"*) wire signed [4:0] c30210,c31210,c32210,c33210,c34210,c35210,c36210,c37210,c38210,c39210,c3A210,c3B210,c3C210,c3D210,c3E210,c3F210;
(*DONT_TOUCH="true"*) wire signed [4:0] c30220,c31220,c32220,c33220,c34220,c35220,c36220,c37220,c38220,c39220,c3A220,c3B220,c3C220,c3D220,c3E220,c3F220;
(*DONT_TOUCH="true"*) wire signed [4:0] c30001,c31001,c32001,c33001,c34001,c35001,c36001,c37001,c38001,c39001,c3A001,c3B001,c3C001,c3D001,c3E001,c3F001;
(*DONT_TOUCH="true"*) wire signed [4:0] c30011,c31011,c32011,c33011,c34011,c35011,c36011,c37011,c38011,c39011,c3A011,c3B011,c3C011,c3D011,c3E011,c3F011;
(*DONT_TOUCH="true"*) wire signed [4:0] c30021,c31021,c32021,c33021,c34021,c35021,c36021,c37021,c38021,c39021,c3A021,c3B021,c3C021,c3D021,c3E021,c3F021;
(*DONT_TOUCH="true"*) wire signed [4:0] c30101,c31101,c32101,c33101,c34101,c35101,c36101,c37101,c38101,c39101,c3A101,c3B101,c3C101,c3D101,c3E101,c3F101;
(*DONT_TOUCH="true"*) wire signed [4:0] c30111,c31111,c32111,c33111,c34111,c35111,c36111,c37111,c38111,c39111,c3A111,c3B111,c3C111,c3D111,c3E111,c3F111;
(*DONT_TOUCH="true"*) wire signed [4:0] c30121,c31121,c32121,c33121,c34121,c35121,c36121,c37121,c38121,c39121,c3A121,c3B121,c3C121,c3D121,c3E121,c3F121;
(*DONT_TOUCH="true"*) wire signed [4:0] c30201,c31201,c32201,c33201,c34201,c35201,c36201,c37201,c38201,c39201,c3A201,c3B201,c3C201,c3D201,c3E201,c3F201;
(*DONT_TOUCH="true"*) wire signed [4:0] c30211,c31211,c32211,c33211,c34211,c35211,c36211,c37211,c38211,c39211,c3A211,c3B211,c3C211,c3D211,c3E211,c3F211;
(*DONT_TOUCH="true"*) wire signed [4:0] c30221,c31221,c32221,c33221,c34221,c35221,c36221,c37221,c38221,c39221,c3A221,c3B221,c3C221,c3D221,c3E221,c3F221;
(*DONT_TOUCH="true"*) wire signed [4:0] c30002,c31002,c32002,c33002,c34002,c35002,c36002,c37002,c38002,c39002,c3A002,c3B002,c3C002,c3D002,c3E002,c3F002;
(*DONT_TOUCH="true"*) wire signed [4:0] c30012,c31012,c32012,c33012,c34012,c35012,c36012,c37012,c38012,c39012,c3A012,c3B012,c3C012,c3D012,c3E012,c3F012;
(*DONT_TOUCH="true"*) wire signed [4:0] c30022,c31022,c32022,c33022,c34022,c35022,c36022,c37022,c38022,c39022,c3A022,c3B022,c3C022,c3D022,c3E022,c3F022;
(*DONT_TOUCH="true"*) wire signed [4:0] c30102,c31102,c32102,c33102,c34102,c35102,c36102,c37102,c38102,c39102,c3A102,c3B102,c3C102,c3D102,c3E102,c3F102;
(*DONT_TOUCH="true"*) wire signed [4:0] c30112,c31112,c32112,c33112,c34112,c35112,c36112,c37112,c38112,c39112,c3A112,c3B112,c3C112,c3D112,c3E112,c3F112;
(*DONT_TOUCH="true"*) wire signed [4:0] c30122,c31122,c32122,c33122,c34122,c35122,c36122,c37122,c38122,c39122,c3A122,c3B122,c3C122,c3D122,c3E122,c3F122;
(*DONT_TOUCH="true"*) wire signed [4:0] c30202,c31202,c32202,c33202,c34202,c35202,c36202,c37202,c38202,c39202,c3A202,c3B202,c3C202,c3D202,c3E202,c3F202;
(*DONT_TOUCH="true"*) wire signed [4:0] c30212,c31212,c32212,c33212,c34212,c35212,c36212,c37212,c38212,c39212,c3A212,c3B212,c3C212,c3D212,c3E212,c3F212;
(*DONT_TOUCH="true"*) wire signed [4:0] c30222,c31222,c32222,c33222,c34222,c35222,c36222,c37222,c38222,c39222,c3A222,c3B222,c3C222,c3D222,c3E222,c3F222;
(*DONT_TOUCH="true"*) wire signed [4:0] c30003,c31003,c32003,c33003,c34003,c35003,c36003,c37003,c38003,c39003,c3A003,c3B003,c3C003,c3D003,c3E003,c3F003;
(*DONT_TOUCH="true"*) wire signed [4:0] c30013,c31013,c32013,c33013,c34013,c35013,c36013,c37013,c38013,c39013,c3A013,c3B013,c3C013,c3D013,c3E013,c3F013;
(*DONT_TOUCH="true"*) wire signed [4:0] c30023,c31023,c32023,c33023,c34023,c35023,c36023,c37023,c38023,c39023,c3A023,c3B023,c3C023,c3D023,c3E023,c3F023;
(*DONT_TOUCH="true"*) wire signed [4:0] c30103,c31103,c32103,c33103,c34103,c35103,c36103,c37103,c38103,c39103,c3A103,c3B103,c3C103,c3D103,c3E103,c3F103;
(*DONT_TOUCH="true"*) wire signed [4:0] c30113,c31113,c32113,c33113,c34113,c35113,c36113,c37113,c38113,c39113,c3A113,c3B113,c3C113,c3D113,c3E113,c3F113;
(*DONT_TOUCH="true"*) wire signed [4:0] c30123,c31123,c32123,c33123,c34123,c35123,c36123,c37123,c38123,c39123,c3A123,c3B123,c3C123,c3D123,c3E123,c3F123;
(*DONT_TOUCH="true"*) wire signed [4:0] c30203,c31203,c32203,c33203,c34203,c35203,c36203,c37203,c38203,c39203,c3A203,c3B203,c3C203,c3D203,c3E203,c3F203;
(*DONT_TOUCH="true"*) wire signed [4:0] c30213,c31213,c32213,c33213,c34213,c35213,c36213,c37213,c38213,c39213,c3A213,c3B213,c3C213,c3D213,c3E213,c3F213;
(*DONT_TOUCH="true"*) wire signed [4:0] c30223,c31223,c32223,c33223,c34223,c35223,c36223,c37223,c38223,c39223,c3A223,c3B223,c3C223,c3D223,c3E223,c3F223;
(*DONT_TOUCH="true"*) wire signed [4:0] c30004,c31004,c32004,c33004,c34004,c35004,c36004,c37004,c38004,c39004,c3A004,c3B004,c3C004,c3D004,c3E004,c3F004;
(*DONT_TOUCH="true"*) wire signed [4:0] c30014,c31014,c32014,c33014,c34014,c35014,c36014,c37014,c38014,c39014,c3A014,c3B014,c3C014,c3D014,c3E014,c3F014;
(*DONT_TOUCH="true"*) wire signed [4:0] c30024,c31024,c32024,c33024,c34024,c35024,c36024,c37024,c38024,c39024,c3A024,c3B024,c3C024,c3D024,c3E024,c3F024;
(*DONT_TOUCH="true"*) wire signed [4:0] c30104,c31104,c32104,c33104,c34104,c35104,c36104,c37104,c38104,c39104,c3A104,c3B104,c3C104,c3D104,c3E104,c3F104;
(*DONT_TOUCH="true"*) wire signed [4:0] c30114,c31114,c32114,c33114,c34114,c35114,c36114,c37114,c38114,c39114,c3A114,c3B114,c3C114,c3D114,c3E114,c3F114;
(*DONT_TOUCH="true"*) wire signed [4:0] c30124,c31124,c32124,c33124,c34124,c35124,c36124,c37124,c38124,c39124,c3A124,c3B124,c3C124,c3D124,c3E124,c3F124;
(*DONT_TOUCH="true"*) wire signed [4:0] c30204,c31204,c32204,c33204,c34204,c35204,c36204,c37204,c38204,c39204,c3A204,c3B204,c3C204,c3D204,c3E204,c3F204;
(*DONT_TOUCH="true"*) wire signed [4:0] c30214,c31214,c32214,c33214,c34214,c35214,c36214,c37214,c38214,c39214,c3A214,c3B214,c3C214,c3D214,c3E214,c3F214;
(*DONT_TOUCH="true"*) wire signed [4:0] c30224,c31224,c32224,c33224,c34224,c35224,c36224,c37224,c38224,c39224,c3A224,c3B224,c3C224,c3D224,c3E224,c3F224;
(*DONT_TOUCH="true"*) wire signed [4:0] c30005,c31005,c32005,c33005,c34005,c35005,c36005,c37005,c38005,c39005,c3A005,c3B005,c3C005,c3D005,c3E005,c3F005;
(*DONT_TOUCH="true"*) wire signed [4:0] c30015,c31015,c32015,c33015,c34015,c35015,c36015,c37015,c38015,c39015,c3A015,c3B015,c3C015,c3D015,c3E015,c3F015;
(*DONT_TOUCH="true"*) wire signed [4:0] c30025,c31025,c32025,c33025,c34025,c35025,c36025,c37025,c38025,c39025,c3A025,c3B025,c3C025,c3D025,c3E025,c3F025;
(*DONT_TOUCH="true"*) wire signed [4:0] c30105,c31105,c32105,c33105,c34105,c35105,c36105,c37105,c38105,c39105,c3A105,c3B105,c3C105,c3D105,c3E105,c3F105;
(*DONT_TOUCH="true"*) wire signed [4:0] c30115,c31115,c32115,c33115,c34115,c35115,c36115,c37115,c38115,c39115,c3A115,c3B115,c3C115,c3D115,c3E115,c3F115;
(*DONT_TOUCH="true"*) wire signed [4:0] c30125,c31125,c32125,c33125,c34125,c35125,c36125,c37125,c38125,c39125,c3A125,c3B125,c3C125,c3D125,c3E125,c3F125;
(*DONT_TOUCH="true"*) wire signed [4:0] c30205,c31205,c32205,c33205,c34205,c35205,c36205,c37205,c38205,c39205,c3A205,c3B205,c3C205,c3D205,c3E205,c3F205;
(*DONT_TOUCH="true"*) wire signed [4:0] c30215,c31215,c32215,c33215,c34215,c35215,c36215,c37215,c38215,c39215,c3A215,c3B215,c3C215,c3D215,c3E215,c3F215;
(*DONT_TOUCH="true"*) wire signed [4:0] c30225,c31225,c32225,c33225,c34225,c35225,c36225,c37225,c38225,c39225,c3A225,c3B225,c3C225,c3D225,c3E225,c3F225;
(*DONT_TOUCH="true"*) wire signed [4:0] c30006,c31006,c32006,c33006,c34006,c35006,c36006,c37006,c38006,c39006,c3A006,c3B006,c3C006,c3D006,c3E006,c3F006;
(*DONT_TOUCH="true"*) wire signed [4:0] c30016,c31016,c32016,c33016,c34016,c35016,c36016,c37016,c38016,c39016,c3A016,c3B016,c3C016,c3D016,c3E016,c3F016;
(*DONT_TOUCH="true"*) wire signed [4:0] c30026,c31026,c32026,c33026,c34026,c35026,c36026,c37026,c38026,c39026,c3A026,c3B026,c3C026,c3D026,c3E026,c3F026;
(*DONT_TOUCH="true"*) wire signed [4:0] c30106,c31106,c32106,c33106,c34106,c35106,c36106,c37106,c38106,c39106,c3A106,c3B106,c3C106,c3D106,c3E106,c3F106;
(*DONT_TOUCH="true"*) wire signed [4:0] c30116,c31116,c32116,c33116,c34116,c35116,c36116,c37116,c38116,c39116,c3A116,c3B116,c3C116,c3D116,c3E116,c3F116;
(*DONT_TOUCH="true"*) wire signed [4:0] c30126,c31126,c32126,c33126,c34126,c35126,c36126,c37126,c38126,c39126,c3A126,c3B126,c3C126,c3D126,c3E126,c3F126;
(*DONT_TOUCH="true"*) wire signed [4:0] c30206,c31206,c32206,c33206,c34206,c35206,c36206,c37206,c38206,c39206,c3A206,c3B206,c3C206,c3D206,c3E206,c3F206;
(*DONT_TOUCH="true"*) wire signed [4:0] c30216,c31216,c32216,c33216,c34216,c35216,c36216,c37216,c38216,c39216,c3A216,c3B216,c3C216,c3D216,c3E216,c3F216;
(*DONT_TOUCH="true"*) wire signed [4:0] c30226,c31226,c32226,c33226,c34226,c35226,c36226,c37226,c38226,c39226,c3A226,c3B226,c3C226,c3D226,c3E226,c3F226;
(*DONT_TOUCH="true"*) wire signed [4:0] c30007,c31007,c32007,c33007,c34007,c35007,c36007,c37007,c38007,c39007,c3A007,c3B007,c3C007,c3D007,c3E007,c3F007;
(*DONT_TOUCH="true"*) wire signed [4:0] c30017,c31017,c32017,c33017,c34017,c35017,c36017,c37017,c38017,c39017,c3A017,c3B017,c3C017,c3D017,c3E017,c3F017;
(*DONT_TOUCH="true"*) wire signed [4:0] c30027,c31027,c32027,c33027,c34027,c35027,c36027,c37027,c38027,c39027,c3A027,c3B027,c3C027,c3D027,c3E027,c3F027;
(*DONT_TOUCH="true"*) wire signed [4:0] c30107,c31107,c32107,c33107,c34107,c35107,c36107,c37107,c38107,c39107,c3A107,c3B107,c3C107,c3D107,c3E107,c3F107;
(*DONT_TOUCH="true"*) wire signed [4:0] c30117,c31117,c32117,c33117,c34117,c35117,c36117,c37117,c38117,c39117,c3A117,c3B117,c3C117,c3D117,c3E117,c3F117;
(*DONT_TOUCH="true"*) wire signed [4:0] c30127,c31127,c32127,c33127,c34127,c35127,c36127,c37127,c38127,c39127,c3A127,c3B127,c3C127,c3D127,c3E127,c3F127;
(*DONT_TOUCH="true"*) wire signed [4:0] c30207,c31207,c32207,c33207,c34207,c35207,c36207,c37207,c38207,c39207,c3A207,c3B207,c3C207,c3D207,c3E207,c3F207;
(*DONT_TOUCH="true"*) wire signed [4:0] c30217,c31217,c32217,c33217,c34217,c35217,c36217,c37217,c38217,c39217,c3A217,c3B217,c3C217,c3D217,c3E217,c3F217;
(*DONT_TOUCH="true"*) wire signed [4:0] c30227,c31227,c32227,c33227,c34227,c35227,c36227,c37227,c38227,c39227,c3A227,c3B227,c3C227,c3D227,c3E227,c3F227;
(*DONT_TOUCH="true"*) wire signed [4:0] c30008,c31008,c32008,c33008,c34008,c35008,c36008,c37008,c38008,c39008,c3A008,c3B008,c3C008,c3D008,c3E008,c3F008;
(*DONT_TOUCH="true"*) wire signed [4:0] c30018,c31018,c32018,c33018,c34018,c35018,c36018,c37018,c38018,c39018,c3A018,c3B018,c3C018,c3D018,c3E018,c3F018;
(*DONT_TOUCH="true"*) wire signed [4:0] c30028,c31028,c32028,c33028,c34028,c35028,c36028,c37028,c38028,c39028,c3A028,c3B028,c3C028,c3D028,c3E028,c3F028;
(*DONT_TOUCH="true"*) wire signed [4:0] c30108,c31108,c32108,c33108,c34108,c35108,c36108,c37108,c38108,c39108,c3A108,c3B108,c3C108,c3D108,c3E108,c3F108;
(*DONT_TOUCH="true"*) wire signed [4:0] c30118,c31118,c32118,c33118,c34118,c35118,c36118,c37118,c38118,c39118,c3A118,c3B118,c3C118,c3D118,c3E118,c3F118;
(*DONT_TOUCH="true"*) wire signed [4:0] c30128,c31128,c32128,c33128,c34128,c35128,c36128,c37128,c38128,c39128,c3A128,c3B128,c3C128,c3D128,c3E128,c3F128;
(*DONT_TOUCH="true"*) wire signed [4:0] c30208,c31208,c32208,c33208,c34208,c35208,c36208,c37208,c38208,c39208,c3A208,c3B208,c3C208,c3D208,c3E208,c3F208;
(*DONT_TOUCH="true"*) wire signed [4:0] c30218,c31218,c32218,c33218,c34218,c35218,c36218,c37218,c38218,c39218,c3A218,c3B218,c3C218,c3D218,c3E218,c3F218;
(*DONT_TOUCH="true"*) wire signed [4:0] c30228,c31228,c32228,c33228,c34228,c35228,c36228,c37228,c38228,c39228,c3A228,c3B228,c3C228,c3D228,c3E228,c3F228;
(*DONT_TOUCH="true"*) wire signed [4:0] c30009,c31009,c32009,c33009,c34009,c35009,c36009,c37009,c38009,c39009,c3A009,c3B009,c3C009,c3D009,c3E009,c3F009;
(*DONT_TOUCH="true"*) wire signed [4:0] c30019,c31019,c32019,c33019,c34019,c35019,c36019,c37019,c38019,c39019,c3A019,c3B019,c3C019,c3D019,c3E019,c3F019;
(*DONT_TOUCH="true"*) wire signed [4:0] c30029,c31029,c32029,c33029,c34029,c35029,c36029,c37029,c38029,c39029,c3A029,c3B029,c3C029,c3D029,c3E029,c3F029;
(*DONT_TOUCH="true"*) wire signed [4:0] c30109,c31109,c32109,c33109,c34109,c35109,c36109,c37109,c38109,c39109,c3A109,c3B109,c3C109,c3D109,c3E109,c3F109;
(*DONT_TOUCH="true"*) wire signed [4:0] c30119,c31119,c32119,c33119,c34119,c35119,c36119,c37119,c38119,c39119,c3A119,c3B119,c3C119,c3D119,c3E119,c3F119;
(*DONT_TOUCH="true"*) wire signed [4:0] c30129,c31129,c32129,c33129,c34129,c35129,c36129,c37129,c38129,c39129,c3A129,c3B129,c3C129,c3D129,c3E129,c3F129;
(*DONT_TOUCH="true"*) wire signed [4:0] c30209,c31209,c32209,c33209,c34209,c35209,c36209,c37209,c38209,c39209,c3A209,c3B209,c3C209,c3D209,c3E209,c3F209;
(*DONT_TOUCH="true"*) wire signed [4:0] c30219,c31219,c32219,c33219,c34219,c35219,c36219,c37219,c38219,c39219,c3A219,c3B219,c3C219,c3D219,c3E219,c3F219;
(*DONT_TOUCH="true"*) wire signed [4:0] c30229,c31229,c32229,c33229,c34229,c35229,c36229,c37229,c38229,c39229,c3A229,c3B229,c3C229,c3D229,c3E229,c3F229;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000A,c3100A,c3200A,c3300A,c3400A,c3500A,c3600A,c3700A,c3800A,c3900A,c3A00A,c3B00A,c3C00A,c3D00A,c3E00A,c3F00A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001A,c3101A,c3201A,c3301A,c3401A,c3501A,c3601A,c3701A,c3801A,c3901A,c3A01A,c3B01A,c3C01A,c3D01A,c3E01A,c3F01A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002A,c3102A,c3202A,c3302A,c3402A,c3502A,c3602A,c3702A,c3802A,c3902A,c3A02A,c3B02A,c3C02A,c3D02A,c3E02A,c3F02A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010A,c3110A,c3210A,c3310A,c3410A,c3510A,c3610A,c3710A,c3810A,c3910A,c3A10A,c3B10A,c3C10A,c3D10A,c3E10A,c3F10A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011A,c3111A,c3211A,c3311A,c3411A,c3511A,c3611A,c3711A,c3811A,c3911A,c3A11A,c3B11A,c3C11A,c3D11A,c3E11A,c3F11A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012A,c3112A,c3212A,c3312A,c3412A,c3512A,c3612A,c3712A,c3812A,c3912A,c3A12A,c3B12A,c3C12A,c3D12A,c3E12A,c3F12A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020A,c3120A,c3220A,c3320A,c3420A,c3520A,c3620A,c3720A,c3820A,c3920A,c3A20A,c3B20A,c3C20A,c3D20A,c3E20A,c3F20A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021A,c3121A,c3221A,c3321A,c3421A,c3521A,c3621A,c3721A,c3821A,c3921A,c3A21A,c3B21A,c3C21A,c3D21A,c3E21A,c3F21A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022A,c3122A,c3222A,c3322A,c3422A,c3522A,c3622A,c3722A,c3822A,c3922A,c3A22A,c3B22A,c3C22A,c3D22A,c3E22A,c3F22A;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000B,c3100B,c3200B,c3300B,c3400B,c3500B,c3600B,c3700B,c3800B,c3900B,c3A00B,c3B00B,c3C00B,c3D00B,c3E00B,c3F00B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001B,c3101B,c3201B,c3301B,c3401B,c3501B,c3601B,c3701B,c3801B,c3901B,c3A01B,c3B01B,c3C01B,c3D01B,c3E01B,c3F01B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002B,c3102B,c3202B,c3302B,c3402B,c3502B,c3602B,c3702B,c3802B,c3902B,c3A02B,c3B02B,c3C02B,c3D02B,c3E02B,c3F02B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010B,c3110B,c3210B,c3310B,c3410B,c3510B,c3610B,c3710B,c3810B,c3910B,c3A10B,c3B10B,c3C10B,c3D10B,c3E10B,c3F10B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011B,c3111B,c3211B,c3311B,c3411B,c3511B,c3611B,c3711B,c3811B,c3911B,c3A11B,c3B11B,c3C11B,c3D11B,c3E11B,c3F11B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012B,c3112B,c3212B,c3312B,c3412B,c3512B,c3612B,c3712B,c3812B,c3912B,c3A12B,c3B12B,c3C12B,c3D12B,c3E12B,c3F12B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020B,c3120B,c3220B,c3320B,c3420B,c3520B,c3620B,c3720B,c3820B,c3920B,c3A20B,c3B20B,c3C20B,c3D20B,c3E20B,c3F20B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021B,c3121B,c3221B,c3321B,c3421B,c3521B,c3621B,c3721B,c3821B,c3921B,c3A21B,c3B21B,c3C21B,c3D21B,c3E21B,c3F21B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022B,c3122B,c3222B,c3322B,c3422B,c3522B,c3622B,c3722B,c3822B,c3922B,c3A22B,c3B22B,c3C22B,c3D22B,c3E22B,c3F22B;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000C,c3100C,c3200C,c3300C,c3400C,c3500C,c3600C,c3700C,c3800C,c3900C,c3A00C,c3B00C,c3C00C,c3D00C,c3E00C,c3F00C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001C,c3101C,c3201C,c3301C,c3401C,c3501C,c3601C,c3701C,c3801C,c3901C,c3A01C,c3B01C,c3C01C,c3D01C,c3E01C,c3F01C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002C,c3102C,c3202C,c3302C,c3402C,c3502C,c3602C,c3702C,c3802C,c3902C,c3A02C,c3B02C,c3C02C,c3D02C,c3E02C,c3F02C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010C,c3110C,c3210C,c3310C,c3410C,c3510C,c3610C,c3710C,c3810C,c3910C,c3A10C,c3B10C,c3C10C,c3D10C,c3E10C,c3F10C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011C,c3111C,c3211C,c3311C,c3411C,c3511C,c3611C,c3711C,c3811C,c3911C,c3A11C,c3B11C,c3C11C,c3D11C,c3E11C,c3F11C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012C,c3112C,c3212C,c3312C,c3412C,c3512C,c3612C,c3712C,c3812C,c3912C,c3A12C,c3B12C,c3C12C,c3D12C,c3E12C,c3F12C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020C,c3120C,c3220C,c3320C,c3420C,c3520C,c3620C,c3720C,c3820C,c3920C,c3A20C,c3B20C,c3C20C,c3D20C,c3E20C,c3F20C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021C,c3121C,c3221C,c3321C,c3421C,c3521C,c3621C,c3721C,c3821C,c3921C,c3A21C,c3B21C,c3C21C,c3D21C,c3E21C,c3F21C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022C,c3122C,c3222C,c3322C,c3422C,c3522C,c3622C,c3722C,c3822C,c3922C,c3A22C,c3B22C,c3C22C,c3D22C,c3E22C,c3F22C;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000D,c3100D,c3200D,c3300D,c3400D,c3500D,c3600D,c3700D,c3800D,c3900D,c3A00D,c3B00D,c3C00D,c3D00D,c3E00D,c3F00D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001D,c3101D,c3201D,c3301D,c3401D,c3501D,c3601D,c3701D,c3801D,c3901D,c3A01D,c3B01D,c3C01D,c3D01D,c3E01D,c3F01D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002D,c3102D,c3202D,c3302D,c3402D,c3502D,c3602D,c3702D,c3802D,c3902D,c3A02D,c3B02D,c3C02D,c3D02D,c3E02D,c3F02D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010D,c3110D,c3210D,c3310D,c3410D,c3510D,c3610D,c3710D,c3810D,c3910D,c3A10D,c3B10D,c3C10D,c3D10D,c3E10D,c3F10D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011D,c3111D,c3211D,c3311D,c3411D,c3511D,c3611D,c3711D,c3811D,c3911D,c3A11D,c3B11D,c3C11D,c3D11D,c3E11D,c3F11D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012D,c3112D,c3212D,c3312D,c3412D,c3512D,c3612D,c3712D,c3812D,c3912D,c3A12D,c3B12D,c3C12D,c3D12D,c3E12D,c3F12D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020D,c3120D,c3220D,c3320D,c3420D,c3520D,c3620D,c3720D,c3820D,c3920D,c3A20D,c3B20D,c3C20D,c3D20D,c3E20D,c3F20D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021D,c3121D,c3221D,c3321D,c3421D,c3521D,c3621D,c3721D,c3821D,c3921D,c3A21D,c3B21D,c3C21D,c3D21D,c3E21D,c3F21D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022D,c3122D,c3222D,c3322D,c3422D,c3522D,c3622D,c3722D,c3822D,c3922D,c3A22D,c3B22D,c3C22D,c3D22D,c3E22D,c3F22D;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000E,c3100E,c3200E,c3300E,c3400E,c3500E,c3600E,c3700E,c3800E,c3900E,c3A00E,c3B00E,c3C00E,c3D00E,c3E00E,c3F00E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001E,c3101E,c3201E,c3301E,c3401E,c3501E,c3601E,c3701E,c3801E,c3901E,c3A01E,c3B01E,c3C01E,c3D01E,c3E01E,c3F01E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002E,c3102E,c3202E,c3302E,c3402E,c3502E,c3602E,c3702E,c3802E,c3902E,c3A02E,c3B02E,c3C02E,c3D02E,c3E02E,c3F02E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010E,c3110E,c3210E,c3310E,c3410E,c3510E,c3610E,c3710E,c3810E,c3910E,c3A10E,c3B10E,c3C10E,c3D10E,c3E10E,c3F10E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011E,c3111E,c3211E,c3311E,c3411E,c3511E,c3611E,c3711E,c3811E,c3911E,c3A11E,c3B11E,c3C11E,c3D11E,c3E11E,c3F11E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012E,c3112E,c3212E,c3312E,c3412E,c3512E,c3612E,c3712E,c3812E,c3912E,c3A12E,c3B12E,c3C12E,c3D12E,c3E12E,c3F12E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020E,c3120E,c3220E,c3320E,c3420E,c3520E,c3620E,c3720E,c3820E,c3920E,c3A20E,c3B20E,c3C20E,c3D20E,c3E20E,c3F20E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021E,c3121E,c3221E,c3321E,c3421E,c3521E,c3621E,c3721E,c3821E,c3921E,c3A21E,c3B21E,c3C21E,c3D21E,c3E21E,c3F21E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022E,c3122E,c3222E,c3322E,c3422E,c3522E,c3622E,c3722E,c3822E,c3922E,c3A22E,c3B22E,c3C22E,c3D22E,c3E22E,c3F22E;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000F,c3100F,c3200F,c3300F,c3400F,c3500F,c3600F,c3700F,c3800F,c3900F,c3A00F,c3B00F,c3C00F,c3D00F,c3E00F,c3F00F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001F,c3101F,c3201F,c3301F,c3401F,c3501F,c3601F,c3701F,c3801F,c3901F,c3A01F,c3B01F,c3C01F,c3D01F,c3E01F,c3F01F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002F,c3102F,c3202F,c3302F,c3402F,c3502F,c3602F,c3702F,c3802F,c3902F,c3A02F,c3B02F,c3C02F,c3D02F,c3E02F,c3F02F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010F,c3110F,c3210F,c3310F,c3410F,c3510F,c3610F,c3710F,c3810F,c3910F,c3A10F,c3B10F,c3C10F,c3D10F,c3E10F,c3F10F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011F,c3111F,c3211F,c3311F,c3411F,c3511F,c3611F,c3711F,c3811F,c3911F,c3A11F,c3B11F,c3C11F,c3D11F,c3E11F,c3F11F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012F,c3112F,c3212F,c3312F,c3412F,c3512F,c3612F,c3712F,c3812F,c3912F,c3A12F,c3B12F,c3C12F,c3D12F,c3E12F,c3F12F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020F,c3120F,c3220F,c3320F,c3420F,c3520F,c3620F,c3720F,c3820F,c3920F,c3A20F,c3B20F,c3C20F,c3D20F,c3E20F,c3F20F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021F,c3121F,c3221F,c3321F,c3421F,c3521F,c3621F,c3721F,c3821F,c3921F,c3A21F,c3B21F,c3C21F,c3D21F,c3E21F,c3F21F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022F,c3122F,c3222F,c3322F,c3422F,c3522F,c3622F,c3722F,c3822F,c3922F,c3A22F,c3B22F,c3C22F,c3D22F,c3E22F,c3F22F;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000G,c3100G,c3200G,c3300G,c3400G,c3500G,c3600G,c3700G,c3800G,c3900G,c3A00G,c3B00G,c3C00G,c3D00G,c3E00G,c3F00G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001G,c3101G,c3201G,c3301G,c3401G,c3501G,c3601G,c3701G,c3801G,c3901G,c3A01G,c3B01G,c3C01G,c3D01G,c3E01G,c3F01G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002G,c3102G,c3202G,c3302G,c3402G,c3502G,c3602G,c3702G,c3802G,c3902G,c3A02G,c3B02G,c3C02G,c3D02G,c3E02G,c3F02G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010G,c3110G,c3210G,c3310G,c3410G,c3510G,c3610G,c3710G,c3810G,c3910G,c3A10G,c3B10G,c3C10G,c3D10G,c3E10G,c3F10G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011G,c3111G,c3211G,c3311G,c3411G,c3511G,c3611G,c3711G,c3811G,c3911G,c3A11G,c3B11G,c3C11G,c3D11G,c3E11G,c3F11G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012G,c3112G,c3212G,c3312G,c3412G,c3512G,c3612G,c3712G,c3812G,c3912G,c3A12G,c3B12G,c3C12G,c3D12G,c3E12G,c3F12G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020G,c3120G,c3220G,c3320G,c3420G,c3520G,c3620G,c3720G,c3820G,c3920G,c3A20G,c3B20G,c3C20G,c3D20G,c3E20G,c3F20G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021G,c3121G,c3221G,c3321G,c3421G,c3521G,c3621G,c3721G,c3821G,c3921G,c3A21G,c3B21G,c3C21G,c3D21G,c3E21G,c3F21G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022G,c3122G,c3222G,c3322G,c3422G,c3522G,c3622G,c3722G,c3822G,c3922G,c3A22G,c3B22G,c3C22G,c3D22G,c3E22G,c3F22G;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000H,c3100H,c3200H,c3300H,c3400H,c3500H,c3600H,c3700H,c3800H,c3900H,c3A00H,c3B00H,c3C00H,c3D00H,c3E00H,c3F00H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001H,c3101H,c3201H,c3301H,c3401H,c3501H,c3601H,c3701H,c3801H,c3901H,c3A01H,c3B01H,c3C01H,c3D01H,c3E01H,c3F01H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002H,c3102H,c3202H,c3302H,c3402H,c3502H,c3602H,c3702H,c3802H,c3902H,c3A02H,c3B02H,c3C02H,c3D02H,c3E02H,c3F02H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010H,c3110H,c3210H,c3310H,c3410H,c3510H,c3610H,c3710H,c3810H,c3910H,c3A10H,c3B10H,c3C10H,c3D10H,c3E10H,c3F10H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011H,c3111H,c3211H,c3311H,c3411H,c3511H,c3611H,c3711H,c3811H,c3911H,c3A11H,c3B11H,c3C11H,c3D11H,c3E11H,c3F11H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012H,c3112H,c3212H,c3312H,c3412H,c3512H,c3612H,c3712H,c3812H,c3912H,c3A12H,c3B12H,c3C12H,c3D12H,c3E12H,c3F12H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020H,c3120H,c3220H,c3320H,c3420H,c3520H,c3620H,c3720H,c3820H,c3920H,c3A20H,c3B20H,c3C20H,c3D20H,c3E20H,c3F20H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021H,c3121H,c3221H,c3321H,c3421H,c3521H,c3621H,c3721H,c3821H,c3921H,c3A21H,c3B21H,c3C21H,c3D21H,c3E21H,c3F21H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022H,c3122H,c3222H,c3322H,c3422H,c3522H,c3622H,c3722H,c3822H,c3922H,c3A22H,c3B22H,c3C22H,c3D22H,c3E22H,c3F22H;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000I,c3100I,c3200I,c3300I,c3400I,c3500I,c3600I,c3700I,c3800I,c3900I,c3A00I,c3B00I,c3C00I,c3D00I,c3E00I,c3F00I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001I,c3101I,c3201I,c3301I,c3401I,c3501I,c3601I,c3701I,c3801I,c3901I,c3A01I,c3B01I,c3C01I,c3D01I,c3E01I,c3F01I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002I,c3102I,c3202I,c3302I,c3402I,c3502I,c3602I,c3702I,c3802I,c3902I,c3A02I,c3B02I,c3C02I,c3D02I,c3E02I,c3F02I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010I,c3110I,c3210I,c3310I,c3410I,c3510I,c3610I,c3710I,c3810I,c3910I,c3A10I,c3B10I,c3C10I,c3D10I,c3E10I,c3F10I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011I,c3111I,c3211I,c3311I,c3411I,c3511I,c3611I,c3711I,c3811I,c3911I,c3A11I,c3B11I,c3C11I,c3D11I,c3E11I,c3F11I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012I,c3112I,c3212I,c3312I,c3412I,c3512I,c3612I,c3712I,c3812I,c3912I,c3A12I,c3B12I,c3C12I,c3D12I,c3E12I,c3F12I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020I,c3120I,c3220I,c3320I,c3420I,c3520I,c3620I,c3720I,c3820I,c3920I,c3A20I,c3B20I,c3C20I,c3D20I,c3E20I,c3F20I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021I,c3121I,c3221I,c3321I,c3421I,c3521I,c3621I,c3721I,c3821I,c3921I,c3A21I,c3B21I,c3C21I,c3D21I,c3E21I,c3F21I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022I,c3122I,c3222I,c3322I,c3422I,c3522I,c3622I,c3722I,c3822I,c3922I,c3A22I,c3B22I,c3C22I,c3D22I,c3E22I,c3F22I;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000J,c3100J,c3200J,c3300J,c3400J,c3500J,c3600J,c3700J,c3800J,c3900J,c3A00J,c3B00J,c3C00J,c3D00J,c3E00J,c3F00J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001J,c3101J,c3201J,c3301J,c3401J,c3501J,c3601J,c3701J,c3801J,c3901J,c3A01J,c3B01J,c3C01J,c3D01J,c3E01J,c3F01J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002J,c3102J,c3202J,c3302J,c3402J,c3502J,c3602J,c3702J,c3802J,c3902J,c3A02J,c3B02J,c3C02J,c3D02J,c3E02J,c3F02J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010J,c3110J,c3210J,c3310J,c3410J,c3510J,c3610J,c3710J,c3810J,c3910J,c3A10J,c3B10J,c3C10J,c3D10J,c3E10J,c3F10J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011J,c3111J,c3211J,c3311J,c3411J,c3511J,c3611J,c3711J,c3811J,c3911J,c3A11J,c3B11J,c3C11J,c3D11J,c3E11J,c3F11J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012J,c3112J,c3212J,c3312J,c3412J,c3512J,c3612J,c3712J,c3812J,c3912J,c3A12J,c3B12J,c3C12J,c3D12J,c3E12J,c3F12J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020J,c3120J,c3220J,c3320J,c3420J,c3520J,c3620J,c3720J,c3820J,c3920J,c3A20J,c3B20J,c3C20J,c3D20J,c3E20J,c3F20J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021J,c3121J,c3221J,c3321J,c3421J,c3521J,c3621J,c3721J,c3821J,c3921J,c3A21J,c3B21J,c3C21J,c3D21J,c3E21J,c3F21J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022J,c3122J,c3222J,c3322J,c3422J,c3522J,c3622J,c3722J,c3822J,c3922J,c3A22J,c3B22J,c3C22J,c3D22J,c3E22J,c3F22J;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000K,c3100K,c3200K,c3300K,c3400K,c3500K,c3600K,c3700K,c3800K,c3900K,c3A00K,c3B00K,c3C00K,c3D00K,c3E00K,c3F00K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001K,c3101K,c3201K,c3301K,c3401K,c3501K,c3601K,c3701K,c3801K,c3901K,c3A01K,c3B01K,c3C01K,c3D01K,c3E01K,c3F01K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002K,c3102K,c3202K,c3302K,c3402K,c3502K,c3602K,c3702K,c3802K,c3902K,c3A02K,c3B02K,c3C02K,c3D02K,c3E02K,c3F02K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010K,c3110K,c3210K,c3310K,c3410K,c3510K,c3610K,c3710K,c3810K,c3910K,c3A10K,c3B10K,c3C10K,c3D10K,c3E10K,c3F10K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011K,c3111K,c3211K,c3311K,c3411K,c3511K,c3611K,c3711K,c3811K,c3911K,c3A11K,c3B11K,c3C11K,c3D11K,c3E11K,c3F11K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012K,c3112K,c3212K,c3312K,c3412K,c3512K,c3612K,c3712K,c3812K,c3912K,c3A12K,c3B12K,c3C12K,c3D12K,c3E12K,c3F12K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020K,c3120K,c3220K,c3320K,c3420K,c3520K,c3620K,c3720K,c3820K,c3920K,c3A20K,c3B20K,c3C20K,c3D20K,c3E20K,c3F20K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021K,c3121K,c3221K,c3321K,c3421K,c3521K,c3621K,c3721K,c3821K,c3921K,c3A21K,c3B21K,c3C21K,c3D21K,c3E21K,c3F21K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022K,c3122K,c3222K,c3322K,c3422K,c3522K,c3622K,c3722K,c3822K,c3922K,c3A22K,c3B22K,c3C22K,c3D22K,c3E22K,c3F22K;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000L,c3100L,c3200L,c3300L,c3400L,c3500L,c3600L,c3700L,c3800L,c3900L,c3A00L,c3B00L,c3C00L,c3D00L,c3E00L,c3F00L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001L,c3101L,c3201L,c3301L,c3401L,c3501L,c3601L,c3701L,c3801L,c3901L,c3A01L,c3B01L,c3C01L,c3D01L,c3E01L,c3F01L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002L,c3102L,c3202L,c3302L,c3402L,c3502L,c3602L,c3702L,c3802L,c3902L,c3A02L,c3B02L,c3C02L,c3D02L,c3E02L,c3F02L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010L,c3110L,c3210L,c3310L,c3410L,c3510L,c3610L,c3710L,c3810L,c3910L,c3A10L,c3B10L,c3C10L,c3D10L,c3E10L,c3F10L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011L,c3111L,c3211L,c3311L,c3411L,c3511L,c3611L,c3711L,c3811L,c3911L,c3A11L,c3B11L,c3C11L,c3D11L,c3E11L,c3F11L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012L,c3112L,c3212L,c3312L,c3412L,c3512L,c3612L,c3712L,c3812L,c3912L,c3A12L,c3B12L,c3C12L,c3D12L,c3E12L,c3F12L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020L,c3120L,c3220L,c3320L,c3420L,c3520L,c3620L,c3720L,c3820L,c3920L,c3A20L,c3B20L,c3C20L,c3D20L,c3E20L,c3F20L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021L,c3121L,c3221L,c3321L,c3421L,c3521L,c3621L,c3721L,c3821L,c3921L,c3A21L,c3B21L,c3C21L,c3D21L,c3E21L,c3F21L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022L,c3122L,c3222L,c3322L,c3422L,c3522L,c3622L,c3722L,c3822L,c3922L,c3A22L,c3B22L,c3C22L,c3D22L,c3E22L,c3F22L;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000M,c3100M,c3200M,c3300M,c3400M,c3500M,c3600M,c3700M,c3800M,c3900M,c3A00M,c3B00M,c3C00M,c3D00M,c3E00M,c3F00M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001M,c3101M,c3201M,c3301M,c3401M,c3501M,c3601M,c3701M,c3801M,c3901M,c3A01M,c3B01M,c3C01M,c3D01M,c3E01M,c3F01M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002M,c3102M,c3202M,c3302M,c3402M,c3502M,c3602M,c3702M,c3802M,c3902M,c3A02M,c3B02M,c3C02M,c3D02M,c3E02M,c3F02M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010M,c3110M,c3210M,c3310M,c3410M,c3510M,c3610M,c3710M,c3810M,c3910M,c3A10M,c3B10M,c3C10M,c3D10M,c3E10M,c3F10M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011M,c3111M,c3211M,c3311M,c3411M,c3511M,c3611M,c3711M,c3811M,c3911M,c3A11M,c3B11M,c3C11M,c3D11M,c3E11M,c3F11M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012M,c3112M,c3212M,c3312M,c3412M,c3512M,c3612M,c3712M,c3812M,c3912M,c3A12M,c3B12M,c3C12M,c3D12M,c3E12M,c3F12M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020M,c3120M,c3220M,c3320M,c3420M,c3520M,c3620M,c3720M,c3820M,c3920M,c3A20M,c3B20M,c3C20M,c3D20M,c3E20M,c3F20M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021M,c3121M,c3221M,c3321M,c3421M,c3521M,c3621M,c3721M,c3821M,c3921M,c3A21M,c3B21M,c3C21M,c3D21M,c3E21M,c3F21M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022M,c3122M,c3222M,c3322M,c3422M,c3522M,c3622M,c3722M,c3822M,c3922M,c3A22M,c3B22M,c3C22M,c3D22M,c3E22M,c3F22M;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000N,c3100N,c3200N,c3300N,c3400N,c3500N,c3600N,c3700N,c3800N,c3900N,c3A00N,c3B00N,c3C00N,c3D00N,c3E00N,c3F00N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001N,c3101N,c3201N,c3301N,c3401N,c3501N,c3601N,c3701N,c3801N,c3901N,c3A01N,c3B01N,c3C01N,c3D01N,c3E01N,c3F01N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002N,c3102N,c3202N,c3302N,c3402N,c3502N,c3602N,c3702N,c3802N,c3902N,c3A02N,c3B02N,c3C02N,c3D02N,c3E02N,c3F02N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010N,c3110N,c3210N,c3310N,c3410N,c3510N,c3610N,c3710N,c3810N,c3910N,c3A10N,c3B10N,c3C10N,c3D10N,c3E10N,c3F10N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011N,c3111N,c3211N,c3311N,c3411N,c3511N,c3611N,c3711N,c3811N,c3911N,c3A11N,c3B11N,c3C11N,c3D11N,c3E11N,c3F11N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012N,c3112N,c3212N,c3312N,c3412N,c3512N,c3612N,c3712N,c3812N,c3912N,c3A12N,c3B12N,c3C12N,c3D12N,c3E12N,c3F12N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020N,c3120N,c3220N,c3320N,c3420N,c3520N,c3620N,c3720N,c3820N,c3920N,c3A20N,c3B20N,c3C20N,c3D20N,c3E20N,c3F20N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021N,c3121N,c3221N,c3321N,c3421N,c3521N,c3621N,c3721N,c3821N,c3921N,c3A21N,c3B21N,c3C21N,c3D21N,c3E21N,c3F21N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022N,c3122N,c3222N,c3322N,c3422N,c3522N,c3622N,c3722N,c3822N,c3922N,c3A22N,c3B22N,c3C22N,c3D22N,c3E22N,c3F22N;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000O,c3100O,c3200O,c3300O,c3400O,c3500O,c3600O,c3700O,c3800O,c3900O,c3A00O,c3B00O,c3C00O,c3D00O,c3E00O,c3F00O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001O,c3101O,c3201O,c3301O,c3401O,c3501O,c3601O,c3701O,c3801O,c3901O,c3A01O,c3B01O,c3C01O,c3D01O,c3E01O,c3F01O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002O,c3102O,c3202O,c3302O,c3402O,c3502O,c3602O,c3702O,c3802O,c3902O,c3A02O,c3B02O,c3C02O,c3D02O,c3E02O,c3F02O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010O,c3110O,c3210O,c3310O,c3410O,c3510O,c3610O,c3710O,c3810O,c3910O,c3A10O,c3B10O,c3C10O,c3D10O,c3E10O,c3F10O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011O,c3111O,c3211O,c3311O,c3411O,c3511O,c3611O,c3711O,c3811O,c3911O,c3A11O,c3B11O,c3C11O,c3D11O,c3E11O,c3F11O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012O,c3112O,c3212O,c3312O,c3412O,c3512O,c3612O,c3712O,c3812O,c3912O,c3A12O,c3B12O,c3C12O,c3D12O,c3E12O,c3F12O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020O,c3120O,c3220O,c3320O,c3420O,c3520O,c3620O,c3720O,c3820O,c3920O,c3A20O,c3B20O,c3C20O,c3D20O,c3E20O,c3F20O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021O,c3121O,c3221O,c3321O,c3421O,c3521O,c3621O,c3721O,c3821O,c3921O,c3A21O,c3B21O,c3C21O,c3D21O,c3E21O,c3F21O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022O,c3122O,c3222O,c3322O,c3422O,c3522O,c3622O,c3722O,c3822O,c3922O,c3A22O,c3B22O,c3C22O,c3D22O,c3E22O,c3F22O;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000P,c3100P,c3200P,c3300P,c3400P,c3500P,c3600P,c3700P,c3800P,c3900P,c3A00P,c3B00P,c3C00P,c3D00P,c3E00P,c3F00P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001P,c3101P,c3201P,c3301P,c3401P,c3501P,c3601P,c3701P,c3801P,c3901P,c3A01P,c3B01P,c3C01P,c3D01P,c3E01P,c3F01P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002P,c3102P,c3202P,c3302P,c3402P,c3502P,c3602P,c3702P,c3802P,c3902P,c3A02P,c3B02P,c3C02P,c3D02P,c3E02P,c3F02P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010P,c3110P,c3210P,c3310P,c3410P,c3510P,c3610P,c3710P,c3810P,c3910P,c3A10P,c3B10P,c3C10P,c3D10P,c3E10P,c3F10P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011P,c3111P,c3211P,c3311P,c3411P,c3511P,c3611P,c3711P,c3811P,c3911P,c3A11P,c3B11P,c3C11P,c3D11P,c3E11P,c3F11P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012P,c3112P,c3212P,c3312P,c3412P,c3512P,c3612P,c3712P,c3812P,c3912P,c3A12P,c3B12P,c3C12P,c3D12P,c3E12P,c3F12P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020P,c3120P,c3220P,c3320P,c3420P,c3520P,c3620P,c3720P,c3820P,c3920P,c3A20P,c3B20P,c3C20P,c3D20P,c3E20P,c3F20P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021P,c3121P,c3221P,c3321P,c3421P,c3521P,c3621P,c3721P,c3821P,c3921P,c3A21P,c3B21P,c3C21P,c3D21P,c3E21P,c3F21P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022P,c3122P,c3222P,c3322P,c3422P,c3522P,c3622P,c3722P,c3822P,c3922P,c3A22P,c3B22P,c3C22P,c3D22P,c3E22P,c3F22P;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000Q,c3100Q,c3200Q,c3300Q,c3400Q,c3500Q,c3600Q,c3700Q,c3800Q,c3900Q,c3A00Q,c3B00Q,c3C00Q,c3D00Q,c3E00Q,c3F00Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001Q,c3101Q,c3201Q,c3301Q,c3401Q,c3501Q,c3601Q,c3701Q,c3801Q,c3901Q,c3A01Q,c3B01Q,c3C01Q,c3D01Q,c3E01Q,c3F01Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002Q,c3102Q,c3202Q,c3302Q,c3402Q,c3502Q,c3602Q,c3702Q,c3802Q,c3902Q,c3A02Q,c3B02Q,c3C02Q,c3D02Q,c3E02Q,c3F02Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010Q,c3110Q,c3210Q,c3310Q,c3410Q,c3510Q,c3610Q,c3710Q,c3810Q,c3910Q,c3A10Q,c3B10Q,c3C10Q,c3D10Q,c3E10Q,c3F10Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011Q,c3111Q,c3211Q,c3311Q,c3411Q,c3511Q,c3611Q,c3711Q,c3811Q,c3911Q,c3A11Q,c3B11Q,c3C11Q,c3D11Q,c3E11Q,c3F11Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012Q,c3112Q,c3212Q,c3312Q,c3412Q,c3512Q,c3612Q,c3712Q,c3812Q,c3912Q,c3A12Q,c3B12Q,c3C12Q,c3D12Q,c3E12Q,c3F12Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020Q,c3120Q,c3220Q,c3320Q,c3420Q,c3520Q,c3620Q,c3720Q,c3820Q,c3920Q,c3A20Q,c3B20Q,c3C20Q,c3D20Q,c3E20Q,c3F20Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021Q,c3121Q,c3221Q,c3321Q,c3421Q,c3521Q,c3621Q,c3721Q,c3821Q,c3921Q,c3A21Q,c3B21Q,c3C21Q,c3D21Q,c3E21Q,c3F21Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022Q,c3122Q,c3222Q,c3322Q,c3422Q,c3522Q,c3622Q,c3722Q,c3822Q,c3922Q,c3A22Q,c3B22Q,c3C22Q,c3D22Q,c3E22Q,c3F22Q;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000R,c3100R,c3200R,c3300R,c3400R,c3500R,c3600R,c3700R,c3800R,c3900R,c3A00R,c3B00R,c3C00R,c3D00R,c3E00R,c3F00R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001R,c3101R,c3201R,c3301R,c3401R,c3501R,c3601R,c3701R,c3801R,c3901R,c3A01R,c3B01R,c3C01R,c3D01R,c3E01R,c3F01R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002R,c3102R,c3202R,c3302R,c3402R,c3502R,c3602R,c3702R,c3802R,c3902R,c3A02R,c3B02R,c3C02R,c3D02R,c3E02R,c3F02R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010R,c3110R,c3210R,c3310R,c3410R,c3510R,c3610R,c3710R,c3810R,c3910R,c3A10R,c3B10R,c3C10R,c3D10R,c3E10R,c3F10R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011R,c3111R,c3211R,c3311R,c3411R,c3511R,c3611R,c3711R,c3811R,c3911R,c3A11R,c3B11R,c3C11R,c3D11R,c3E11R,c3F11R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012R,c3112R,c3212R,c3312R,c3412R,c3512R,c3612R,c3712R,c3812R,c3912R,c3A12R,c3B12R,c3C12R,c3D12R,c3E12R,c3F12R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020R,c3120R,c3220R,c3320R,c3420R,c3520R,c3620R,c3720R,c3820R,c3920R,c3A20R,c3B20R,c3C20R,c3D20R,c3E20R,c3F20R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021R,c3121R,c3221R,c3321R,c3421R,c3521R,c3621R,c3721R,c3821R,c3921R,c3A21R,c3B21R,c3C21R,c3D21R,c3E21R,c3F21R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022R,c3122R,c3222R,c3322R,c3422R,c3522R,c3622R,c3722R,c3822R,c3922R,c3A22R,c3B22R,c3C22R,c3D22R,c3E22R,c3F22R;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000S,c3100S,c3200S,c3300S,c3400S,c3500S,c3600S,c3700S,c3800S,c3900S,c3A00S,c3B00S,c3C00S,c3D00S,c3E00S,c3F00S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001S,c3101S,c3201S,c3301S,c3401S,c3501S,c3601S,c3701S,c3801S,c3901S,c3A01S,c3B01S,c3C01S,c3D01S,c3E01S,c3F01S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002S,c3102S,c3202S,c3302S,c3402S,c3502S,c3602S,c3702S,c3802S,c3902S,c3A02S,c3B02S,c3C02S,c3D02S,c3E02S,c3F02S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010S,c3110S,c3210S,c3310S,c3410S,c3510S,c3610S,c3710S,c3810S,c3910S,c3A10S,c3B10S,c3C10S,c3D10S,c3E10S,c3F10S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011S,c3111S,c3211S,c3311S,c3411S,c3511S,c3611S,c3711S,c3811S,c3911S,c3A11S,c3B11S,c3C11S,c3D11S,c3E11S,c3F11S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012S,c3112S,c3212S,c3312S,c3412S,c3512S,c3612S,c3712S,c3812S,c3912S,c3A12S,c3B12S,c3C12S,c3D12S,c3E12S,c3F12S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020S,c3120S,c3220S,c3320S,c3420S,c3520S,c3620S,c3720S,c3820S,c3920S,c3A20S,c3B20S,c3C20S,c3D20S,c3E20S,c3F20S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021S,c3121S,c3221S,c3321S,c3421S,c3521S,c3621S,c3721S,c3821S,c3921S,c3A21S,c3B21S,c3C21S,c3D21S,c3E21S,c3F21S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022S,c3122S,c3222S,c3322S,c3422S,c3522S,c3622S,c3722S,c3822S,c3922S,c3A22S,c3B22S,c3C22S,c3D22S,c3E22S,c3F22S;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000T,c3100T,c3200T,c3300T,c3400T,c3500T,c3600T,c3700T,c3800T,c3900T,c3A00T,c3B00T,c3C00T,c3D00T,c3E00T,c3F00T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001T,c3101T,c3201T,c3301T,c3401T,c3501T,c3601T,c3701T,c3801T,c3901T,c3A01T,c3B01T,c3C01T,c3D01T,c3E01T,c3F01T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002T,c3102T,c3202T,c3302T,c3402T,c3502T,c3602T,c3702T,c3802T,c3902T,c3A02T,c3B02T,c3C02T,c3D02T,c3E02T,c3F02T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010T,c3110T,c3210T,c3310T,c3410T,c3510T,c3610T,c3710T,c3810T,c3910T,c3A10T,c3B10T,c3C10T,c3D10T,c3E10T,c3F10T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011T,c3111T,c3211T,c3311T,c3411T,c3511T,c3611T,c3711T,c3811T,c3911T,c3A11T,c3B11T,c3C11T,c3D11T,c3E11T,c3F11T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012T,c3112T,c3212T,c3312T,c3412T,c3512T,c3612T,c3712T,c3812T,c3912T,c3A12T,c3B12T,c3C12T,c3D12T,c3E12T,c3F12T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020T,c3120T,c3220T,c3320T,c3420T,c3520T,c3620T,c3720T,c3820T,c3920T,c3A20T,c3B20T,c3C20T,c3D20T,c3E20T,c3F20T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021T,c3121T,c3221T,c3321T,c3421T,c3521T,c3621T,c3721T,c3821T,c3921T,c3A21T,c3B21T,c3C21T,c3D21T,c3E21T,c3F21T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022T,c3122T,c3222T,c3322T,c3422T,c3522T,c3622T,c3722T,c3822T,c3922T,c3A22T,c3B22T,c3C22T,c3D22T,c3E22T,c3F22T;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000U,c3100U,c3200U,c3300U,c3400U,c3500U,c3600U,c3700U,c3800U,c3900U,c3A00U,c3B00U,c3C00U,c3D00U,c3E00U,c3F00U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001U,c3101U,c3201U,c3301U,c3401U,c3501U,c3601U,c3701U,c3801U,c3901U,c3A01U,c3B01U,c3C01U,c3D01U,c3E01U,c3F01U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002U,c3102U,c3202U,c3302U,c3402U,c3502U,c3602U,c3702U,c3802U,c3902U,c3A02U,c3B02U,c3C02U,c3D02U,c3E02U,c3F02U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010U,c3110U,c3210U,c3310U,c3410U,c3510U,c3610U,c3710U,c3810U,c3910U,c3A10U,c3B10U,c3C10U,c3D10U,c3E10U,c3F10U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011U,c3111U,c3211U,c3311U,c3411U,c3511U,c3611U,c3711U,c3811U,c3911U,c3A11U,c3B11U,c3C11U,c3D11U,c3E11U,c3F11U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012U,c3112U,c3212U,c3312U,c3412U,c3512U,c3612U,c3712U,c3812U,c3912U,c3A12U,c3B12U,c3C12U,c3D12U,c3E12U,c3F12U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020U,c3120U,c3220U,c3320U,c3420U,c3520U,c3620U,c3720U,c3820U,c3920U,c3A20U,c3B20U,c3C20U,c3D20U,c3E20U,c3F20U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021U,c3121U,c3221U,c3321U,c3421U,c3521U,c3621U,c3721U,c3821U,c3921U,c3A21U,c3B21U,c3C21U,c3D21U,c3E21U,c3F21U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022U,c3122U,c3222U,c3322U,c3422U,c3522U,c3622U,c3722U,c3822U,c3922U,c3A22U,c3B22U,c3C22U,c3D22U,c3E22U,c3F22U;
(*DONT_TOUCH="true"*) wire signed [4:0] c3000V,c3100V,c3200V,c3300V,c3400V,c3500V,c3600V,c3700V,c3800V,c3900V,c3A00V,c3B00V,c3C00V,c3D00V,c3E00V,c3F00V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3001V,c3101V,c3201V,c3301V,c3401V,c3501V,c3601V,c3701V,c3801V,c3901V,c3A01V,c3B01V,c3C01V,c3D01V,c3E01V,c3F01V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3002V,c3102V,c3202V,c3302V,c3402V,c3502V,c3602V,c3702V,c3802V,c3902V,c3A02V,c3B02V,c3C02V,c3D02V,c3E02V,c3F02V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3010V,c3110V,c3210V,c3310V,c3410V,c3510V,c3610V,c3710V,c3810V,c3910V,c3A10V,c3B10V,c3C10V,c3D10V,c3E10V,c3F10V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3011V,c3111V,c3211V,c3311V,c3411V,c3511V,c3611V,c3711V,c3811V,c3911V,c3A11V,c3B11V,c3C11V,c3D11V,c3E11V,c3F11V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3012V,c3112V,c3212V,c3312V,c3412V,c3512V,c3612V,c3712V,c3812V,c3912V,c3A12V,c3B12V,c3C12V,c3D12V,c3E12V,c3F12V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3020V,c3120V,c3220V,c3320V,c3420V,c3520V,c3620V,c3720V,c3820V,c3920V,c3A20V,c3B20V,c3C20V,c3D20V,c3E20V,c3F20V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3021V,c3121V,c3221V,c3321V,c3421V,c3521V,c3621V,c3721V,c3821V,c3921V,c3A21V,c3B21V,c3C21V,c3D21V,c3E21V,c3F21V;
(*DONT_TOUCH="true"*) wire signed [4:0] c3022V,c3122V,c3222V,c3322V,c3422V,c3522V,c3622V,c3722V,c3822V,c3922V,c3A22V,c3B22V,c3C22V,c3D22V,c3E22V,c3F22V;
(*DONT_TOUCH="true"*) wire signed [8:0] C3000;
(*DONT_TOUCH="true"*) wire A3000;
(*DONT_TOUCH="true"*) wire signed [8:0] C3010;
(*DONT_TOUCH="true"*) wire A3010;
(*DONT_TOUCH="true"*) wire signed [8:0] C3020;
(*DONT_TOUCH="true"*) wire A3020;
(*DONT_TOUCH="true"*) wire signed [8:0] C3100;
(*DONT_TOUCH="true"*) wire A3100;
(*DONT_TOUCH="true"*) wire signed [8:0] C3110;
(*DONT_TOUCH="true"*) wire A3110;
(*DONT_TOUCH="true"*) wire signed [8:0] C3120;
(*DONT_TOUCH="true"*) wire A3120;
(*DONT_TOUCH="true"*) wire signed [8:0] C3200;
(*DONT_TOUCH="true"*) wire A3200;
(*DONT_TOUCH="true"*) wire signed [8:0] C3210;
(*DONT_TOUCH="true"*) wire A3210;
(*DONT_TOUCH="true"*) wire signed [8:0] C3220;
(*DONT_TOUCH="true"*) wire A3220;
(*DONT_TOUCH="true"*) wire signed [8:0] C3001;
(*DONT_TOUCH="true"*) wire A3001;
(*DONT_TOUCH="true"*) wire signed [8:0] C3011;
(*DONT_TOUCH="true"*) wire A3011;
(*DONT_TOUCH="true"*) wire signed [8:0] C3021;
(*DONT_TOUCH="true"*) wire A3021;
(*DONT_TOUCH="true"*) wire signed [8:0] C3101;
(*DONT_TOUCH="true"*) wire A3101;
(*DONT_TOUCH="true"*) wire signed [8:0] C3111;
(*DONT_TOUCH="true"*) wire A3111;
(*DONT_TOUCH="true"*) wire signed [8:0] C3121;
(*DONT_TOUCH="true"*) wire A3121;
(*DONT_TOUCH="true"*) wire signed [8:0] C3201;
(*DONT_TOUCH="true"*) wire A3201;
(*DONT_TOUCH="true"*) wire signed [8:0] C3211;
(*DONT_TOUCH="true"*) wire A3211;
(*DONT_TOUCH="true"*) wire signed [8:0] C3221;
(*DONT_TOUCH="true"*) wire A3221;
(*DONT_TOUCH="true"*) wire signed [8:0] C3002;
(*DONT_TOUCH="true"*) wire A3002;
(*DONT_TOUCH="true"*) wire signed [8:0] C3012;
(*DONT_TOUCH="true"*) wire A3012;
(*DONT_TOUCH="true"*) wire signed [8:0] C3022;
(*DONT_TOUCH="true"*) wire A3022;
(*DONT_TOUCH="true"*) wire signed [8:0] C3102;
(*DONT_TOUCH="true"*) wire A3102;
(*DONT_TOUCH="true"*) wire signed [8:0] C3112;
(*DONT_TOUCH="true"*) wire A3112;
(*DONT_TOUCH="true"*) wire signed [8:0] C3122;
(*DONT_TOUCH="true"*) wire A3122;
(*DONT_TOUCH="true"*) wire signed [8:0] C3202;
(*DONT_TOUCH="true"*) wire A3202;
(*DONT_TOUCH="true"*) wire signed [8:0] C3212;
(*DONT_TOUCH="true"*) wire A3212;
(*DONT_TOUCH="true"*) wire signed [8:0] C3222;
(*DONT_TOUCH="true"*) wire A3222;
(*DONT_TOUCH="true"*) wire signed [8:0] C3003;
(*DONT_TOUCH="true"*) wire A3003;
(*DONT_TOUCH="true"*) wire signed [8:0] C3013;
(*DONT_TOUCH="true"*) wire A3013;
(*DONT_TOUCH="true"*) wire signed [8:0] C3023;
(*DONT_TOUCH="true"*) wire A3023;
(*DONT_TOUCH="true"*) wire signed [8:0] C3103;
(*DONT_TOUCH="true"*) wire A3103;
(*DONT_TOUCH="true"*) wire signed [8:0] C3113;
(*DONT_TOUCH="true"*) wire A3113;
(*DONT_TOUCH="true"*) wire signed [8:0] C3123;
(*DONT_TOUCH="true"*) wire A3123;
(*DONT_TOUCH="true"*) wire signed [8:0] C3203;
(*DONT_TOUCH="true"*) wire A3203;
(*DONT_TOUCH="true"*) wire signed [8:0] C3213;
(*DONT_TOUCH="true"*) wire A3213;
(*DONT_TOUCH="true"*) wire signed [8:0] C3223;
(*DONT_TOUCH="true"*) wire A3223;
(*DONT_TOUCH="true"*) wire signed [8:0] C3004;
(*DONT_TOUCH="true"*) wire A3004;
(*DONT_TOUCH="true"*) wire signed [8:0] C3014;
(*DONT_TOUCH="true"*) wire A3014;
(*DONT_TOUCH="true"*) wire signed [8:0] C3024;
(*DONT_TOUCH="true"*) wire A3024;
(*DONT_TOUCH="true"*) wire signed [8:0] C3104;
(*DONT_TOUCH="true"*) wire A3104;
(*DONT_TOUCH="true"*) wire signed [8:0] C3114;
(*DONT_TOUCH="true"*) wire A3114;
(*DONT_TOUCH="true"*) wire signed [8:0] C3124;
(*DONT_TOUCH="true"*) wire A3124;
(*DONT_TOUCH="true"*) wire signed [8:0] C3204;
(*DONT_TOUCH="true"*) wire A3204;
(*DONT_TOUCH="true"*) wire signed [8:0] C3214;
(*DONT_TOUCH="true"*) wire A3214;
(*DONT_TOUCH="true"*) wire signed [8:0] C3224;
(*DONT_TOUCH="true"*) wire A3224;
(*DONT_TOUCH="true"*) wire signed [8:0] C3005;
(*DONT_TOUCH="true"*) wire A3005;
(*DONT_TOUCH="true"*) wire signed [8:0] C3015;
(*DONT_TOUCH="true"*) wire A3015;
(*DONT_TOUCH="true"*) wire signed [8:0] C3025;
(*DONT_TOUCH="true"*) wire A3025;
(*DONT_TOUCH="true"*) wire signed [8:0] C3105;
(*DONT_TOUCH="true"*) wire A3105;
(*DONT_TOUCH="true"*) wire signed [8:0] C3115;
(*DONT_TOUCH="true"*) wire A3115;
(*DONT_TOUCH="true"*) wire signed [8:0] C3125;
(*DONT_TOUCH="true"*) wire A3125;
(*DONT_TOUCH="true"*) wire signed [8:0] C3205;
(*DONT_TOUCH="true"*) wire A3205;
(*DONT_TOUCH="true"*) wire signed [8:0] C3215;
(*DONT_TOUCH="true"*) wire A3215;
(*DONT_TOUCH="true"*) wire signed [8:0] C3225;
(*DONT_TOUCH="true"*) wire A3225;
(*DONT_TOUCH="true"*) wire signed [8:0] C3006;
(*DONT_TOUCH="true"*) wire A3006;
(*DONT_TOUCH="true"*) wire signed [8:0] C3016;
(*DONT_TOUCH="true"*) wire A3016;
(*DONT_TOUCH="true"*) wire signed [8:0] C3026;
(*DONT_TOUCH="true"*) wire A3026;
(*DONT_TOUCH="true"*) wire signed [8:0] C3106;
(*DONT_TOUCH="true"*) wire A3106;
(*DONT_TOUCH="true"*) wire signed [8:0] C3116;
(*DONT_TOUCH="true"*) wire A3116;
(*DONT_TOUCH="true"*) wire signed [8:0] C3126;
(*DONT_TOUCH="true"*) wire A3126;
(*DONT_TOUCH="true"*) wire signed [8:0] C3206;
(*DONT_TOUCH="true"*) wire A3206;
(*DONT_TOUCH="true"*) wire signed [8:0] C3216;
(*DONT_TOUCH="true"*) wire A3216;
(*DONT_TOUCH="true"*) wire signed [8:0] C3226;
(*DONT_TOUCH="true"*) wire A3226;
(*DONT_TOUCH="true"*) wire signed [8:0] C3007;
(*DONT_TOUCH="true"*) wire A3007;
(*DONT_TOUCH="true"*) wire signed [8:0] C3017;
(*DONT_TOUCH="true"*) wire A3017;
(*DONT_TOUCH="true"*) wire signed [8:0] C3027;
(*DONT_TOUCH="true"*) wire A3027;
(*DONT_TOUCH="true"*) wire signed [8:0] C3107;
(*DONT_TOUCH="true"*) wire A3107;
(*DONT_TOUCH="true"*) wire signed [8:0] C3117;
(*DONT_TOUCH="true"*) wire A3117;
(*DONT_TOUCH="true"*) wire signed [8:0] C3127;
(*DONT_TOUCH="true"*) wire A3127;
(*DONT_TOUCH="true"*) wire signed [8:0] C3207;
(*DONT_TOUCH="true"*) wire A3207;
(*DONT_TOUCH="true"*) wire signed [8:0] C3217;
(*DONT_TOUCH="true"*) wire A3217;
(*DONT_TOUCH="true"*) wire signed [8:0] C3227;
(*DONT_TOUCH="true"*) wire A3227;
(*DONT_TOUCH="true"*) wire signed [8:0] C3008;
(*DONT_TOUCH="true"*) wire A3008;
(*DONT_TOUCH="true"*) wire signed [8:0] C3018;
(*DONT_TOUCH="true"*) wire A3018;
(*DONT_TOUCH="true"*) wire signed [8:0] C3028;
(*DONT_TOUCH="true"*) wire A3028;
(*DONT_TOUCH="true"*) wire signed [8:0] C3108;
(*DONT_TOUCH="true"*) wire A3108;
(*DONT_TOUCH="true"*) wire signed [8:0] C3118;
(*DONT_TOUCH="true"*) wire A3118;
(*DONT_TOUCH="true"*) wire signed [8:0] C3128;
(*DONT_TOUCH="true"*) wire A3128;
(*DONT_TOUCH="true"*) wire signed [8:0] C3208;
(*DONT_TOUCH="true"*) wire A3208;
(*DONT_TOUCH="true"*) wire signed [8:0] C3218;
(*DONT_TOUCH="true"*) wire A3218;
(*DONT_TOUCH="true"*) wire signed [8:0] C3228;
(*DONT_TOUCH="true"*) wire A3228;
(*DONT_TOUCH="true"*) wire signed [8:0] C3009;
(*DONT_TOUCH="true"*) wire A3009;
(*DONT_TOUCH="true"*) wire signed [8:0] C3019;
(*DONT_TOUCH="true"*) wire A3019;
(*DONT_TOUCH="true"*) wire signed [8:0] C3029;
(*DONT_TOUCH="true"*) wire A3029;
(*DONT_TOUCH="true"*) wire signed [8:0] C3109;
(*DONT_TOUCH="true"*) wire A3109;
(*DONT_TOUCH="true"*) wire signed [8:0] C3119;
(*DONT_TOUCH="true"*) wire A3119;
(*DONT_TOUCH="true"*) wire signed [8:0] C3129;
(*DONT_TOUCH="true"*) wire A3129;
(*DONT_TOUCH="true"*) wire signed [8:0] C3209;
(*DONT_TOUCH="true"*) wire A3209;
(*DONT_TOUCH="true"*) wire signed [8:0] C3219;
(*DONT_TOUCH="true"*) wire A3219;
(*DONT_TOUCH="true"*) wire signed [8:0] C3229;
(*DONT_TOUCH="true"*) wire A3229;
(*DONT_TOUCH="true"*) wire signed [8:0] C300A;
(*DONT_TOUCH="true"*) wire A300A;
(*DONT_TOUCH="true"*) wire signed [8:0] C301A;
(*DONT_TOUCH="true"*) wire A301A;
(*DONT_TOUCH="true"*) wire signed [8:0] C302A;
(*DONT_TOUCH="true"*) wire A302A;
(*DONT_TOUCH="true"*) wire signed [8:0] C310A;
(*DONT_TOUCH="true"*) wire A310A;
(*DONT_TOUCH="true"*) wire signed [8:0] C311A;
(*DONT_TOUCH="true"*) wire A311A;
(*DONT_TOUCH="true"*) wire signed [8:0] C312A;
(*DONT_TOUCH="true"*) wire A312A;
(*DONT_TOUCH="true"*) wire signed [8:0] C320A;
(*DONT_TOUCH="true"*) wire A320A;
(*DONT_TOUCH="true"*) wire signed [8:0] C321A;
(*DONT_TOUCH="true"*) wire A321A;
(*DONT_TOUCH="true"*) wire signed [8:0] C322A;
(*DONT_TOUCH="true"*) wire A322A;
(*DONT_TOUCH="true"*) wire signed [8:0] C300B;
(*DONT_TOUCH="true"*) wire A300B;
(*DONT_TOUCH="true"*) wire signed [8:0] C301B;
(*DONT_TOUCH="true"*) wire A301B;
(*DONT_TOUCH="true"*) wire signed [8:0] C302B;
(*DONT_TOUCH="true"*) wire A302B;
(*DONT_TOUCH="true"*) wire signed [8:0] C310B;
(*DONT_TOUCH="true"*) wire A310B;
(*DONT_TOUCH="true"*) wire signed [8:0] C311B;
(*DONT_TOUCH="true"*) wire A311B;
(*DONT_TOUCH="true"*) wire signed [8:0] C312B;
(*DONT_TOUCH="true"*) wire A312B;
(*DONT_TOUCH="true"*) wire signed [8:0] C320B;
(*DONT_TOUCH="true"*) wire A320B;
(*DONT_TOUCH="true"*) wire signed [8:0] C321B;
(*DONT_TOUCH="true"*) wire A321B;
(*DONT_TOUCH="true"*) wire signed [8:0] C322B;
(*DONT_TOUCH="true"*) wire A322B;
(*DONT_TOUCH="true"*) wire signed [8:0] C300C;
(*DONT_TOUCH="true"*) wire A300C;
(*DONT_TOUCH="true"*) wire signed [8:0] C301C;
(*DONT_TOUCH="true"*) wire A301C;
(*DONT_TOUCH="true"*) wire signed [8:0] C302C;
(*DONT_TOUCH="true"*) wire A302C;
(*DONT_TOUCH="true"*) wire signed [8:0] C310C;
(*DONT_TOUCH="true"*) wire A310C;
(*DONT_TOUCH="true"*) wire signed [8:0] C311C;
(*DONT_TOUCH="true"*) wire A311C;
(*DONT_TOUCH="true"*) wire signed [8:0] C312C;
(*DONT_TOUCH="true"*) wire A312C;
(*DONT_TOUCH="true"*) wire signed [8:0] C320C;
(*DONT_TOUCH="true"*) wire A320C;
(*DONT_TOUCH="true"*) wire signed [8:0] C321C;
(*DONT_TOUCH="true"*) wire A321C;
(*DONT_TOUCH="true"*) wire signed [8:0] C322C;
(*DONT_TOUCH="true"*) wire A322C;
(*DONT_TOUCH="true"*) wire signed [8:0] C300D;
(*DONT_TOUCH="true"*) wire A300D;
(*DONT_TOUCH="true"*) wire signed [8:0] C301D;
(*DONT_TOUCH="true"*) wire A301D;
(*DONT_TOUCH="true"*) wire signed [8:0] C302D;
(*DONT_TOUCH="true"*) wire A302D;
(*DONT_TOUCH="true"*) wire signed [8:0] C310D;
(*DONT_TOUCH="true"*) wire A310D;
(*DONT_TOUCH="true"*) wire signed [8:0] C311D;
(*DONT_TOUCH="true"*) wire A311D;
(*DONT_TOUCH="true"*) wire signed [8:0] C312D;
(*DONT_TOUCH="true"*) wire A312D;
(*DONT_TOUCH="true"*) wire signed [8:0] C320D;
(*DONT_TOUCH="true"*) wire A320D;
(*DONT_TOUCH="true"*) wire signed [8:0] C321D;
(*DONT_TOUCH="true"*) wire A321D;
(*DONT_TOUCH="true"*) wire signed [8:0] C322D;
(*DONT_TOUCH="true"*) wire A322D;
(*DONT_TOUCH="true"*) wire signed [8:0] C300E;
(*DONT_TOUCH="true"*) wire A300E;
(*DONT_TOUCH="true"*) wire signed [8:0] C301E;
(*DONT_TOUCH="true"*) wire A301E;
(*DONT_TOUCH="true"*) wire signed [8:0] C302E;
(*DONT_TOUCH="true"*) wire A302E;
(*DONT_TOUCH="true"*) wire signed [8:0] C310E;
(*DONT_TOUCH="true"*) wire A310E;
(*DONT_TOUCH="true"*) wire signed [8:0] C311E;
(*DONT_TOUCH="true"*) wire A311E;
(*DONT_TOUCH="true"*) wire signed [8:0] C312E;
(*DONT_TOUCH="true"*) wire A312E;
(*DONT_TOUCH="true"*) wire signed [8:0] C320E;
(*DONT_TOUCH="true"*) wire A320E;
(*DONT_TOUCH="true"*) wire signed [8:0] C321E;
(*DONT_TOUCH="true"*) wire A321E;
(*DONT_TOUCH="true"*) wire signed [8:0] C322E;
(*DONT_TOUCH="true"*) wire A322E;
(*DONT_TOUCH="true"*) wire signed [8:0] C300F;
(*DONT_TOUCH="true"*) wire A300F;
(*DONT_TOUCH="true"*) wire signed [8:0] C301F;
(*DONT_TOUCH="true"*) wire A301F;
(*DONT_TOUCH="true"*) wire signed [8:0] C302F;
(*DONT_TOUCH="true"*) wire A302F;
(*DONT_TOUCH="true"*) wire signed [8:0] C310F;
(*DONT_TOUCH="true"*) wire A310F;
(*DONT_TOUCH="true"*) wire signed [8:0] C311F;
(*DONT_TOUCH="true"*) wire A311F;
(*DONT_TOUCH="true"*) wire signed [8:0] C312F;
(*DONT_TOUCH="true"*) wire A312F;
(*DONT_TOUCH="true"*) wire signed [8:0] C320F;
(*DONT_TOUCH="true"*) wire A320F;
(*DONT_TOUCH="true"*) wire signed [8:0] C321F;
(*DONT_TOUCH="true"*) wire A321F;
(*DONT_TOUCH="true"*) wire signed [8:0] C322F;
(*DONT_TOUCH="true"*) wire A322F;
(*DONT_TOUCH="true"*) wire signed [8:0] C300G;
(*DONT_TOUCH="true"*) wire A300G;
(*DONT_TOUCH="true"*) wire signed [8:0] C301G;
(*DONT_TOUCH="true"*) wire A301G;
(*DONT_TOUCH="true"*) wire signed [8:0] C302G;
(*DONT_TOUCH="true"*) wire A302G;
(*DONT_TOUCH="true"*) wire signed [8:0] C310G;
(*DONT_TOUCH="true"*) wire A310G;
(*DONT_TOUCH="true"*) wire signed [8:0] C311G;
(*DONT_TOUCH="true"*) wire A311G;
(*DONT_TOUCH="true"*) wire signed [8:0] C312G;
(*DONT_TOUCH="true"*) wire A312G;
(*DONT_TOUCH="true"*) wire signed [8:0] C320G;
(*DONT_TOUCH="true"*) wire A320G;
(*DONT_TOUCH="true"*) wire signed [8:0] C321G;
(*DONT_TOUCH="true"*) wire A321G;
(*DONT_TOUCH="true"*) wire signed [8:0] C322G;
(*DONT_TOUCH="true"*) wire A322G;
(*DONT_TOUCH="true"*) wire signed [8:0] C300H;
(*DONT_TOUCH="true"*) wire A300H;
(*DONT_TOUCH="true"*) wire signed [8:0] C301H;
(*DONT_TOUCH="true"*) wire A301H;
(*DONT_TOUCH="true"*) wire signed [8:0] C302H;
(*DONT_TOUCH="true"*) wire A302H;
(*DONT_TOUCH="true"*) wire signed [8:0] C310H;
(*DONT_TOUCH="true"*) wire A310H;
(*DONT_TOUCH="true"*) wire signed [8:0] C311H;
(*DONT_TOUCH="true"*) wire A311H;
(*DONT_TOUCH="true"*) wire signed [8:0] C312H;
(*DONT_TOUCH="true"*) wire A312H;
(*DONT_TOUCH="true"*) wire signed [8:0] C320H;
(*DONT_TOUCH="true"*) wire A320H;
(*DONT_TOUCH="true"*) wire signed [8:0] C321H;
(*DONT_TOUCH="true"*) wire A321H;
(*DONT_TOUCH="true"*) wire signed [8:0] C322H;
(*DONT_TOUCH="true"*) wire A322H;
(*DONT_TOUCH="true"*) wire signed [8:0] C300I;
(*DONT_TOUCH="true"*) wire A300I;
(*DONT_TOUCH="true"*) wire signed [8:0] C301I;
(*DONT_TOUCH="true"*) wire A301I;
(*DONT_TOUCH="true"*) wire signed [8:0] C302I;
(*DONT_TOUCH="true"*) wire A302I;
(*DONT_TOUCH="true"*) wire signed [8:0] C310I;
(*DONT_TOUCH="true"*) wire A310I;
(*DONT_TOUCH="true"*) wire signed [8:0] C311I;
(*DONT_TOUCH="true"*) wire A311I;
(*DONT_TOUCH="true"*) wire signed [8:0] C312I;
(*DONT_TOUCH="true"*) wire A312I;
(*DONT_TOUCH="true"*) wire signed [8:0] C320I;
(*DONT_TOUCH="true"*) wire A320I;
(*DONT_TOUCH="true"*) wire signed [8:0] C321I;
(*DONT_TOUCH="true"*) wire A321I;
(*DONT_TOUCH="true"*) wire signed [8:0] C322I;
(*DONT_TOUCH="true"*) wire A322I;
(*DONT_TOUCH="true"*) wire signed [8:0] C300J;
(*DONT_TOUCH="true"*) wire A300J;
(*DONT_TOUCH="true"*) wire signed [8:0] C301J;
(*DONT_TOUCH="true"*) wire A301J;
(*DONT_TOUCH="true"*) wire signed [8:0] C302J;
(*DONT_TOUCH="true"*) wire A302J;
(*DONT_TOUCH="true"*) wire signed [8:0] C310J;
(*DONT_TOUCH="true"*) wire A310J;
(*DONT_TOUCH="true"*) wire signed [8:0] C311J;
(*DONT_TOUCH="true"*) wire A311J;
(*DONT_TOUCH="true"*) wire signed [8:0] C312J;
(*DONT_TOUCH="true"*) wire A312J;
(*DONT_TOUCH="true"*) wire signed [8:0] C320J;
(*DONT_TOUCH="true"*) wire A320J;
(*DONT_TOUCH="true"*) wire signed [8:0] C321J;
(*DONT_TOUCH="true"*) wire A321J;
(*DONT_TOUCH="true"*) wire signed [8:0] C322J;
(*DONT_TOUCH="true"*) wire A322J;
(*DONT_TOUCH="true"*) wire signed [8:0] C300K;
(*DONT_TOUCH="true"*) wire A300K;
(*DONT_TOUCH="true"*) wire signed [8:0] C301K;
(*DONT_TOUCH="true"*) wire A301K;
(*DONT_TOUCH="true"*) wire signed [8:0] C302K;
(*DONT_TOUCH="true"*) wire A302K;
(*DONT_TOUCH="true"*) wire signed [8:0] C310K;
(*DONT_TOUCH="true"*) wire A310K;
(*DONT_TOUCH="true"*) wire signed [8:0] C311K;
(*DONT_TOUCH="true"*) wire A311K;
(*DONT_TOUCH="true"*) wire signed [8:0] C312K;
(*DONT_TOUCH="true"*) wire A312K;
(*DONT_TOUCH="true"*) wire signed [8:0] C320K;
(*DONT_TOUCH="true"*) wire A320K;
(*DONT_TOUCH="true"*) wire signed [8:0] C321K;
(*DONT_TOUCH="true"*) wire A321K;
(*DONT_TOUCH="true"*) wire signed [8:0] C322K;
(*DONT_TOUCH="true"*) wire A322K;
(*DONT_TOUCH="true"*) wire signed [8:0] C300L;
(*DONT_TOUCH="true"*) wire A300L;
(*DONT_TOUCH="true"*) wire signed [8:0] C301L;
(*DONT_TOUCH="true"*) wire A301L;
(*DONT_TOUCH="true"*) wire signed [8:0] C302L;
(*DONT_TOUCH="true"*) wire A302L;
(*DONT_TOUCH="true"*) wire signed [8:0] C310L;
(*DONT_TOUCH="true"*) wire A310L;
(*DONT_TOUCH="true"*) wire signed [8:0] C311L;
(*DONT_TOUCH="true"*) wire A311L;
(*DONT_TOUCH="true"*) wire signed [8:0] C312L;
(*DONT_TOUCH="true"*) wire A312L;
(*DONT_TOUCH="true"*) wire signed [8:0] C320L;
(*DONT_TOUCH="true"*) wire A320L;
(*DONT_TOUCH="true"*) wire signed [8:0] C321L;
(*DONT_TOUCH="true"*) wire A321L;
(*DONT_TOUCH="true"*) wire signed [8:0] C322L;
(*DONT_TOUCH="true"*) wire A322L;
(*DONT_TOUCH="true"*) wire signed [8:0] C300M;
(*DONT_TOUCH="true"*) wire A300M;
(*DONT_TOUCH="true"*) wire signed [8:0] C301M;
(*DONT_TOUCH="true"*) wire A301M;
(*DONT_TOUCH="true"*) wire signed [8:0] C302M;
(*DONT_TOUCH="true"*) wire A302M;
(*DONT_TOUCH="true"*) wire signed [8:0] C310M;
(*DONT_TOUCH="true"*) wire A310M;
(*DONT_TOUCH="true"*) wire signed [8:0] C311M;
(*DONT_TOUCH="true"*) wire A311M;
(*DONT_TOUCH="true"*) wire signed [8:0] C312M;
(*DONT_TOUCH="true"*) wire A312M;
(*DONT_TOUCH="true"*) wire signed [8:0] C320M;
(*DONT_TOUCH="true"*) wire A320M;
(*DONT_TOUCH="true"*) wire signed [8:0] C321M;
(*DONT_TOUCH="true"*) wire A321M;
(*DONT_TOUCH="true"*) wire signed [8:0] C322M;
(*DONT_TOUCH="true"*) wire A322M;
(*DONT_TOUCH="true"*) wire signed [8:0] C300N;
(*DONT_TOUCH="true"*) wire A300N;
(*DONT_TOUCH="true"*) wire signed [8:0] C301N;
(*DONT_TOUCH="true"*) wire A301N;
(*DONT_TOUCH="true"*) wire signed [8:0] C302N;
(*DONT_TOUCH="true"*) wire A302N;
(*DONT_TOUCH="true"*) wire signed [8:0] C310N;
(*DONT_TOUCH="true"*) wire A310N;
(*DONT_TOUCH="true"*) wire signed [8:0] C311N;
(*DONT_TOUCH="true"*) wire A311N;
(*DONT_TOUCH="true"*) wire signed [8:0] C312N;
(*DONT_TOUCH="true"*) wire A312N;
(*DONT_TOUCH="true"*) wire signed [8:0] C320N;
(*DONT_TOUCH="true"*) wire A320N;
(*DONT_TOUCH="true"*) wire signed [8:0] C321N;
(*DONT_TOUCH="true"*) wire A321N;
(*DONT_TOUCH="true"*) wire signed [8:0] C322N;
(*DONT_TOUCH="true"*) wire A322N;
(*DONT_TOUCH="true"*) wire signed [8:0] C300O;
(*DONT_TOUCH="true"*) wire A300O;
(*DONT_TOUCH="true"*) wire signed [8:0] C301O;
(*DONT_TOUCH="true"*) wire A301O;
(*DONT_TOUCH="true"*) wire signed [8:0] C302O;
(*DONT_TOUCH="true"*) wire A302O;
(*DONT_TOUCH="true"*) wire signed [8:0] C310O;
(*DONT_TOUCH="true"*) wire A310O;
(*DONT_TOUCH="true"*) wire signed [8:0] C311O;
(*DONT_TOUCH="true"*) wire A311O;
(*DONT_TOUCH="true"*) wire signed [8:0] C312O;
(*DONT_TOUCH="true"*) wire A312O;
(*DONT_TOUCH="true"*) wire signed [8:0] C320O;
(*DONT_TOUCH="true"*) wire A320O;
(*DONT_TOUCH="true"*) wire signed [8:0] C321O;
(*DONT_TOUCH="true"*) wire A321O;
(*DONT_TOUCH="true"*) wire signed [8:0] C322O;
(*DONT_TOUCH="true"*) wire A322O;
(*DONT_TOUCH="true"*) wire signed [8:0] C300P;
(*DONT_TOUCH="true"*) wire A300P;
(*DONT_TOUCH="true"*) wire signed [8:0] C301P;
(*DONT_TOUCH="true"*) wire A301P;
(*DONT_TOUCH="true"*) wire signed [8:0] C302P;
(*DONT_TOUCH="true"*) wire A302P;
(*DONT_TOUCH="true"*) wire signed [8:0] C310P;
(*DONT_TOUCH="true"*) wire A310P;
(*DONT_TOUCH="true"*) wire signed [8:0] C311P;
(*DONT_TOUCH="true"*) wire A311P;
(*DONT_TOUCH="true"*) wire signed [8:0] C312P;
(*DONT_TOUCH="true"*) wire A312P;
(*DONT_TOUCH="true"*) wire signed [8:0] C320P;
(*DONT_TOUCH="true"*) wire A320P;
(*DONT_TOUCH="true"*) wire signed [8:0] C321P;
(*DONT_TOUCH="true"*) wire A321P;
(*DONT_TOUCH="true"*) wire signed [8:0] C322P;
(*DONT_TOUCH="true"*) wire A322P;
(*DONT_TOUCH="true"*) wire signed [8:0] C300Q;
(*DONT_TOUCH="true"*) wire A300Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C301Q;
(*DONT_TOUCH="true"*) wire A301Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C302Q;
(*DONT_TOUCH="true"*) wire A302Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C310Q;
(*DONT_TOUCH="true"*) wire A310Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C311Q;
(*DONT_TOUCH="true"*) wire A311Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C312Q;
(*DONT_TOUCH="true"*) wire A312Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C320Q;
(*DONT_TOUCH="true"*) wire A320Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C321Q;
(*DONT_TOUCH="true"*) wire A321Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C322Q;
(*DONT_TOUCH="true"*) wire A322Q;
(*DONT_TOUCH="true"*) wire signed [8:0] C300R;
(*DONT_TOUCH="true"*) wire A300R;
(*DONT_TOUCH="true"*) wire signed [8:0] C301R;
(*DONT_TOUCH="true"*) wire A301R;
(*DONT_TOUCH="true"*) wire signed [8:0] C302R;
(*DONT_TOUCH="true"*) wire A302R;
(*DONT_TOUCH="true"*) wire signed [8:0] C310R;
(*DONT_TOUCH="true"*) wire A310R;
(*DONT_TOUCH="true"*) wire signed [8:0] C311R;
(*DONT_TOUCH="true"*) wire A311R;
(*DONT_TOUCH="true"*) wire signed [8:0] C312R;
(*DONT_TOUCH="true"*) wire A312R;
(*DONT_TOUCH="true"*) wire signed [8:0] C320R;
(*DONT_TOUCH="true"*) wire A320R;
(*DONT_TOUCH="true"*) wire signed [8:0] C321R;
(*DONT_TOUCH="true"*) wire A321R;
(*DONT_TOUCH="true"*) wire signed [8:0] C322R;
(*DONT_TOUCH="true"*) wire A322R;
(*DONT_TOUCH="true"*) wire signed [8:0] C300S;
(*DONT_TOUCH="true"*) wire A300S;
(*DONT_TOUCH="true"*) wire signed [8:0] C301S;
(*DONT_TOUCH="true"*) wire A301S;
(*DONT_TOUCH="true"*) wire signed [8:0] C302S;
(*DONT_TOUCH="true"*) wire A302S;
(*DONT_TOUCH="true"*) wire signed [8:0] C310S;
(*DONT_TOUCH="true"*) wire A310S;
(*DONT_TOUCH="true"*) wire signed [8:0] C311S;
(*DONT_TOUCH="true"*) wire A311S;
(*DONT_TOUCH="true"*) wire signed [8:0] C312S;
(*DONT_TOUCH="true"*) wire A312S;
(*DONT_TOUCH="true"*) wire signed [8:0] C320S;
(*DONT_TOUCH="true"*) wire A320S;
(*DONT_TOUCH="true"*) wire signed [8:0] C321S;
(*DONT_TOUCH="true"*) wire A321S;
(*DONT_TOUCH="true"*) wire signed [8:0] C322S;
(*DONT_TOUCH="true"*) wire A322S;
(*DONT_TOUCH="true"*) wire signed [8:0] C300T;
(*DONT_TOUCH="true"*) wire A300T;
(*DONT_TOUCH="true"*) wire signed [8:0] C301T;
(*DONT_TOUCH="true"*) wire A301T;
(*DONT_TOUCH="true"*) wire signed [8:0] C302T;
(*DONT_TOUCH="true"*) wire A302T;
(*DONT_TOUCH="true"*) wire signed [8:0] C310T;
(*DONT_TOUCH="true"*) wire A310T;
(*DONT_TOUCH="true"*) wire signed [8:0] C311T;
(*DONT_TOUCH="true"*) wire A311T;
(*DONT_TOUCH="true"*) wire signed [8:0] C312T;
(*DONT_TOUCH="true"*) wire A312T;
(*DONT_TOUCH="true"*) wire signed [8:0] C320T;
(*DONT_TOUCH="true"*) wire A320T;
(*DONT_TOUCH="true"*) wire signed [8:0] C321T;
(*DONT_TOUCH="true"*) wire A321T;
(*DONT_TOUCH="true"*) wire signed [8:0] C322T;
(*DONT_TOUCH="true"*) wire A322T;
(*DONT_TOUCH="true"*) wire signed [8:0] C300U;
(*DONT_TOUCH="true"*) wire A300U;
(*DONT_TOUCH="true"*) wire signed [8:0] C301U;
(*DONT_TOUCH="true"*) wire A301U;
(*DONT_TOUCH="true"*) wire signed [8:0] C302U;
(*DONT_TOUCH="true"*) wire A302U;
(*DONT_TOUCH="true"*) wire signed [8:0] C310U;
(*DONT_TOUCH="true"*) wire A310U;
(*DONT_TOUCH="true"*) wire signed [8:0] C311U;
(*DONT_TOUCH="true"*) wire A311U;
(*DONT_TOUCH="true"*) wire signed [8:0] C312U;
(*DONT_TOUCH="true"*) wire A312U;
(*DONT_TOUCH="true"*) wire signed [8:0] C320U;
(*DONT_TOUCH="true"*) wire A320U;
(*DONT_TOUCH="true"*) wire signed [8:0] C321U;
(*DONT_TOUCH="true"*) wire A321U;
(*DONT_TOUCH="true"*) wire signed [8:0] C322U;
(*DONT_TOUCH="true"*) wire A322U;
(*DONT_TOUCH="true"*) wire signed [8:0] C300V;
(*DONT_TOUCH="true"*) wire A300V;
(*DONT_TOUCH="true"*) wire signed [8:0] C301V;
(*DONT_TOUCH="true"*) wire A301V;
(*DONT_TOUCH="true"*) wire signed [8:0] C302V;
(*DONT_TOUCH="true"*) wire A302V;
(*DONT_TOUCH="true"*) wire signed [8:0] C310V;
(*DONT_TOUCH="true"*) wire A310V;
(*DONT_TOUCH="true"*) wire signed [8:0] C311V;
(*DONT_TOUCH="true"*) wire A311V;
(*DONT_TOUCH="true"*) wire signed [8:0] C312V;
(*DONT_TOUCH="true"*) wire A312V;
(*DONT_TOUCH="true"*) wire signed [8:0] C320V;
(*DONT_TOUCH="true"*) wire A320V;
(*DONT_TOUCH="true"*) wire signed [8:0] C321V;
(*DONT_TOUCH="true"*) wire A321V;
(*DONT_TOUCH="true"*) wire signed [8:0] C322V;
(*DONT_TOUCH="true"*) wire A322V;
DFF_save_fm DFF_W1152(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30000));
DFF_save_fm DFF_W1153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30010));
DFF_save_fm DFF_W1154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30020));
DFF_save_fm DFF_W1155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30100));
DFF_save_fm DFF_W1156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30110));
DFF_save_fm DFF_W1157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30120));
DFF_save_fm DFF_W1158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30200));
DFF_save_fm DFF_W1159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30210));
DFF_save_fm DFF_W1160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30220));
DFF_save_fm DFF_W1161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30001));
DFF_save_fm DFF_W1162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30011));
DFF_save_fm DFF_W1163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30021));
DFF_save_fm DFF_W1164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30101));
DFF_save_fm DFF_W1165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30111));
DFF_save_fm DFF_W1166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30121));
DFF_save_fm DFF_W1167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30201));
DFF_save_fm DFF_W1168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30211));
DFF_save_fm DFF_W1169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30221));
DFF_save_fm DFF_W1170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30002));
DFF_save_fm DFF_W1171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30012));
DFF_save_fm DFF_W1172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30022));
DFF_save_fm DFF_W1173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30102));
DFF_save_fm DFF_W1174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30112));
DFF_save_fm DFF_W1175(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30122));
DFF_save_fm DFF_W1176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30202));
DFF_save_fm DFF_W1177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30212));
DFF_save_fm DFF_W1178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30222));
DFF_save_fm DFF_W1179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30003));
DFF_save_fm DFF_W1180(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30013));
DFF_save_fm DFF_W1181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30023));
DFF_save_fm DFF_W1182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30103));
DFF_save_fm DFF_W1183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30113));
DFF_save_fm DFF_W1184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30123));
DFF_save_fm DFF_W1185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30203));
DFF_save_fm DFF_W1186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30213));
DFF_save_fm DFF_W1187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30223));
DFF_save_fm DFF_W1188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30004));
DFF_save_fm DFF_W1189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30014));
DFF_save_fm DFF_W1190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30024));
DFF_save_fm DFF_W1191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30104));
DFF_save_fm DFF_W1192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30114));
DFF_save_fm DFF_W1193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30124));
DFF_save_fm DFF_W1194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30204));
DFF_save_fm DFF_W1195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30214));
DFF_save_fm DFF_W1196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30224));
DFF_save_fm DFF_W1197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30005));
DFF_save_fm DFF_W1198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30015));
DFF_save_fm DFF_W1199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30025));
DFF_save_fm DFF_W1200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30105));
DFF_save_fm DFF_W1201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30115));
DFF_save_fm DFF_W1202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30125));
DFF_save_fm DFF_W1203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30205));
DFF_save_fm DFF_W1204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30215));
DFF_save_fm DFF_W1205(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30225));
DFF_save_fm DFF_W1206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30006));
DFF_save_fm DFF_W1207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30016));
DFF_save_fm DFF_W1208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30026));
DFF_save_fm DFF_W1209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30106));
DFF_save_fm DFF_W1210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30116));
DFF_save_fm DFF_W1211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30126));
DFF_save_fm DFF_W1212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30206));
DFF_save_fm DFF_W1213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30216));
DFF_save_fm DFF_W1214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30226));
DFF_save_fm DFF_W1215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30007));
DFF_save_fm DFF_W1216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30017));
DFF_save_fm DFF_W1217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30027));
DFF_save_fm DFF_W1218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30107));
DFF_save_fm DFF_W1219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30117));
DFF_save_fm DFF_W1220(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30127));
DFF_save_fm DFF_W1221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30207));
DFF_save_fm DFF_W1222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30217));
DFF_save_fm DFF_W1223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30227));
DFF_save_fm DFF_W1224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30008));
DFF_save_fm DFF_W1225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30018));
DFF_save_fm DFF_W1226(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30028));
DFF_save_fm DFF_W1227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30108));
DFF_save_fm DFF_W1228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30118));
DFF_save_fm DFF_W1229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30128));
DFF_save_fm DFF_W1230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30208));
DFF_save_fm DFF_W1231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30218));
DFF_save_fm DFF_W1232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30228));
DFF_save_fm DFF_W1233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30009));
DFF_save_fm DFF_W1234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30019));
DFF_save_fm DFF_W1235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30029));
DFF_save_fm DFF_W1236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30109));
DFF_save_fm DFF_W1237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30119));
DFF_save_fm DFF_W1238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30129));
DFF_save_fm DFF_W1239(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30209));
DFF_save_fm DFF_W1240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30219));
DFF_save_fm DFF_W1241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30229));
DFF_save_fm DFF_W1242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000A));
DFF_save_fm DFF_W1243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001A));
DFF_save_fm DFF_W1244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002A));
DFF_save_fm DFF_W1245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010A));
DFF_save_fm DFF_W1246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011A));
DFF_save_fm DFF_W1247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012A));
DFF_save_fm DFF_W1248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020A));
DFF_save_fm DFF_W1249(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021A));
DFF_save_fm DFF_W1250(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022A));
DFF_save_fm DFF_W1251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000B));
DFF_save_fm DFF_W1252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001B));
DFF_save_fm DFF_W1253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002B));
DFF_save_fm DFF_W1254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010B));
DFF_save_fm DFF_W1255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011B));
DFF_save_fm DFF_W1256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012B));
DFF_save_fm DFF_W1257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020B));
DFF_save_fm DFF_W1258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021B));
DFF_save_fm DFF_W1259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022B));
DFF_save_fm DFF_W1260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000C));
DFF_save_fm DFF_W1261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001C));
DFF_save_fm DFF_W1262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002C));
DFF_save_fm DFF_W1263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010C));
DFF_save_fm DFF_W1264(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011C));
DFF_save_fm DFF_W1265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012C));
DFF_save_fm DFF_W1266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020C));
DFF_save_fm DFF_W1267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021C));
DFF_save_fm DFF_W1268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022C));
DFF_save_fm DFF_W1269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000D));
DFF_save_fm DFF_W1270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001D));
DFF_save_fm DFF_W1271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002D));
DFF_save_fm DFF_W1272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010D));
DFF_save_fm DFF_W1273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011D));
DFF_save_fm DFF_W1274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012D));
DFF_save_fm DFF_W1275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020D));
DFF_save_fm DFF_W1276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021D));
DFF_save_fm DFF_W1277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022D));
DFF_save_fm DFF_W1278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000E));
DFF_save_fm DFF_W1279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001E));
DFF_save_fm DFF_W1280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002E));
DFF_save_fm DFF_W1281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010E));
DFF_save_fm DFF_W1282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011E));
DFF_save_fm DFF_W1283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012E));
DFF_save_fm DFF_W1284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020E));
DFF_save_fm DFF_W1285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021E));
DFF_save_fm DFF_W1286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022E));
DFF_save_fm DFF_W1287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000F));
DFF_save_fm DFF_W1288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001F));
DFF_save_fm DFF_W1289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002F));
DFF_save_fm DFF_W1290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010F));
DFF_save_fm DFF_W1291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011F));
DFF_save_fm DFF_W1292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012F));
DFF_save_fm DFF_W1293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020F));
DFF_save_fm DFF_W1294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021F));
DFF_save_fm DFF_W1295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022F));
DFF_save_fm DFF_W1296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31000));
DFF_save_fm DFF_W1297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31010));
DFF_save_fm DFF_W1298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31020));
DFF_save_fm DFF_W1299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31100));
DFF_save_fm DFF_W1300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31110));
DFF_save_fm DFF_W1301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31120));
DFF_save_fm DFF_W1302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31200));
DFF_save_fm DFF_W1303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31210));
DFF_save_fm DFF_W1304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31220));
DFF_save_fm DFF_W1305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31001));
DFF_save_fm DFF_W1306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31011));
DFF_save_fm DFF_W1307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31021));
DFF_save_fm DFF_W1308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31101));
DFF_save_fm DFF_W1309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31111));
DFF_save_fm DFF_W1310(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31121));
DFF_save_fm DFF_W1311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31201));
DFF_save_fm DFF_W1312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31211));
DFF_save_fm DFF_W1313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31221));
DFF_save_fm DFF_W1314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31002));
DFF_save_fm DFF_W1315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31012));
DFF_save_fm DFF_W1316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31022));
DFF_save_fm DFF_W1317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31102));
DFF_save_fm DFF_W1318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31112));
DFF_save_fm DFF_W1319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31122));
DFF_save_fm DFF_W1320(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31202));
DFF_save_fm DFF_W1321(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31212));
DFF_save_fm DFF_W1322(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31222));
DFF_save_fm DFF_W1323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31003));
DFF_save_fm DFF_W1324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31013));
DFF_save_fm DFF_W1325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31023));
DFF_save_fm DFF_W1326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31103));
DFF_save_fm DFF_W1327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31113));
DFF_save_fm DFF_W1328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31123));
DFF_save_fm DFF_W1329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31203));
DFF_save_fm DFF_W1330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31213));
DFF_save_fm DFF_W1331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31223));
DFF_save_fm DFF_W1332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31004));
DFF_save_fm DFF_W1333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31014));
DFF_save_fm DFF_W1334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31024));
DFF_save_fm DFF_W1335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31104));
DFF_save_fm DFF_W1336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31114));
DFF_save_fm DFF_W1337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31124));
DFF_save_fm DFF_W1338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31204));
DFF_save_fm DFF_W1339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31214));
DFF_save_fm DFF_W1340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31224));
DFF_save_fm DFF_W1341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31005));
DFF_save_fm DFF_W1342(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31015));
DFF_save_fm DFF_W1343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31025));
DFF_save_fm DFF_W1344(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31105));
DFF_save_fm DFF_W1345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31115));
DFF_save_fm DFF_W1346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31125));
DFF_save_fm DFF_W1347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31205));
DFF_save_fm DFF_W1348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31215));
DFF_save_fm DFF_W1349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31225));
DFF_save_fm DFF_W1350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31006));
DFF_save_fm DFF_W1351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31016));
DFF_save_fm DFF_W1352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31026));
DFF_save_fm DFF_W1353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31106));
DFF_save_fm DFF_W1354(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31116));
DFF_save_fm DFF_W1355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31126));
DFF_save_fm DFF_W1356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31206));
DFF_save_fm DFF_W1357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31216));
DFF_save_fm DFF_W1358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31226));
DFF_save_fm DFF_W1359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31007));
DFF_save_fm DFF_W1360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31017));
DFF_save_fm DFF_W1361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31027));
DFF_save_fm DFF_W1362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31107));
DFF_save_fm DFF_W1363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31117));
DFF_save_fm DFF_W1364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31127));
DFF_save_fm DFF_W1365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31207));
DFF_save_fm DFF_W1366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31217));
DFF_save_fm DFF_W1367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31227));
DFF_save_fm DFF_W1368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31008));
DFF_save_fm DFF_W1369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31018));
DFF_save_fm DFF_W1370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31028));
DFF_save_fm DFF_W1371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31108));
DFF_save_fm DFF_W1372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31118));
DFF_save_fm DFF_W1373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31128));
DFF_save_fm DFF_W1374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31208));
DFF_save_fm DFF_W1375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31218));
DFF_save_fm DFF_W1376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31228));
DFF_save_fm DFF_W1377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31009));
DFF_save_fm DFF_W1378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31019));
DFF_save_fm DFF_W1379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31029));
DFF_save_fm DFF_W1380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31109));
DFF_save_fm DFF_W1381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31119));
DFF_save_fm DFF_W1382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31129));
DFF_save_fm DFF_W1383(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31209));
DFF_save_fm DFF_W1384(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31219));
DFF_save_fm DFF_W1385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31229));
DFF_save_fm DFF_W1386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100A));
DFF_save_fm DFF_W1387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101A));
DFF_save_fm DFF_W1388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102A));
DFF_save_fm DFF_W1389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110A));
DFF_save_fm DFF_W1390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111A));
DFF_save_fm DFF_W1391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112A));
DFF_save_fm DFF_W1392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120A));
DFF_save_fm DFF_W1393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121A));
DFF_save_fm DFF_W1394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122A));
DFF_save_fm DFF_W1395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100B));
DFF_save_fm DFF_W1396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101B));
DFF_save_fm DFF_W1397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102B));
DFF_save_fm DFF_W1398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110B));
DFF_save_fm DFF_W1399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111B));
DFF_save_fm DFF_W1400(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112B));
DFF_save_fm DFF_W1401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120B));
DFF_save_fm DFF_W1402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121B));
DFF_save_fm DFF_W1403(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122B));
DFF_save_fm DFF_W1404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100C));
DFF_save_fm DFF_W1405(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101C));
DFF_save_fm DFF_W1406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102C));
DFF_save_fm DFF_W1407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110C));
DFF_save_fm DFF_W1408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111C));
DFF_save_fm DFF_W1409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112C));
DFF_save_fm DFF_W1410(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120C));
DFF_save_fm DFF_W1411(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121C));
DFF_save_fm DFF_W1412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122C));
DFF_save_fm DFF_W1413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100D));
DFF_save_fm DFF_W1414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101D));
DFF_save_fm DFF_W1415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102D));
DFF_save_fm DFF_W1416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110D));
DFF_save_fm DFF_W1417(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111D));
DFF_save_fm DFF_W1418(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112D));
DFF_save_fm DFF_W1419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120D));
DFF_save_fm DFF_W1420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121D));
DFF_save_fm DFF_W1421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122D));
DFF_save_fm DFF_W1422(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100E));
DFF_save_fm DFF_W1423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101E));
DFF_save_fm DFF_W1424(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102E));
DFF_save_fm DFF_W1425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110E));
DFF_save_fm DFF_W1426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111E));
DFF_save_fm DFF_W1427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112E));
DFF_save_fm DFF_W1428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120E));
DFF_save_fm DFF_W1429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121E));
DFF_save_fm DFF_W1430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122E));
DFF_save_fm DFF_W1431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100F));
DFF_save_fm DFF_W1432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101F));
DFF_save_fm DFF_W1433(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102F));
DFF_save_fm DFF_W1434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110F));
DFF_save_fm DFF_W1435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111F));
DFF_save_fm DFF_W1436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112F));
DFF_save_fm DFF_W1437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120F));
DFF_save_fm DFF_W1438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121F));
DFF_save_fm DFF_W1439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122F));
DFF_save_fm DFF_W1440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32000));
DFF_save_fm DFF_W1441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32010));
DFF_save_fm DFF_W1442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32020));
DFF_save_fm DFF_W1443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32100));
DFF_save_fm DFF_W1444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32110));
DFF_save_fm DFF_W1445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32120));
DFF_save_fm DFF_W1446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32200));
DFF_save_fm DFF_W1447(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32210));
DFF_save_fm DFF_W1448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32220));
DFF_save_fm DFF_W1449(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32001));
DFF_save_fm DFF_W1450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32011));
DFF_save_fm DFF_W1451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32021));
DFF_save_fm DFF_W1452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32101));
DFF_save_fm DFF_W1453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32111));
DFF_save_fm DFF_W1454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32121));
DFF_save_fm DFF_W1455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32201));
DFF_save_fm DFF_W1456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32211));
DFF_save_fm DFF_W1457(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32221));
DFF_save_fm DFF_W1458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32002));
DFF_save_fm DFF_W1459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32012));
DFF_save_fm DFF_W1460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32022));
DFF_save_fm DFF_W1461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32102));
DFF_save_fm DFF_W1462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32112));
DFF_save_fm DFF_W1463(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32122));
DFF_save_fm DFF_W1464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32202));
DFF_save_fm DFF_W1465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32212));
DFF_save_fm DFF_W1466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32222));
DFF_save_fm DFF_W1467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32003));
DFF_save_fm DFF_W1468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32013));
DFF_save_fm DFF_W1469(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32023));
DFF_save_fm DFF_W1470(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32103));
DFF_save_fm DFF_W1471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32113));
DFF_save_fm DFF_W1472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32123));
DFF_save_fm DFF_W1473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32203));
DFF_save_fm DFF_W1474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32213));
DFF_save_fm DFF_W1475(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32223));
DFF_save_fm DFF_W1476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32004));
DFF_save_fm DFF_W1477(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32014));
DFF_save_fm DFF_W1478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32024));
DFF_save_fm DFF_W1479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32104));
DFF_save_fm DFF_W1480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32114));
DFF_save_fm DFF_W1481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32124));
DFF_save_fm DFF_W1482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32204));
DFF_save_fm DFF_W1483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32214));
DFF_save_fm DFF_W1484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32224));
DFF_save_fm DFF_W1485(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32005));
DFF_save_fm DFF_W1486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32015));
DFF_save_fm DFF_W1487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32025));
DFF_save_fm DFF_W1488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32105));
DFF_save_fm DFF_W1489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32115));
DFF_save_fm DFF_W1490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32125));
DFF_save_fm DFF_W1491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32205));
DFF_save_fm DFF_W1492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32215));
DFF_save_fm DFF_W1493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32225));
DFF_save_fm DFF_W1494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32006));
DFF_save_fm DFF_W1495(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32016));
DFF_save_fm DFF_W1496(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32026));
DFF_save_fm DFF_W1497(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32106));
DFF_save_fm DFF_W1498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32116));
DFF_save_fm DFF_W1499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32126));
DFF_save_fm DFF_W1500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32206));
DFF_save_fm DFF_W1501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32216));
DFF_save_fm DFF_W1502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32226));
DFF_save_fm DFF_W1503(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32007));
DFF_save_fm DFF_W1504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32017));
DFF_save_fm DFF_W1505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32027));
DFF_save_fm DFF_W1506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32107));
DFF_save_fm DFF_W1507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32117));
DFF_save_fm DFF_W1508(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32127));
DFF_save_fm DFF_W1509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32207));
DFF_save_fm DFF_W1510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32217));
DFF_save_fm DFF_W1511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32227));
DFF_save_fm DFF_W1512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32008));
DFF_save_fm DFF_W1513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32018));
DFF_save_fm DFF_W1514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32028));
DFF_save_fm DFF_W1515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32108));
DFF_save_fm DFF_W1516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32118));
DFF_save_fm DFF_W1517(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32128));
DFF_save_fm DFF_W1518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32208));
DFF_save_fm DFF_W1519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32218));
DFF_save_fm DFF_W1520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32228));
DFF_save_fm DFF_W1521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32009));
DFF_save_fm DFF_W1522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32019));
DFF_save_fm DFF_W1523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32029));
DFF_save_fm DFF_W1524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32109));
DFF_save_fm DFF_W1525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32119));
DFF_save_fm DFF_W1526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W32129));
DFF_save_fm DFF_W1527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32209));
DFF_save_fm DFF_W1528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32219));
DFF_save_fm DFF_W1529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W32229));
DFF_save_fm DFF_W1530(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3200A));
DFF_save_fm DFF_W1531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3201A));
DFF_save_fm DFF_W1532(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3202A));
DFF_save_fm DFF_W1533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3210A));
DFF_save_fm DFF_W1534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3211A));
DFF_save_fm DFF_W1535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3212A));
DFF_save_fm DFF_W1536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3220A));
DFF_save_fm DFF_W1537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3221A));
DFF_save_fm DFF_W1538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3222A));
DFF_save_fm DFF_W1539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3200B));
DFF_save_fm DFF_W1540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3201B));
DFF_save_fm DFF_W1541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3202B));
DFF_save_fm DFF_W1542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3210B));
DFF_save_fm DFF_W1543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3211B));
DFF_save_fm DFF_W1544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3212B));
DFF_save_fm DFF_W1545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3220B));
DFF_save_fm DFF_W1546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3221B));
DFF_save_fm DFF_W1547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3222B));
DFF_save_fm DFF_W1548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3200C));
DFF_save_fm DFF_W1549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3201C));
DFF_save_fm DFF_W1550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3202C));
DFF_save_fm DFF_W1551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3210C));
DFF_save_fm DFF_W1552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3211C));
DFF_save_fm DFF_W1553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3212C));
DFF_save_fm DFF_W1554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3220C));
DFF_save_fm DFF_W1555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3221C));
DFF_save_fm DFF_W1556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3222C));
DFF_save_fm DFF_W1557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3200D));
DFF_save_fm DFF_W1558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3201D));
DFF_save_fm DFF_W1559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3202D));
DFF_save_fm DFF_W1560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3210D));
DFF_save_fm DFF_W1561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3211D));
DFF_save_fm DFF_W1562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3212D));
DFF_save_fm DFF_W1563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3220D));
DFF_save_fm DFF_W1564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3221D));
DFF_save_fm DFF_W1565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3222D));
DFF_save_fm DFF_W1566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3200E));
DFF_save_fm DFF_W1567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3201E));
DFF_save_fm DFF_W1568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3202E));
DFF_save_fm DFF_W1569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3210E));
DFF_save_fm DFF_W1570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3211E));
DFF_save_fm DFF_W1571(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3212E));
DFF_save_fm DFF_W1572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3220E));
DFF_save_fm DFF_W1573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3221E));
DFF_save_fm DFF_W1574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3222E));
DFF_save_fm DFF_W1575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3200F));
DFF_save_fm DFF_W1576(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3201F));
DFF_save_fm DFF_W1577(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3202F));
DFF_save_fm DFF_W1578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3210F));
DFF_save_fm DFF_W1579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3211F));
DFF_save_fm DFF_W1580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3212F));
DFF_save_fm DFF_W1581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3220F));
DFF_save_fm DFF_W1582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3221F));
DFF_save_fm DFF_W1583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3222F));
DFF_save_fm DFF_W1584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33000));
DFF_save_fm DFF_W1585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33010));
DFF_save_fm DFF_W1586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33020));
DFF_save_fm DFF_W1587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33100));
DFF_save_fm DFF_W1588(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33110));
DFF_save_fm DFF_W1589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33120));
DFF_save_fm DFF_W1590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33200));
DFF_save_fm DFF_W1591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33210));
DFF_save_fm DFF_W1592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33220));
DFF_save_fm DFF_W1593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33001));
DFF_save_fm DFF_W1594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33011));
DFF_save_fm DFF_W1595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33021));
DFF_save_fm DFF_W1596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33101));
DFF_save_fm DFF_W1597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33111));
DFF_save_fm DFF_W1598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33121));
DFF_save_fm DFF_W1599(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33201));
DFF_save_fm DFF_W1600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33211));
DFF_save_fm DFF_W1601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33221));
DFF_save_fm DFF_W1602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33002));
DFF_save_fm DFF_W1603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33012));
DFF_save_fm DFF_W1604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33022));
DFF_save_fm DFF_W1605(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33102));
DFF_save_fm DFF_W1606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33112));
DFF_save_fm DFF_W1607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33122));
DFF_save_fm DFF_W1608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33202));
DFF_save_fm DFF_W1609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33212));
DFF_save_fm DFF_W1610(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33222));
DFF_save_fm DFF_W1611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33003));
DFF_save_fm DFF_W1612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33013));
DFF_save_fm DFF_W1613(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33023));
DFF_save_fm DFF_W1614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33103));
DFF_save_fm DFF_W1615(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33113));
DFF_save_fm DFF_W1616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33123));
DFF_save_fm DFF_W1617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33203));
DFF_save_fm DFF_W1618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33213));
DFF_save_fm DFF_W1619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33223));
DFF_save_fm DFF_W1620(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33004));
DFF_save_fm DFF_W1621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33014));
DFF_save_fm DFF_W1622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33024));
DFF_save_fm DFF_W1623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33104));
DFF_save_fm DFF_W1624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33114));
DFF_save_fm DFF_W1625(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33124));
DFF_save_fm DFF_W1626(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33204));
DFF_save_fm DFF_W1627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33214));
DFF_save_fm DFF_W1628(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33224));
DFF_save_fm DFF_W1629(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33005));
DFF_save_fm DFF_W1630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33015));
DFF_save_fm DFF_W1631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33025));
DFF_save_fm DFF_W1632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33105));
DFF_save_fm DFF_W1633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33115));
DFF_save_fm DFF_W1634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33125));
DFF_save_fm DFF_W1635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33205));
DFF_save_fm DFF_W1636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33215));
DFF_save_fm DFF_W1637(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33225));
DFF_save_fm DFF_W1638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33006));
DFF_save_fm DFF_W1639(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33016));
DFF_save_fm DFF_W1640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33026));
DFF_save_fm DFF_W1641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33106));
DFF_save_fm DFF_W1642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33116));
DFF_save_fm DFF_W1643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33126));
DFF_save_fm DFF_W1644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33206));
DFF_save_fm DFF_W1645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33216));
DFF_save_fm DFF_W1646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33226));
DFF_save_fm DFF_W1647(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33007));
DFF_save_fm DFF_W1648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33017));
DFF_save_fm DFF_W1649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33027));
DFF_save_fm DFF_W1650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33107));
DFF_save_fm DFF_W1651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33117));
DFF_save_fm DFF_W1652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33127));
DFF_save_fm DFF_W1653(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33207));
DFF_save_fm DFF_W1654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33217));
DFF_save_fm DFF_W1655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33227));
DFF_save_fm DFF_W1656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33008));
DFF_save_fm DFF_W1657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33018));
DFF_save_fm DFF_W1658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33028));
DFF_save_fm DFF_W1659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33108));
DFF_save_fm DFF_W1660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33118));
DFF_save_fm DFF_W1661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33128));
DFF_save_fm DFF_W1662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33208));
DFF_save_fm DFF_W1663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33218));
DFF_save_fm DFF_W1664(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33228));
DFF_save_fm DFF_W1665(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33009));
DFF_save_fm DFF_W1666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33019));
DFF_save_fm DFF_W1667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33029));
DFF_save_fm DFF_W1668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33109));
DFF_save_fm DFF_W1669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33119));
DFF_save_fm DFF_W1670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33129));
DFF_save_fm DFF_W1671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W33209));
DFF_save_fm DFF_W1672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33219));
DFF_save_fm DFF_W1673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W33229));
DFF_save_fm DFF_W1674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3300A));
DFF_save_fm DFF_W1675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3301A));
DFF_save_fm DFF_W1676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3302A));
DFF_save_fm DFF_W1677(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3310A));
DFF_save_fm DFF_W1678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3311A));
DFF_save_fm DFF_W1679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3312A));
DFF_save_fm DFF_W1680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3320A));
DFF_save_fm DFF_W1681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3321A));
DFF_save_fm DFF_W1682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3322A));
DFF_save_fm DFF_W1683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3300B));
DFF_save_fm DFF_W1684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3301B));
DFF_save_fm DFF_W1685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3302B));
DFF_save_fm DFF_W1686(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3310B));
DFF_save_fm DFF_W1687(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3311B));
DFF_save_fm DFF_W1688(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3312B));
DFF_save_fm DFF_W1689(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3320B));
DFF_save_fm DFF_W1690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3321B));
DFF_save_fm DFF_W1691(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3322B));
DFF_save_fm DFF_W1692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3300C));
DFF_save_fm DFF_W1693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3301C));
DFF_save_fm DFF_W1694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3302C));
DFF_save_fm DFF_W1695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3310C));
DFF_save_fm DFF_W1696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3311C));
DFF_save_fm DFF_W1697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3312C));
DFF_save_fm DFF_W1698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3320C));
DFF_save_fm DFF_W1699(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3321C));
DFF_save_fm DFF_W1700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3322C));
DFF_save_fm DFF_W1701(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3300D));
DFF_save_fm DFF_W1702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3301D));
DFF_save_fm DFF_W1703(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3302D));
DFF_save_fm DFF_W1704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3310D));
DFF_save_fm DFF_W1705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3311D));
DFF_save_fm DFF_W1706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3312D));
DFF_save_fm DFF_W1707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3320D));
DFF_save_fm DFF_W1708(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3321D));
DFF_save_fm DFF_W1709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3322D));
DFF_save_fm DFF_W1710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3300E));
DFF_save_fm DFF_W1711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3301E));
DFF_save_fm DFF_W1712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3302E));
DFF_save_fm DFF_W1713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3310E));
DFF_save_fm DFF_W1714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3311E));
DFF_save_fm DFF_W1715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3312E));
DFF_save_fm DFF_W1716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3320E));
DFF_save_fm DFF_W1717(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3321E));
DFF_save_fm DFF_W1718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3322E));
DFF_save_fm DFF_W1719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3300F));
DFF_save_fm DFF_W1720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3301F));
DFF_save_fm DFF_W1721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3302F));
DFF_save_fm DFF_W1722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3310F));
DFF_save_fm DFF_W1723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3311F));
DFF_save_fm DFF_W1724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3312F));
DFF_save_fm DFF_W1725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3320F));
DFF_save_fm DFF_W1726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3321F));
DFF_save_fm DFF_W1727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3322F));
DFF_save_fm DFF_W1728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34000));
DFF_save_fm DFF_W1729(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34010));
DFF_save_fm DFF_W1730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34020));
DFF_save_fm DFF_W1731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34100));
DFF_save_fm DFF_W1732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34110));
DFF_save_fm DFF_W1733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34120));
DFF_save_fm DFF_W1734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34200));
DFF_save_fm DFF_W1735(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34210));
DFF_save_fm DFF_W1736(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34220));
DFF_save_fm DFF_W1737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34001));
DFF_save_fm DFF_W1738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34011));
DFF_save_fm DFF_W1739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34021));
DFF_save_fm DFF_W1740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34101));
DFF_save_fm DFF_W1741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34111));
DFF_save_fm DFF_W1742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34121));
DFF_save_fm DFF_W1743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34201));
DFF_save_fm DFF_W1744(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34211));
DFF_save_fm DFF_W1745(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34221));
DFF_save_fm DFF_W1746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34002));
DFF_save_fm DFF_W1747(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34012));
DFF_save_fm DFF_W1748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34022));
DFF_save_fm DFF_W1749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34102));
DFF_save_fm DFF_W1750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34112));
DFF_save_fm DFF_W1751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34122));
DFF_save_fm DFF_W1752(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34202));
DFF_save_fm DFF_W1753(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34212));
DFF_save_fm DFF_W1754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34222));
DFF_save_fm DFF_W1755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34003));
DFF_save_fm DFF_W1756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34013));
DFF_save_fm DFF_W1757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34023));
DFF_save_fm DFF_W1758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34103));
DFF_save_fm DFF_W1759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34113));
DFF_save_fm DFF_W1760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34123));
DFF_save_fm DFF_W1761(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34203));
DFF_save_fm DFF_W1762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34213));
DFF_save_fm DFF_W1763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34223));
DFF_save_fm DFF_W1764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34004));
DFF_save_fm DFF_W1765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34014));
DFF_save_fm DFF_W1766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34024));
DFF_save_fm DFF_W1767(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34104));
DFF_save_fm DFF_W1768(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34114));
DFF_save_fm DFF_W1769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34124));
DFF_save_fm DFF_W1770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34204));
DFF_save_fm DFF_W1771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34214));
DFF_save_fm DFF_W1772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34224));
DFF_save_fm DFF_W1773(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34005));
DFF_save_fm DFF_W1774(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34015));
DFF_save_fm DFF_W1775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34025));
DFF_save_fm DFF_W1776(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34105));
DFF_save_fm DFF_W1777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34115));
DFF_save_fm DFF_W1778(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34125));
DFF_save_fm DFF_W1779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34205));
DFF_save_fm DFF_W1780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34215));
DFF_save_fm DFF_W1781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34225));
DFF_save_fm DFF_W1782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34006));
DFF_save_fm DFF_W1783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34016));
DFF_save_fm DFF_W1784(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34026));
DFF_save_fm DFF_W1785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34106));
DFF_save_fm DFF_W1786(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34116));
DFF_save_fm DFF_W1787(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34126));
DFF_save_fm DFF_W1788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34206));
DFF_save_fm DFF_W1789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34216));
DFF_save_fm DFF_W1790(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34226));
DFF_save_fm DFF_W1791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34007));
DFF_save_fm DFF_W1792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34017));
DFF_save_fm DFF_W1793(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34027));
DFF_save_fm DFF_W1794(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34107));
DFF_save_fm DFF_W1795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34117));
DFF_save_fm DFF_W1796(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34127));
DFF_save_fm DFF_W1797(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34207));
DFF_save_fm DFF_W1798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34217));
DFF_save_fm DFF_W1799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34227));
DFF_save_fm DFF_W1800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34008));
DFF_save_fm DFF_W1801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34018));
DFF_save_fm DFF_W1802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34028));
DFF_save_fm DFF_W1803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34108));
DFF_save_fm DFF_W1804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34118));
DFF_save_fm DFF_W1805(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34128));
DFF_save_fm DFF_W1806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34208));
DFF_save_fm DFF_W1807(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34218));
DFF_save_fm DFF_W1808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34228));
DFF_save_fm DFF_W1809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34009));
DFF_save_fm DFF_W1810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34019));
DFF_save_fm DFF_W1811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34029));
DFF_save_fm DFF_W1812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34109));
DFF_save_fm DFF_W1813(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34119));
DFF_save_fm DFF_W1814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34129));
DFF_save_fm DFF_W1815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W34209));
DFF_save_fm DFF_W1816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34219));
DFF_save_fm DFF_W1817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W34229));
DFF_save_fm DFF_W1818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3400A));
DFF_save_fm DFF_W1819(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3401A));
DFF_save_fm DFF_W1820(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3402A));
DFF_save_fm DFF_W1821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3410A));
DFF_save_fm DFF_W1822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3411A));
DFF_save_fm DFF_W1823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3412A));
DFF_save_fm DFF_W1824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3420A));
DFF_save_fm DFF_W1825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3421A));
DFF_save_fm DFF_W1826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3422A));
DFF_save_fm DFF_W1827(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3400B));
DFF_save_fm DFF_W1828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3401B));
DFF_save_fm DFF_W1829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3402B));
DFF_save_fm DFF_W1830(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3410B));
DFF_save_fm DFF_W1831(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3411B));
DFF_save_fm DFF_W1832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3412B));
DFF_save_fm DFF_W1833(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3420B));
DFF_save_fm DFF_W1834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3421B));
DFF_save_fm DFF_W1835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3422B));
DFF_save_fm DFF_W1836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3400C));
DFF_save_fm DFF_W1837(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3401C));
DFF_save_fm DFF_W1838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3402C));
DFF_save_fm DFF_W1839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3410C));
DFF_save_fm DFF_W1840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3411C));
DFF_save_fm DFF_W1841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3412C));
DFF_save_fm DFF_W1842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3420C));
DFF_save_fm DFF_W1843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3421C));
DFF_save_fm DFF_W1844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3422C));
DFF_save_fm DFF_W1845(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3400D));
DFF_save_fm DFF_W1846(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3401D));
DFF_save_fm DFF_W1847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3402D));
DFF_save_fm DFF_W1848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3410D));
DFF_save_fm DFF_W1849(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3411D));
DFF_save_fm DFF_W1850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3412D));
DFF_save_fm DFF_W1851(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3420D));
DFF_save_fm DFF_W1852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3421D));
DFF_save_fm DFF_W1853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3422D));
DFF_save_fm DFF_W1854(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3400E));
DFF_save_fm DFF_W1855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3401E));
DFF_save_fm DFF_W1856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3402E));
DFF_save_fm DFF_W1857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3410E));
DFF_save_fm DFF_W1858(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3411E));
DFF_save_fm DFF_W1859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3412E));
DFF_save_fm DFF_W1860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3420E));
DFF_save_fm DFF_W1861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3421E));
DFF_save_fm DFF_W1862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3422E));
DFF_save_fm DFF_W1863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3400F));
DFF_save_fm DFF_W1864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3401F));
DFF_save_fm DFF_W1865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3402F));
DFF_save_fm DFF_W1866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3410F));
DFF_save_fm DFF_W1867(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3411F));
DFF_save_fm DFF_W1868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3412F));
DFF_save_fm DFF_W1869(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3420F));
DFF_save_fm DFF_W1870(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3421F));
DFF_save_fm DFF_W1871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3422F));
DFF_save_fm DFF_W1872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35000));
DFF_save_fm DFF_W1873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35010));
DFF_save_fm DFF_W1874(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35020));
DFF_save_fm DFF_W1875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35100));
DFF_save_fm DFF_W1876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35110));
DFF_save_fm DFF_W1877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35120));
DFF_save_fm DFF_W1878(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35200));
DFF_save_fm DFF_W1879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35210));
DFF_save_fm DFF_W1880(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35220));
DFF_save_fm DFF_W1881(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35001));
DFF_save_fm DFF_W1882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35011));
DFF_save_fm DFF_W1883(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35021));
DFF_save_fm DFF_W1884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35101));
DFF_save_fm DFF_W1885(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35111));
DFF_save_fm DFF_W1886(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35121));
DFF_save_fm DFF_W1887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35201));
DFF_save_fm DFF_W1888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35211));
DFF_save_fm DFF_W1889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35221));
DFF_save_fm DFF_W1890(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35002));
DFF_save_fm DFF_W1891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35012));
DFF_save_fm DFF_W1892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35022));
DFF_save_fm DFF_W1893(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35102));
DFF_save_fm DFF_W1894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35112));
DFF_save_fm DFF_W1895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35122));
DFF_save_fm DFF_W1896(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35202));
DFF_save_fm DFF_W1897(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35212));
DFF_save_fm DFF_W1898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35222));
DFF_save_fm DFF_W1899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35003));
DFF_save_fm DFF_W1900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35013));
DFF_save_fm DFF_W1901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35023));
DFF_save_fm DFF_W1902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35103));
DFF_save_fm DFF_W1903(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35113));
DFF_save_fm DFF_W1904(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35123));
DFF_save_fm DFF_W1905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35203));
DFF_save_fm DFF_W1906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35213));
DFF_save_fm DFF_W1907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35223));
DFF_save_fm DFF_W1908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35004));
DFF_save_fm DFF_W1909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35014));
DFF_save_fm DFF_W1910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35024));
DFF_save_fm DFF_W1911(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35104));
DFF_save_fm DFF_W1912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35114));
DFF_save_fm DFF_W1913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35124));
DFF_save_fm DFF_W1914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35204));
DFF_save_fm DFF_W1915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35214));
DFF_save_fm DFF_W1916(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35224));
DFF_save_fm DFF_W1917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35005));
DFF_save_fm DFF_W1918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35015));
DFF_save_fm DFF_W1919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35025));
DFF_save_fm DFF_W1920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35105));
DFF_save_fm DFF_W1921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35115));
DFF_save_fm DFF_W1922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35125));
DFF_save_fm DFF_W1923(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35205));
DFF_save_fm DFF_W1924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35215));
DFF_save_fm DFF_W1925(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35225));
DFF_save_fm DFF_W1926(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35006));
DFF_save_fm DFF_W1927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35016));
DFF_save_fm DFF_W1928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35026));
DFF_save_fm DFF_W1929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35106));
DFF_save_fm DFF_W1930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35116));
DFF_save_fm DFF_W1931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35126));
DFF_save_fm DFF_W1932(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35206));
DFF_save_fm DFF_W1933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35216));
DFF_save_fm DFF_W1934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35226));
DFF_save_fm DFF_W1935(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35007));
DFF_save_fm DFF_W1936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35017));
DFF_save_fm DFF_W1937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35027));
DFF_save_fm DFF_W1938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35107));
DFF_save_fm DFF_W1939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35117));
DFF_save_fm DFF_W1940(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35127));
DFF_save_fm DFF_W1941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35207));
DFF_save_fm DFF_W1942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35217));
DFF_save_fm DFF_W1943(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35227));
DFF_save_fm DFF_W1944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35008));
DFF_save_fm DFF_W1945(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35018));
DFF_save_fm DFF_W1946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35028));
DFF_save_fm DFF_W1947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35108));
DFF_save_fm DFF_W1948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35118));
DFF_save_fm DFF_W1949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35128));
DFF_save_fm DFF_W1950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35208));
DFF_save_fm DFF_W1951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35218));
DFF_save_fm DFF_W1952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35228));
DFF_save_fm DFF_W1953(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35009));
DFF_save_fm DFF_W1954(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35019));
DFF_save_fm DFF_W1955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35029));
DFF_save_fm DFF_W1956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35109));
DFF_save_fm DFF_W1957(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35119));
DFF_save_fm DFF_W1958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35129));
DFF_save_fm DFF_W1959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35209));
DFF_save_fm DFF_W1960(.clk(clk),.rstn(rstn),.reset_value(1),.q(W35219));
DFF_save_fm DFF_W1961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W35229));
DFF_save_fm DFF_W1962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3500A));
DFF_save_fm DFF_W1963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3501A));
DFF_save_fm DFF_W1964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3502A));
DFF_save_fm DFF_W1965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3510A));
DFF_save_fm DFF_W1966(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3511A));
DFF_save_fm DFF_W1967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3512A));
DFF_save_fm DFF_W1968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3520A));
DFF_save_fm DFF_W1969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3521A));
DFF_save_fm DFF_W1970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3522A));
DFF_save_fm DFF_W1971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3500B));
DFF_save_fm DFF_W1972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3501B));
DFF_save_fm DFF_W1973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3502B));
DFF_save_fm DFF_W1974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3510B));
DFF_save_fm DFF_W1975(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3511B));
DFF_save_fm DFF_W1976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3512B));
DFF_save_fm DFF_W1977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3520B));
DFF_save_fm DFF_W1978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3521B));
DFF_save_fm DFF_W1979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3522B));
DFF_save_fm DFF_W1980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3500C));
DFF_save_fm DFF_W1981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3501C));
DFF_save_fm DFF_W1982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3502C));
DFF_save_fm DFF_W1983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3510C));
DFF_save_fm DFF_W1984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3511C));
DFF_save_fm DFF_W1985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3512C));
DFF_save_fm DFF_W1986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3520C));
DFF_save_fm DFF_W1987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3521C));
DFF_save_fm DFF_W1988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3522C));
DFF_save_fm DFF_W1989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3500D));
DFF_save_fm DFF_W1990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3501D));
DFF_save_fm DFF_W1991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3502D));
DFF_save_fm DFF_W1992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3510D));
DFF_save_fm DFF_W1993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3511D));
DFF_save_fm DFF_W1994(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3512D));
DFF_save_fm DFF_W1995(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3520D));
DFF_save_fm DFF_W1996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3521D));
DFF_save_fm DFF_W1997(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3522D));
DFF_save_fm DFF_W1998(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3500E));
DFF_save_fm DFF_W1999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3501E));
DFF_save_fm DFF_W2000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3502E));
DFF_save_fm DFF_W2001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3510E));
DFF_save_fm DFF_W2002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3511E));
DFF_save_fm DFF_W2003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3512E));
DFF_save_fm DFF_W2004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3520E));
DFF_save_fm DFF_W2005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3521E));
DFF_save_fm DFF_W2006(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3522E));
DFF_save_fm DFF_W2007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3500F));
DFF_save_fm DFF_W2008(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3501F));
DFF_save_fm DFF_W2009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3502F));
DFF_save_fm DFF_W2010(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3510F));
DFF_save_fm DFF_W2011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3511F));
DFF_save_fm DFF_W2012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3512F));
DFF_save_fm DFF_W2013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3520F));
DFF_save_fm DFF_W2014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3521F));
DFF_save_fm DFF_W2015(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3522F));
DFF_save_fm DFF_W2016(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36000));
DFF_save_fm DFF_W2017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36010));
DFF_save_fm DFF_W2018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36020));
DFF_save_fm DFF_W2019(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36100));
DFF_save_fm DFF_W2020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36110));
DFF_save_fm DFF_W2021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36120));
DFF_save_fm DFF_W2022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36200));
DFF_save_fm DFF_W2023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36210));
DFF_save_fm DFF_W2024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36220));
DFF_save_fm DFF_W2025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36001));
DFF_save_fm DFF_W2026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36011));
DFF_save_fm DFF_W2027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36021));
DFF_save_fm DFF_W2028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36101));
DFF_save_fm DFF_W2029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36111));
DFF_save_fm DFF_W2030(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36121));
DFF_save_fm DFF_W2031(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36201));
DFF_save_fm DFF_W2032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36211));
DFF_save_fm DFF_W2033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36221));
DFF_save_fm DFF_W2034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36002));
DFF_save_fm DFF_W2035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36012));
DFF_save_fm DFF_W2036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36022));
DFF_save_fm DFF_W2037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36102));
DFF_save_fm DFF_W2038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36112));
DFF_save_fm DFF_W2039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36122));
DFF_save_fm DFF_W2040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36202));
DFF_save_fm DFF_W2041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36212));
DFF_save_fm DFF_W2042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36222));
DFF_save_fm DFF_W2043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36003));
DFF_save_fm DFF_W2044(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36013));
DFF_save_fm DFF_W2045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36023));
DFF_save_fm DFF_W2046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36103));
DFF_save_fm DFF_W2047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36113));
DFF_save_fm DFF_W2048(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36123));
DFF_save_fm DFF_W2049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36203));
DFF_save_fm DFF_W2050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36213));
DFF_save_fm DFF_W2051(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36223));
DFF_save_fm DFF_W2052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36004));
DFF_save_fm DFF_W2053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36014));
DFF_save_fm DFF_W2054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36024));
DFF_save_fm DFF_W2055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36104));
DFF_save_fm DFF_W2056(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36114));
DFF_save_fm DFF_W2057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36124));
DFF_save_fm DFF_W2058(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36204));
DFF_save_fm DFF_W2059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36214));
DFF_save_fm DFF_W2060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36224));
DFF_save_fm DFF_W2061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36005));
DFF_save_fm DFF_W2062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36015));
DFF_save_fm DFF_W2063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36025));
DFF_save_fm DFF_W2064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36105));
DFF_save_fm DFF_W2065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36115));
DFF_save_fm DFF_W2066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36125));
DFF_save_fm DFF_W2067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36205));
DFF_save_fm DFF_W2068(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36215));
DFF_save_fm DFF_W2069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36225));
DFF_save_fm DFF_W2070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36006));
DFF_save_fm DFF_W2071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36016));
DFF_save_fm DFF_W2072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36026));
DFF_save_fm DFF_W2073(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36106));
DFF_save_fm DFF_W2074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36116));
DFF_save_fm DFF_W2075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36126));
DFF_save_fm DFF_W2076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36206));
DFF_save_fm DFF_W2077(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36216));
DFF_save_fm DFF_W2078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36226));
DFF_save_fm DFF_W2079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36007));
DFF_save_fm DFF_W2080(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36017));
DFF_save_fm DFF_W2081(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36027));
DFF_save_fm DFF_W2082(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36107));
DFF_save_fm DFF_W2083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36117));
DFF_save_fm DFF_W2084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36127));
DFF_save_fm DFF_W2085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36207));
DFF_save_fm DFF_W2086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36217));
DFF_save_fm DFF_W2087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36227));
DFF_save_fm DFF_W2088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36008));
DFF_save_fm DFF_W2089(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36018));
DFF_save_fm DFF_W2090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36028));
DFF_save_fm DFF_W2091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36108));
DFF_save_fm DFF_W2092(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36118));
DFF_save_fm DFF_W2093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36128));
DFF_save_fm DFF_W2094(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36208));
DFF_save_fm DFF_W2095(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36218));
DFF_save_fm DFF_W2096(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36228));
DFF_save_fm DFF_W2097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36009));
DFF_save_fm DFF_W2098(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36019));
DFF_save_fm DFF_W2099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36029));
DFF_save_fm DFF_W2100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36109));
DFF_save_fm DFF_W2101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36119));
DFF_save_fm DFF_W2102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36129));
DFF_save_fm DFF_W2103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36209));
DFF_save_fm DFF_W2104(.clk(clk),.rstn(rstn),.reset_value(1),.q(W36219));
DFF_save_fm DFF_W2105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W36229));
DFF_save_fm DFF_W2106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3600A));
DFF_save_fm DFF_W2107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3601A));
DFF_save_fm DFF_W2108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3602A));
DFF_save_fm DFF_W2109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3610A));
DFF_save_fm DFF_W2110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3611A));
DFF_save_fm DFF_W2111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3612A));
DFF_save_fm DFF_W2112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3620A));
DFF_save_fm DFF_W2113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3621A));
DFF_save_fm DFF_W2114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3622A));
DFF_save_fm DFF_W2115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3600B));
DFF_save_fm DFF_W2116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3601B));
DFF_save_fm DFF_W2117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3602B));
DFF_save_fm DFF_W2118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3610B));
DFF_save_fm DFF_W2119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3611B));
DFF_save_fm DFF_W2120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3612B));
DFF_save_fm DFF_W2121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3620B));
DFF_save_fm DFF_W2122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3621B));
DFF_save_fm DFF_W2123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3622B));
DFF_save_fm DFF_W2124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3600C));
DFF_save_fm DFF_W2125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3601C));
DFF_save_fm DFF_W2126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3602C));
DFF_save_fm DFF_W2127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3610C));
DFF_save_fm DFF_W2128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3611C));
DFF_save_fm DFF_W2129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3612C));
DFF_save_fm DFF_W2130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3620C));
DFF_save_fm DFF_W2131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3621C));
DFF_save_fm DFF_W2132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3622C));
DFF_save_fm DFF_W2133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3600D));
DFF_save_fm DFF_W2134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3601D));
DFF_save_fm DFF_W2135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3602D));
DFF_save_fm DFF_W2136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3610D));
DFF_save_fm DFF_W2137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3611D));
DFF_save_fm DFF_W2138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3612D));
DFF_save_fm DFF_W2139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3620D));
DFF_save_fm DFF_W2140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3621D));
DFF_save_fm DFF_W2141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3622D));
DFF_save_fm DFF_W2142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3600E));
DFF_save_fm DFF_W2143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3601E));
DFF_save_fm DFF_W2144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3602E));
DFF_save_fm DFF_W2145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3610E));
DFF_save_fm DFF_W2146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3611E));
DFF_save_fm DFF_W2147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3612E));
DFF_save_fm DFF_W2148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3620E));
DFF_save_fm DFF_W2149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3621E));
DFF_save_fm DFF_W2150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3622E));
DFF_save_fm DFF_W2151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3600F));
DFF_save_fm DFF_W2152(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3601F));
DFF_save_fm DFF_W2153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3602F));
DFF_save_fm DFF_W2154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3610F));
DFF_save_fm DFF_W2155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3611F));
DFF_save_fm DFF_W2156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3612F));
DFF_save_fm DFF_W2157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3620F));
DFF_save_fm DFF_W2158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3621F));
DFF_save_fm DFF_W2159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3622F));
DFF_save_fm DFF_W2160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37000));
DFF_save_fm DFF_W2161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37010));
DFF_save_fm DFF_W2162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37020));
DFF_save_fm DFF_W2163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37100));
DFF_save_fm DFF_W2164(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37110));
DFF_save_fm DFF_W2165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37120));
DFF_save_fm DFF_W2166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37200));
DFF_save_fm DFF_W2167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37210));
DFF_save_fm DFF_W2168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37220));
DFF_save_fm DFF_W2169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37001));
DFF_save_fm DFF_W2170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37011));
DFF_save_fm DFF_W2171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37021));
DFF_save_fm DFF_W2172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37101));
DFF_save_fm DFF_W2173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37111));
DFF_save_fm DFF_W2174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37121));
DFF_save_fm DFF_W2175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37201));
DFF_save_fm DFF_W2176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37211));
DFF_save_fm DFF_W2177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37221));
DFF_save_fm DFF_W2178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37002));
DFF_save_fm DFF_W2179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37012));
DFF_save_fm DFF_W2180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37022));
DFF_save_fm DFF_W2181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37102));
DFF_save_fm DFF_W2182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37112));
DFF_save_fm DFF_W2183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37122));
DFF_save_fm DFF_W2184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37202));
DFF_save_fm DFF_W2185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37212));
DFF_save_fm DFF_W2186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37222));
DFF_save_fm DFF_W2187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37003));
DFF_save_fm DFF_W2188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37013));
DFF_save_fm DFF_W2189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37023));
DFF_save_fm DFF_W2190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37103));
DFF_save_fm DFF_W2191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37113));
DFF_save_fm DFF_W2192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37123));
DFF_save_fm DFF_W2193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37203));
DFF_save_fm DFF_W2194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37213));
DFF_save_fm DFF_W2195(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37223));
DFF_save_fm DFF_W2196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37004));
DFF_save_fm DFF_W2197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37014));
DFF_save_fm DFF_W2198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37024));
DFF_save_fm DFF_W2199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37104));
DFF_save_fm DFF_W2200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37114));
DFF_save_fm DFF_W2201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37124));
DFF_save_fm DFF_W2202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37204));
DFF_save_fm DFF_W2203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37214));
DFF_save_fm DFF_W2204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37224));
DFF_save_fm DFF_W2205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37005));
DFF_save_fm DFF_W2206(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37015));
DFF_save_fm DFF_W2207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37025));
DFF_save_fm DFF_W2208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37105));
DFF_save_fm DFF_W2209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37115));
DFF_save_fm DFF_W2210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37125));
DFF_save_fm DFF_W2211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37205));
DFF_save_fm DFF_W2212(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37215));
DFF_save_fm DFF_W2213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37225));
DFF_save_fm DFF_W2214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37006));
DFF_save_fm DFF_W2215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37016));
DFF_save_fm DFF_W2216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37026));
DFF_save_fm DFF_W2217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37106));
DFF_save_fm DFF_W2218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37116));
DFF_save_fm DFF_W2219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37126));
DFF_save_fm DFF_W2220(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37206));
DFF_save_fm DFF_W2221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37216));
DFF_save_fm DFF_W2222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37226));
DFF_save_fm DFF_W2223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37007));
DFF_save_fm DFF_W2224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37017));
DFF_save_fm DFF_W2225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37027));
DFF_save_fm DFF_W2226(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37107));
DFF_save_fm DFF_W2227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37117));
DFF_save_fm DFF_W2228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37127));
DFF_save_fm DFF_W2229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37207));
DFF_save_fm DFF_W2230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37217));
DFF_save_fm DFF_W2231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37227));
DFF_save_fm DFF_W2232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37008));
DFF_save_fm DFF_W2233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37018));
DFF_save_fm DFF_W2234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37028));
DFF_save_fm DFF_W2235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37108));
DFF_save_fm DFF_W2236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37118));
DFF_save_fm DFF_W2237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37128));
DFF_save_fm DFF_W2238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37208));
DFF_save_fm DFF_W2239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37218));
DFF_save_fm DFF_W2240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37228));
DFF_save_fm DFF_W2241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37009));
DFF_save_fm DFF_W2242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37019));
DFF_save_fm DFF_W2243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37029));
DFF_save_fm DFF_W2244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37109));
DFF_save_fm DFF_W2245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37119));
DFF_save_fm DFF_W2246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37129));
DFF_save_fm DFF_W2247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37209));
DFF_save_fm DFF_W2248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W37219));
DFF_save_fm DFF_W2249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W37229));
DFF_save_fm DFF_W2250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3700A));
DFF_save_fm DFF_W2251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3701A));
DFF_save_fm DFF_W2252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3702A));
DFF_save_fm DFF_W2253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3710A));
DFF_save_fm DFF_W2254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3711A));
DFF_save_fm DFF_W2255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3712A));
DFF_save_fm DFF_W2256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3720A));
DFF_save_fm DFF_W2257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3721A));
DFF_save_fm DFF_W2258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3722A));
DFF_save_fm DFF_W2259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3700B));
DFF_save_fm DFF_W2260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3701B));
DFF_save_fm DFF_W2261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3702B));
DFF_save_fm DFF_W2262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3710B));
DFF_save_fm DFF_W2263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3711B));
DFF_save_fm DFF_W2264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3712B));
DFF_save_fm DFF_W2265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3720B));
DFF_save_fm DFF_W2266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3721B));
DFF_save_fm DFF_W2267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3722B));
DFF_save_fm DFF_W2268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3700C));
DFF_save_fm DFF_W2269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3701C));
DFF_save_fm DFF_W2270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3702C));
DFF_save_fm DFF_W2271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3710C));
DFF_save_fm DFF_W2272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3711C));
DFF_save_fm DFF_W2273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3712C));
DFF_save_fm DFF_W2274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3720C));
DFF_save_fm DFF_W2275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3721C));
DFF_save_fm DFF_W2276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3722C));
DFF_save_fm DFF_W2277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3700D));
DFF_save_fm DFF_W2278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3701D));
DFF_save_fm DFF_W2279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3702D));
DFF_save_fm DFF_W2280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3710D));
DFF_save_fm DFF_W2281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3711D));
DFF_save_fm DFF_W2282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3712D));
DFF_save_fm DFF_W2283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3720D));
DFF_save_fm DFF_W2284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3721D));
DFF_save_fm DFF_W2285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3722D));
DFF_save_fm DFF_W2286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3700E));
DFF_save_fm DFF_W2287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3701E));
DFF_save_fm DFF_W2288(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3702E));
DFF_save_fm DFF_W2289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3710E));
DFF_save_fm DFF_W2290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3711E));
DFF_save_fm DFF_W2291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3712E));
DFF_save_fm DFF_W2292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3720E));
DFF_save_fm DFF_W2293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3721E));
DFF_save_fm DFF_W2294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3722E));
DFF_save_fm DFF_W2295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3700F));
DFF_save_fm DFF_W2296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3701F));
DFF_save_fm DFF_W2297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3702F));
DFF_save_fm DFF_W2298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3710F));
DFF_save_fm DFF_W2299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3711F));
DFF_save_fm DFF_W2300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3712F));
DFF_save_fm DFF_W2301(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3720F));
DFF_save_fm DFF_W2302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3721F));
DFF_save_fm DFF_W2303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3722F));
DFF_save_fm DFF_W2304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38000));
DFF_save_fm DFF_W2305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38010));
DFF_save_fm DFF_W2306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38020));
DFF_save_fm DFF_W2307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38100));
DFF_save_fm DFF_W2308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38110));
DFF_save_fm DFF_W2309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38120));
DFF_save_fm DFF_W2310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38200));
DFF_save_fm DFF_W2311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38210));
DFF_save_fm DFF_W2312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38220));
DFF_save_fm DFF_W2313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38001));
DFF_save_fm DFF_W2314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38011));
DFF_save_fm DFF_W2315(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38021));
DFF_save_fm DFF_W2316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38101));
DFF_save_fm DFF_W2317(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38111));
DFF_save_fm DFF_W2318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38121));
DFF_save_fm DFF_W2319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38201));
DFF_save_fm DFF_W2320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38211));
DFF_save_fm DFF_W2321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38221));
DFF_save_fm DFF_W2322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38002));
DFF_save_fm DFF_W2323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38012));
DFF_save_fm DFF_W2324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38022));
DFF_save_fm DFF_W2325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38102));
DFF_save_fm DFF_W2326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38112));
DFF_save_fm DFF_W2327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38122));
DFF_save_fm DFF_W2328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38202));
DFF_save_fm DFF_W2329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38212));
DFF_save_fm DFF_W2330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38222));
DFF_save_fm DFF_W2331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38003));
DFF_save_fm DFF_W2332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38013));
DFF_save_fm DFF_W2333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38023));
DFF_save_fm DFF_W2334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38103));
DFF_save_fm DFF_W2335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38113));
DFF_save_fm DFF_W2336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38123));
DFF_save_fm DFF_W2337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38203));
DFF_save_fm DFF_W2338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38213));
DFF_save_fm DFF_W2339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38223));
DFF_save_fm DFF_W2340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38004));
DFF_save_fm DFF_W2341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38014));
DFF_save_fm DFF_W2342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38024));
DFF_save_fm DFF_W2343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38104));
DFF_save_fm DFF_W2344(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38114));
DFF_save_fm DFF_W2345(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38124));
DFF_save_fm DFF_W2346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38204));
DFF_save_fm DFF_W2347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38214));
DFF_save_fm DFF_W2348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38224));
DFF_save_fm DFF_W2349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38005));
DFF_save_fm DFF_W2350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38015));
DFF_save_fm DFF_W2351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38025));
DFF_save_fm DFF_W2352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38105));
DFF_save_fm DFF_W2353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38115));
DFF_save_fm DFF_W2354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38125));
DFF_save_fm DFF_W2355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38205));
DFF_save_fm DFF_W2356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38215));
DFF_save_fm DFF_W2357(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38225));
DFF_save_fm DFF_W2358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38006));
DFF_save_fm DFF_W2359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38016));
DFF_save_fm DFF_W2360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38026));
DFF_save_fm DFF_W2361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38106));
DFF_save_fm DFF_W2362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38116));
DFF_save_fm DFF_W2363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38126));
DFF_save_fm DFF_W2364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38206));
DFF_save_fm DFF_W2365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38216));
DFF_save_fm DFF_W2366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38226));
DFF_save_fm DFF_W2367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38007));
DFF_save_fm DFF_W2368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38017));
DFF_save_fm DFF_W2369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38027));
DFF_save_fm DFF_W2370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38107));
DFF_save_fm DFF_W2371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38117));
DFF_save_fm DFF_W2372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38127));
DFF_save_fm DFF_W2373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38207));
DFF_save_fm DFF_W2374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38217));
DFF_save_fm DFF_W2375(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38227));
DFF_save_fm DFF_W2376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38008));
DFF_save_fm DFF_W2377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38018));
DFF_save_fm DFF_W2378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38028));
DFF_save_fm DFF_W2379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38108));
DFF_save_fm DFF_W2380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38118));
DFF_save_fm DFF_W2381(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38128));
DFF_save_fm DFF_W2382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38208));
DFF_save_fm DFF_W2383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38218));
DFF_save_fm DFF_W2384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38228));
DFF_save_fm DFF_W2385(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38009));
DFF_save_fm DFF_W2386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38019));
DFF_save_fm DFF_W2387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38029));
DFF_save_fm DFF_W2388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38109));
DFF_save_fm DFF_W2389(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38119));
DFF_save_fm DFF_W2390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38129));
DFF_save_fm DFF_W2391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W38209));
DFF_save_fm DFF_W2392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38219));
DFF_save_fm DFF_W2393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W38229));
DFF_save_fm DFF_W2394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3800A));
DFF_save_fm DFF_W2395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3801A));
DFF_save_fm DFF_W2396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3802A));
DFF_save_fm DFF_W2397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3810A));
DFF_save_fm DFF_W2398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3811A));
DFF_save_fm DFF_W2399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3812A));
DFF_save_fm DFF_W2400(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3820A));
DFF_save_fm DFF_W2401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3821A));
DFF_save_fm DFF_W2402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3822A));
DFF_save_fm DFF_W2403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3800B));
DFF_save_fm DFF_W2404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3801B));
DFF_save_fm DFF_W2405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3802B));
DFF_save_fm DFF_W2406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3810B));
DFF_save_fm DFF_W2407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3811B));
DFF_save_fm DFF_W2408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3812B));
DFF_save_fm DFF_W2409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3820B));
DFF_save_fm DFF_W2410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3821B));
DFF_save_fm DFF_W2411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3822B));
DFF_save_fm DFF_W2412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3800C));
DFF_save_fm DFF_W2413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3801C));
DFF_save_fm DFF_W2414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3802C));
DFF_save_fm DFF_W2415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3810C));
DFF_save_fm DFF_W2416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3811C));
DFF_save_fm DFF_W2417(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3812C));
DFF_save_fm DFF_W2418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3820C));
DFF_save_fm DFF_W2419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3821C));
DFF_save_fm DFF_W2420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3822C));
DFF_save_fm DFF_W2421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3800D));
DFF_save_fm DFF_W2422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3801D));
DFF_save_fm DFF_W2423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3802D));
DFF_save_fm DFF_W2424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3810D));
DFF_save_fm DFF_W2425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3811D));
DFF_save_fm DFF_W2426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3812D));
DFF_save_fm DFF_W2427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3820D));
DFF_save_fm DFF_W2428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3821D));
DFF_save_fm DFF_W2429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3822D));
DFF_save_fm DFF_W2430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3800E));
DFF_save_fm DFF_W2431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3801E));
DFF_save_fm DFF_W2432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3802E));
DFF_save_fm DFF_W2433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3810E));
DFF_save_fm DFF_W2434(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3811E));
DFF_save_fm DFF_W2435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3812E));
DFF_save_fm DFF_W2436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3820E));
DFF_save_fm DFF_W2437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3821E));
DFF_save_fm DFF_W2438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3822E));
DFF_save_fm DFF_W2439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3800F));
DFF_save_fm DFF_W2440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3801F));
DFF_save_fm DFF_W2441(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3802F));
DFF_save_fm DFF_W2442(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3810F));
DFF_save_fm DFF_W2443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3811F));
DFF_save_fm DFF_W2444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3812F));
DFF_save_fm DFF_W2445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3820F));
DFF_save_fm DFF_W2446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3821F));
DFF_save_fm DFF_W2447(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3822F));
DFF_save_fm DFF_W2448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39000));
DFF_save_fm DFF_W2449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39010));
DFF_save_fm DFF_W2450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39020));
DFF_save_fm DFF_W2451(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39100));
DFF_save_fm DFF_W2452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39110));
DFF_save_fm DFF_W2453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39120));
DFF_save_fm DFF_W2454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39200));
DFF_save_fm DFF_W2455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39210));
DFF_save_fm DFF_W2456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39220));
DFF_save_fm DFF_W2457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39001));
DFF_save_fm DFF_W2458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39011));
DFF_save_fm DFF_W2459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39021));
DFF_save_fm DFF_W2460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39101));
DFF_save_fm DFF_W2461(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39111));
DFF_save_fm DFF_W2462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39121));
DFF_save_fm DFF_W2463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39201));
DFF_save_fm DFF_W2464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39211));
DFF_save_fm DFF_W2465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39221));
DFF_save_fm DFF_W2466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39002));
DFF_save_fm DFF_W2467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39012));
DFF_save_fm DFF_W2468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39022));
DFF_save_fm DFF_W2469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39102));
DFF_save_fm DFF_W2470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39112));
DFF_save_fm DFF_W2471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39122));
DFF_save_fm DFF_W2472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39202));
DFF_save_fm DFF_W2473(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39212));
DFF_save_fm DFF_W2474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39222));
DFF_save_fm DFF_W2475(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39003));
DFF_save_fm DFF_W2476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39013));
DFF_save_fm DFF_W2477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39023));
DFF_save_fm DFF_W2478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39103));
DFF_save_fm DFF_W2479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39113));
DFF_save_fm DFF_W2480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39123));
DFF_save_fm DFF_W2481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39203));
DFF_save_fm DFF_W2482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39213));
DFF_save_fm DFF_W2483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39223));
DFF_save_fm DFF_W2484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39004));
DFF_save_fm DFF_W2485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39014));
DFF_save_fm DFF_W2486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39024));
DFF_save_fm DFF_W2487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39104));
DFF_save_fm DFF_W2488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39114));
DFF_save_fm DFF_W2489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39124));
DFF_save_fm DFF_W2490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39204));
DFF_save_fm DFF_W2491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39214));
DFF_save_fm DFF_W2492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39224));
DFF_save_fm DFF_W2493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39005));
DFF_save_fm DFF_W2494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39015));
DFF_save_fm DFF_W2495(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39025));
DFF_save_fm DFF_W2496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39105));
DFF_save_fm DFF_W2497(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39115));
DFF_save_fm DFF_W2498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39125));
DFF_save_fm DFF_W2499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39205));
DFF_save_fm DFF_W2500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39215));
DFF_save_fm DFF_W2501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39225));
DFF_save_fm DFF_W2502(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39006));
DFF_save_fm DFF_W2503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39016));
DFF_save_fm DFF_W2504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39026));
DFF_save_fm DFF_W2505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39106));
DFF_save_fm DFF_W2506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39116));
DFF_save_fm DFF_W2507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39126));
DFF_save_fm DFF_W2508(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39206));
DFF_save_fm DFF_W2509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39216));
DFF_save_fm DFF_W2510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39226));
DFF_save_fm DFF_W2511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39007));
DFF_save_fm DFF_W2512(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39017));
DFF_save_fm DFF_W2513(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39027));
DFF_save_fm DFF_W2514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39107));
DFF_save_fm DFF_W2515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39117));
DFF_save_fm DFF_W2516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39127));
DFF_save_fm DFF_W2517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39207));
DFF_save_fm DFF_W2518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39217));
DFF_save_fm DFF_W2519(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39227));
DFF_save_fm DFF_W2520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39008));
DFF_save_fm DFF_W2521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39018));
DFF_save_fm DFF_W2522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39028));
DFF_save_fm DFF_W2523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39108));
DFF_save_fm DFF_W2524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39118));
DFF_save_fm DFF_W2525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39128));
DFF_save_fm DFF_W2526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39208));
DFF_save_fm DFF_W2527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39218));
DFF_save_fm DFF_W2528(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39228));
DFF_save_fm DFF_W2529(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39009));
DFF_save_fm DFF_W2530(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39019));
DFF_save_fm DFF_W2531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39029));
DFF_save_fm DFF_W2532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39109));
DFF_save_fm DFF_W2533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W39119));
DFF_save_fm DFF_W2534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39129));
DFF_save_fm DFF_W2535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39209));
DFF_save_fm DFF_W2536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39219));
DFF_save_fm DFF_W2537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W39229));
DFF_save_fm DFF_W2538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3900A));
DFF_save_fm DFF_W2539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3901A));
DFF_save_fm DFF_W2540(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3902A));
DFF_save_fm DFF_W2541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3910A));
DFF_save_fm DFF_W2542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3911A));
DFF_save_fm DFF_W2543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3912A));
DFF_save_fm DFF_W2544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3920A));
DFF_save_fm DFF_W2545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3921A));
DFF_save_fm DFF_W2546(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3922A));
DFF_save_fm DFF_W2547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3900B));
DFF_save_fm DFF_W2548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3901B));
DFF_save_fm DFF_W2549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3902B));
DFF_save_fm DFF_W2550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3910B));
DFF_save_fm DFF_W2551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3911B));
DFF_save_fm DFF_W2552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3912B));
DFF_save_fm DFF_W2553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3920B));
DFF_save_fm DFF_W2554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3921B));
DFF_save_fm DFF_W2555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3922B));
DFF_save_fm DFF_W2556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3900C));
DFF_save_fm DFF_W2557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3901C));
DFF_save_fm DFF_W2558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3902C));
DFF_save_fm DFF_W2559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3910C));
DFF_save_fm DFF_W2560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3911C));
DFF_save_fm DFF_W2561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3912C));
DFF_save_fm DFF_W2562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3920C));
DFF_save_fm DFF_W2563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3921C));
DFF_save_fm DFF_W2564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3922C));
DFF_save_fm DFF_W2565(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3900D));
DFF_save_fm DFF_W2566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3901D));
DFF_save_fm DFF_W2567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3902D));
DFF_save_fm DFF_W2568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3910D));
DFF_save_fm DFF_W2569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3911D));
DFF_save_fm DFF_W2570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3912D));
DFF_save_fm DFF_W2571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3920D));
DFF_save_fm DFF_W2572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3921D));
DFF_save_fm DFF_W2573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3922D));
DFF_save_fm DFF_W2574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3900E));
DFF_save_fm DFF_W2575(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3901E));
DFF_save_fm DFF_W2576(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3902E));
DFF_save_fm DFF_W2577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3910E));
DFF_save_fm DFF_W2578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3911E));
DFF_save_fm DFF_W2579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3912E));
DFF_save_fm DFF_W2580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3920E));
DFF_save_fm DFF_W2581(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3921E));
DFF_save_fm DFF_W2582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3922E));
DFF_save_fm DFF_W2583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3900F));
DFF_save_fm DFF_W2584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3901F));
DFF_save_fm DFF_W2585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3902F));
DFF_save_fm DFF_W2586(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3910F));
DFF_save_fm DFF_W2587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3911F));
DFF_save_fm DFF_W2588(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3912F));
DFF_save_fm DFF_W2589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3920F));
DFF_save_fm DFF_W2590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3921F));
DFF_save_fm DFF_W2591(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3922F));
DFF_save_fm DFF_W2592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A000));
DFF_save_fm DFF_W2593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A010));
DFF_save_fm DFF_W2594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A020));
DFF_save_fm DFF_W2595(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A100));
DFF_save_fm DFF_W2596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A110));
DFF_save_fm DFF_W2597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A120));
DFF_save_fm DFF_W2598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A200));
DFF_save_fm DFF_W2599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A210));
DFF_save_fm DFF_W2600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A220));
DFF_save_fm DFF_W2601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A001));
DFF_save_fm DFF_W2602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A011));
DFF_save_fm DFF_W2603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A021));
DFF_save_fm DFF_W2604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A101));
DFF_save_fm DFF_W2605(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A111));
DFF_save_fm DFF_W2606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A121));
DFF_save_fm DFF_W2607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A201));
DFF_save_fm DFF_W2608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A211));
DFF_save_fm DFF_W2609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A221));
DFF_save_fm DFF_W2610(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A002));
DFF_save_fm DFF_W2611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A012));
DFF_save_fm DFF_W2612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A022));
DFF_save_fm DFF_W2613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A102));
DFF_save_fm DFF_W2614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A112));
DFF_save_fm DFF_W2615(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A122));
DFF_save_fm DFF_W2616(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A202));
DFF_save_fm DFF_W2617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A212));
DFF_save_fm DFF_W2618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A222));
DFF_save_fm DFF_W2619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A003));
DFF_save_fm DFF_W2620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A013));
DFF_save_fm DFF_W2621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A023));
DFF_save_fm DFF_W2622(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A103));
DFF_save_fm DFF_W2623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A113));
DFF_save_fm DFF_W2624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A123));
DFF_save_fm DFF_W2625(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A203));
DFF_save_fm DFF_W2626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A213));
DFF_save_fm DFF_W2627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A223));
DFF_save_fm DFF_W2628(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A004));
DFF_save_fm DFF_W2629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A014));
DFF_save_fm DFF_W2630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A024));
DFF_save_fm DFF_W2631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A104));
DFF_save_fm DFF_W2632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A114));
DFF_save_fm DFF_W2633(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A124));
DFF_save_fm DFF_W2634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A204));
DFF_save_fm DFF_W2635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A214));
DFF_save_fm DFF_W2636(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A224));
DFF_save_fm DFF_W2637(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A005));
DFF_save_fm DFF_W2638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A015));
DFF_save_fm DFF_W2639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A025));
DFF_save_fm DFF_W2640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A105));
DFF_save_fm DFF_W2641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A115));
DFF_save_fm DFF_W2642(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A125));
DFF_save_fm DFF_W2643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A205));
DFF_save_fm DFF_W2644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A215));
DFF_save_fm DFF_W2645(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A225));
DFF_save_fm DFF_W2646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A006));
DFF_save_fm DFF_W2647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A016));
DFF_save_fm DFF_W2648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A026));
DFF_save_fm DFF_W2649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A106));
DFF_save_fm DFF_W2650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A116));
DFF_save_fm DFF_W2651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A126));
DFF_save_fm DFF_W2652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A206));
DFF_save_fm DFF_W2653(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A216));
DFF_save_fm DFF_W2654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A226));
DFF_save_fm DFF_W2655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A007));
DFF_save_fm DFF_W2656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A017));
DFF_save_fm DFF_W2657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A027));
DFF_save_fm DFF_W2658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A107));
DFF_save_fm DFF_W2659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A117));
DFF_save_fm DFF_W2660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A127));
DFF_save_fm DFF_W2661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A207));
DFF_save_fm DFF_W2662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A217));
DFF_save_fm DFF_W2663(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A227));
DFF_save_fm DFF_W2664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A008));
DFF_save_fm DFF_W2665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A018));
DFF_save_fm DFF_W2666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A028));
DFF_save_fm DFF_W2667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A108));
DFF_save_fm DFF_W2668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A118));
DFF_save_fm DFF_W2669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A128));
DFF_save_fm DFF_W2670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A208));
DFF_save_fm DFF_W2671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A218));
DFF_save_fm DFF_W2672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A228));
DFF_save_fm DFF_W2673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A009));
DFF_save_fm DFF_W2674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A019));
DFF_save_fm DFF_W2675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A029));
DFF_save_fm DFF_W2676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A109));
DFF_save_fm DFF_W2677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A119));
DFF_save_fm DFF_W2678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A129));
DFF_save_fm DFF_W2679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A209));
DFF_save_fm DFF_W2680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A219));
DFF_save_fm DFF_W2681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A229));
DFF_save_fm DFF_W2682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A00A));
DFF_save_fm DFF_W2683(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A01A));
DFF_save_fm DFF_W2684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A02A));
DFF_save_fm DFF_W2685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A10A));
DFF_save_fm DFF_W2686(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A11A));
DFF_save_fm DFF_W2687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A12A));
DFF_save_fm DFF_W2688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A20A));
DFF_save_fm DFF_W2689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A21A));
DFF_save_fm DFF_W2690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A22A));
DFF_save_fm DFF_W2691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A00B));
DFF_save_fm DFF_W2692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A01B));
DFF_save_fm DFF_W2693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A02B));
DFF_save_fm DFF_W2694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A10B));
DFF_save_fm DFF_W2695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A11B));
DFF_save_fm DFF_W2696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A12B));
DFF_save_fm DFF_W2697(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A20B));
DFF_save_fm DFF_W2698(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A21B));
DFF_save_fm DFF_W2699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A22B));
DFF_save_fm DFF_W2700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A00C));
DFF_save_fm DFF_W2701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A01C));
DFF_save_fm DFF_W2702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A02C));
DFF_save_fm DFF_W2703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A10C));
DFF_save_fm DFF_W2704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A11C));
DFF_save_fm DFF_W2705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A12C));
DFF_save_fm DFF_W2706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A20C));
DFF_save_fm DFF_W2707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A21C));
DFF_save_fm DFF_W2708(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A22C));
DFF_save_fm DFF_W2709(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A00D));
DFF_save_fm DFF_W2710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A01D));
DFF_save_fm DFF_W2711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A02D));
DFF_save_fm DFF_W2712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A10D));
DFF_save_fm DFF_W2713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A11D));
DFF_save_fm DFF_W2714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A12D));
DFF_save_fm DFF_W2715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A20D));
DFF_save_fm DFF_W2716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A21D));
DFF_save_fm DFF_W2717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A22D));
DFF_save_fm DFF_W2718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A00E));
DFF_save_fm DFF_W2719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A01E));
DFF_save_fm DFF_W2720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A02E));
DFF_save_fm DFF_W2721(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A10E));
DFF_save_fm DFF_W2722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A11E));
DFF_save_fm DFF_W2723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A12E));
DFF_save_fm DFF_W2724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A20E));
DFF_save_fm DFF_W2725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A21E));
DFF_save_fm DFF_W2726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A22E));
DFF_save_fm DFF_W2727(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A00F));
DFF_save_fm DFF_W2728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A01F));
DFF_save_fm DFF_W2729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A02F));
DFF_save_fm DFF_W2730(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A10F));
DFF_save_fm DFF_W2731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A11F));
DFF_save_fm DFF_W2732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A12F));
DFF_save_fm DFF_W2733(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A20F));
DFF_save_fm DFF_W2734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3A21F));
DFF_save_fm DFF_W2735(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3A22F));
DFF_save_fm DFF_W2736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B000));
DFF_save_fm DFF_W2737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B010));
DFF_save_fm DFF_W2738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B020));
DFF_save_fm DFF_W2739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B100));
DFF_save_fm DFF_W2740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B110));
DFF_save_fm DFF_W2741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B120));
DFF_save_fm DFF_W2742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B200));
DFF_save_fm DFF_W2743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B210));
DFF_save_fm DFF_W2744(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B220));
DFF_save_fm DFF_W2745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B001));
DFF_save_fm DFF_W2746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B011));
DFF_save_fm DFF_W2747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B021));
DFF_save_fm DFF_W2748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B101));
DFF_save_fm DFF_W2749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B111));
DFF_save_fm DFF_W2750(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B121));
DFF_save_fm DFF_W2751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B201));
DFF_save_fm DFF_W2752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B211));
DFF_save_fm DFF_W2753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B221));
DFF_save_fm DFF_W2754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B002));
DFF_save_fm DFF_W2755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B012));
DFF_save_fm DFF_W2756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B022));
DFF_save_fm DFF_W2757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B102));
DFF_save_fm DFF_W2758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B112));
DFF_save_fm DFF_W2759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B122));
DFF_save_fm DFF_W2760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B202));
DFF_save_fm DFF_W2761(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B212));
DFF_save_fm DFF_W2762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B222));
DFF_save_fm DFF_W2763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B003));
DFF_save_fm DFF_W2764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B013));
DFF_save_fm DFF_W2765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B023));
DFF_save_fm DFF_W2766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B103));
DFF_save_fm DFF_W2767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B113));
DFF_save_fm DFF_W2768(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B123));
DFF_save_fm DFF_W2769(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B203));
DFF_save_fm DFF_W2770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B213));
DFF_save_fm DFF_W2771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B223));
DFF_save_fm DFF_W2772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B004));
DFF_save_fm DFF_W2773(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B014));
DFF_save_fm DFF_W2774(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B024));
DFF_save_fm DFF_W2775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B104));
DFF_save_fm DFF_W2776(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B114));
DFF_save_fm DFF_W2777(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B124));
DFF_save_fm DFF_W2778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B204));
DFF_save_fm DFF_W2779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B214));
DFF_save_fm DFF_W2780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B224));
DFF_save_fm DFF_W2781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B005));
DFF_save_fm DFF_W2782(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B015));
DFF_save_fm DFF_W2783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B025));
DFF_save_fm DFF_W2784(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B105));
DFF_save_fm DFF_W2785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B115));
DFF_save_fm DFF_W2786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B125));
DFF_save_fm DFF_W2787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B205));
DFF_save_fm DFF_W2788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B215));
DFF_save_fm DFF_W2789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B225));
DFF_save_fm DFF_W2790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B006));
DFF_save_fm DFF_W2791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B016));
DFF_save_fm DFF_W2792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B026));
DFF_save_fm DFF_W2793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B106));
DFF_save_fm DFF_W2794(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B116));
DFF_save_fm DFF_W2795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B126));
DFF_save_fm DFF_W2796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B206));
DFF_save_fm DFF_W2797(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B216));
DFF_save_fm DFF_W2798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B226));
DFF_save_fm DFF_W2799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B007));
DFF_save_fm DFF_W2800(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B017));
DFF_save_fm DFF_W2801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B027));
DFF_save_fm DFF_W2802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B107));
DFF_save_fm DFF_W2803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B117));
DFF_save_fm DFF_W2804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B127));
DFF_save_fm DFF_W2805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B207));
DFF_save_fm DFF_W2806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B217));
DFF_save_fm DFF_W2807(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B227));
DFF_save_fm DFF_W2808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B008));
DFF_save_fm DFF_W2809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B018));
DFF_save_fm DFF_W2810(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B028));
DFF_save_fm DFF_W2811(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B108));
DFF_save_fm DFF_W2812(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B118));
DFF_save_fm DFF_W2813(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B128));
DFF_save_fm DFF_W2814(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B208));
DFF_save_fm DFF_W2815(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B218));
DFF_save_fm DFF_W2816(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B228));
DFF_save_fm DFF_W2817(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B009));
DFF_save_fm DFF_W2818(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B019));
DFF_save_fm DFF_W2819(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B029));
DFF_save_fm DFF_W2820(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B109));
DFF_save_fm DFF_W2821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B119));
DFF_save_fm DFF_W2822(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B129));
DFF_save_fm DFF_W2823(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B209));
DFF_save_fm DFF_W2824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B219));
DFF_save_fm DFF_W2825(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B229));
DFF_save_fm DFF_W2826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B00A));
DFF_save_fm DFF_W2827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B01A));
DFF_save_fm DFF_W2828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B02A));
DFF_save_fm DFF_W2829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B10A));
DFF_save_fm DFF_W2830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B11A));
DFF_save_fm DFF_W2831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B12A));
DFF_save_fm DFF_W2832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B20A));
DFF_save_fm DFF_W2833(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B21A));
DFF_save_fm DFF_W2834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B22A));
DFF_save_fm DFF_W2835(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B00B));
DFF_save_fm DFF_W2836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B01B));
DFF_save_fm DFF_W2837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B02B));
DFF_save_fm DFF_W2838(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B10B));
DFF_save_fm DFF_W2839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B11B));
DFF_save_fm DFF_W2840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B12B));
DFF_save_fm DFF_W2841(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B20B));
DFF_save_fm DFF_W2842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B21B));
DFF_save_fm DFF_W2843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B22B));
DFF_save_fm DFF_W2844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B00C));
DFF_save_fm DFF_W2845(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B01C));
DFF_save_fm DFF_W2846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B02C));
DFF_save_fm DFF_W2847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B10C));
DFF_save_fm DFF_W2848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B11C));
DFF_save_fm DFF_W2849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B12C));
DFF_save_fm DFF_W2850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B20C));
DFF_save_fm DFF_W2851(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B21C));
DFF_save_fm DFF_W2852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B22C));
DFF_save_fm DFF_W2853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B00D));
DFF_save_fm DFF_W2854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B01D));
DFF_save_fm DFF_W2855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B02D));
DFF_save_fm DFF_W2856(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B10D));
DFF_save_fm DFF_W2857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B11D));
DFF_save_fm DFF_W2858(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B12D));
DFF_save_fm DFF_W2859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B20D));
DFF_save_fm DFF_W2860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B21D));
DFF_save_fm DFF_W2861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B22D));
DFF_save_fm DFF_W2862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B00E));
DFF_save_fm DFF_W2863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B01E));
DFF_save_fm DFF_W2864(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B02E));
DFF_save_fm DFF_W2865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B10E));
DFF_save_fm DFF_W2866(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B11E));
DFF_save_fm DFF_W2867(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B12E));
DFF_save_fm DFF_W2868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B20E));
DFF_save_fm DFF_W2869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B21E));
DFF_save_fm DFF_W2870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B22E));
DFF_save_fm DFF_W2871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B00F));
DFF_save_fm DFF_W2872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B01F));
DFF_save_fm DFF_W2873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B02F));
DFF_save_fm DFF_W2874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B10F));
DFF_save_fm DFF_W2875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B11F));
DFF_save_fm DFF_W2876(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B12F));
DFF_save_fm DFF_W2877(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3B20F));
DFF_save_fm DFF_W2878(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B21F));
DFF_save_fm DFF_W2879(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3B22F));
DFF_save_fm DFF_W2880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C000));
DFF_save_fm DFF_W2881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C010));
DFF_save_fm DFF_W2882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C020));
DFF_save_fm DFF_W2883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C100));
DFF_save_fm DFF_W2884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C110));
DFF_save_fm DFF_W2885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C120));
DFF_save_fm DFF_W2886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C200));
DFF_save_fm DFF_W2887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C210));
DFF_save_fm DFF_W2888(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C220));
DFF_save_fm DFF_W2889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C001));
DFF_save_fm DFF_W2890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C011));
DFF_save_fm DFF_W2891(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C021));
DFF_save_fm DFF_W2892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C101));
DFF_save_fm DFF_W2893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C111));
DFF_save_fm DFF_W2894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C121));
DFF_save_fm DFF_W2895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C201));
DFF_save_fm DFF_W2896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C211));
DFF_save_fm DFF_W2897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C221));
DFF_save_fm DFF_W2898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C002));
DFF_save_fm DFF_W2899(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C012));
DFF_save_fm DFF_W2900(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C022));
DFF_save_fm DFF_W2901(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C102));
DFF_save_fm DFF_W2902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C112));
DFF_save_fm DFF_W2903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C122));
DFF_save_fm DFF_W2904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C202));
DFF_save_fm DFF_W2905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C212));
DFF_save_fm DFF_W2906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C222));
DFF_save_fm DFF_W2907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C003));
DFF_save_fm DFF_W2908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C013));
DFF_save_fm DFF_W2909(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C023));
DFF_save_fm DFF_W2910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C103));
DFF_save_fm DFF_W2911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C113));
DFF_save_fm DFF_W2912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C123));
DFF_save_fm DFF_W2913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C203));
DFF_save_fm DFF_W2914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C213));
DFF_save_fm DFF_W2915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C223));
DFF_save_fm DFF_W2916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C004));
DFF_save_fm DFF_W2917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C014));
DFF_save_fm DFF_W2918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C024));
DFF_save_fm DFF_W2919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C104));
DFF_save_fm DFF_W2920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C114));
DFF_save_fm DFF_W2921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C124));
DFF_save_fm DFF_W2922(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C204));
DFF_save_fm DFF_W2923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C214));
DFF_save_fm DFF_W2924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C224));
DFF_save_fm DFF_W2925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C005));
DFF_save_fm DFF_W2926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C015));
DFF_save_fm DFF_W2927(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C025));
DFF_save_fm DFF_W2928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C105));
DFF_save_fm DFF_W2929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C115));
DFF_save_fm DFF_W2930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C125));
DFF_save_fm DFF_W2931(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C205));
DFF_save_fm DFF_W2932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C215));
DFF_save_fm DFF_W2933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C225));
DFF_save_fm DFF_W2934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C006));
DFF_save_fm DFF_W2935(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C016));
DFF_save_fm DFF_W2936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C026));
DFF_save_fm DFF_W2937(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C106));
DFF_save_fm DFF_W2938(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C116));
DFF_save_fm DFF_W2939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C126));
DFF_save_fm DFF_W2940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C206));
DFF_save_fm DFF_W2941(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C216));
DFF_save_fm DFF_W2942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C226));
DFF_save_fm DFF_W2943(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C007));
DFF_save_fm DFF_W2944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C017));
DFF_save_fm DFF_W2945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C027));
DFF_save_fm DFF_W2946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C107));
DFF_save_fm DFF_W2947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C117));
DFF_save_fm DFF_W2948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C127));
DFF_save_fm DFF_W2949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C207));
DFF_save_fm DFF_W2950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C217));
DFF_save_fm DFF_W2951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C227));
DFF_save_fm DFF_W2952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C008));
DFF_save_fm DFF_W2953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C018));
DFF_save_fm DFF_W2954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C028));
DFF_save_fm DFF_W2955(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C108));
DFF_save_fm DFF_W2956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C118));
DFF_save_fm DFF_W2957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C128));
DFF_save_fm DFF_W2958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C208));
DFF_save_fm DFF_W2959(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C218));
DFF_save_fm DFF_W2960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C228));
DFF_save_fm DFF_W2961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C009));
DFF_save_fm DFF_W2962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C019));
DFF_save_fm DFF_W2963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C029));
DFF_save_fm DFF_W2964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C109));
DFF_save_fm DFF_W2965(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C119));
DFF_save_fm DFF_W2966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C129));
DFF_save_fm DFF_W2967(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C209));
DFF_save_fm DFF_W2968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C219));
DFF_save_fm DFF_W2969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C229));
DFF_save_fm DFF_W2970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C00A));
DFF_save_fm DFF_W2971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C01A));
DFF_save_fm DFF_W2972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C02A));
DFF_save_fm DFF_W2973(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C10A));
DFF_save_fm DFF_W2974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C11A));
DFF_save_fm DFF_W2975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C12A));
DFF_save_fm DFF_W2976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C20A));
DFF_save_fm DFF_W2977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C21A));
DFF_save_fm DFF_W2978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C22A));
DFF_save_fm DFF_W2979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C00B));
DFF_save_fm DFF_W2980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C01B));
DFF_save_fm DFF_W2981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C02B));
DFF_save_fm DFF_W2982(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C10B));
DFF_save_fm DFF_W2983(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C11B));
DFF_save_fm DFF_W2984(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C12B));
DFF_save_fm DFF_W2985(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C20B));
DFF_save_fm DFF_W2986(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C21B));
DFF_save_fm DFF_W2987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C22B));
DFF_save_fm DFF_W2988(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C00C));
DFF_save_fm DFF_W2989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C01C));
DFF_save_fm DFF_W2990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C02C));
DFF_save_fm DFF_W2991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C10C));
DFF_save_fm DFF_W2992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C11C));
DFF_save_fm DFF_W2993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C12C));
DFF_save_fm DFF_W2994(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C20C));
DFF_save_fm DFF_W2995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C21C));
DFF_save_fm DFF_W2996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C22C));
DFF_save_fm DFF_W2997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C00D));
DFF_save_fm DFF_W2998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C01D));
DFF_save_fm DFF_W2999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C02D));
DFF_save_fm DFF_W3000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C10D));
DFF_save_fm DFF_W3001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C11D));
DFF_save_fm DFF_W3002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C12D));
DFF_save_fm DFF_W3003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C20D));
DFF_save_fm DFF_W3004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C21D));
DFF_save_fm DFF_W3005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C22D));
DFF_save_fm DFF_W3006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C00E));
DFF_save_fm DFF_W3007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C01E));
DFF_save_fm DFF_W3008(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C02E));
DFF_save_fm DFF_W3009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C10E));
DFF_save_fm DFF_W3010(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C11E));
DFF_save_fm DFF_W3011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C12E));
DFF_save_fm DFF_W3012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C20E));
DFF_save_fm DFF_W3013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C21E));
DFF_save_fm DFF_W3014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C22E));
DFF_save_fm DFF_W3015(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C00F));
DFF_save_fm DFF_W3016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C01F));
DFF_save_fm DFF_W3017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C02F));
DFF_save_fm DFF_W3018(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C10F));
DFF_save_fm DFF_W3019(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C11F));
DFF_save_fm DFF_W3020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3C12F));
DFF_save_fm DFF_W3021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C20F));
DFF_save_fm DFF_W3022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C21F));
DFF_save_fm DFF_W3023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3C22F));
DFF_save_fm DFF_W3024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D000));
DFF_save_fm DFF_W3025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D010));
DFF_save_fm DFF_W3026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D020));
DFF_save_fm DFF_W3027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D100));
DFF_save_fm DFF_W3028(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D110));
DFF_save_fm DFF_W3029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D120));
DFF_save_fm DFF_W3030(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D200));
DFF_save_fm DFF_W3031(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D210));
DFF_save_fm DFF_W3032(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D220));
DFF_save_fm DFF_W3033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D001));
DFF_save_fm DFF_W3034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D011));
DFF_save_fm DFF_W3035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D021));
DFF_save_fm DFF_W3036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D101));
DFF_save_fm DFF_W3037(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D111));
DFF_save_fm DFF_W3038(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D121));
DFF_save_fm DFF_W3039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D201));
DFF_save_fm DFF_W3040(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D211));
DFF_save_fm DFF_W3041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D221));
DFF_save_fm DFF_W3042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D002));
DFF_save_fm DFF_W3043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D012));
DFF_save_fm DFF_W3044(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D022));
DFF_save_fm DFF_W3045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D102));
DFF_save_fm DFF_W3046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D112));
DFF_save_fm DFF_W3047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D122));
DFF_save_fm DFF_W3048(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D202));
DFF_save_fm DFF_W3049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D212));
DFF_save_fm DFF_W3050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D222));
DFF_save_fm DFF_W3051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D003));
DFF_save_fm DFF_W3052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D013));
DFF_save_fm DFF_W3053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D023));
DFF_save_fm DFF_W3054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D103));
DFF_save_fm DFF_W3055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D113));
DFF_save_fm DFF_W3056(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D123));
DFF_save_fm DFF_W3057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D203));
DFF_save_fm DFF_W3058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D213));
DFF_save_fm DFF_W3059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D223));
DFF_save_fm DFF_W3060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D004));
DFF_save_fm DFF_W3061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D014));
DFF_save_fm DFF_W3062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D024));
DFF_save_fm DFF_W3063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D104));
DFF_save_fm DFF_W3064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D114));
DFF_save_fm DFF_W3065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D124));
DFF_save_fm DFF_W3066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D204));
DFF_save_fm DFF_W3067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D214));
DFF_save_fm DFF_W3068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D224));
DFF_save_fm DFF_W3069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D005));
DFF_save_fm DFF_W3070(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D015));
DFF_save_fm DFF_W3071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D025));
DFF_save_fm DFF_W3072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D105));
DFF_save_fm DFF_W3073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D115));
DFF_save_fm DFF_W3074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D125));
DFF_save_fm DFF_W3075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D205));
DFF_save_fm DFF_W3076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D215));
DFF_save_fm DFF_W3077(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D225));
DFF_save_fm DFF_W3078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D006));
DFF_save_fm DFF_W3079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D016));
DFF_save_fm DFF_W3080(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D026));
DFF_save_fm DFF_W3081(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D106));
DFF_save_fm DFF_W3082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D116));
DFF_save_fm DFF_W3083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D126));
DFF_save_fm DFF_W3084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D206));
DFF_save_fm DFF_W3085(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D216));
DFF_save_fm DFF_W3086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D226));
DFF_save_fm DFF_W3087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D007));
DFF_save_fm DFF_W3088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D017));
DFF_save_fm DFF_W3089(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D027));
DFF_save_fm DFF_W3090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D107));
DFF_save_fm DFF_W3091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D117));
DFF_save_fm DFF_W3092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D127));
DFF_save_fm DFF_W3093(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D207));
DFF_save_fm DFF_W3094(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D217));
DFF_save_fm DFF_W3095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D227));
DFF_save_fm DFF_W3096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D008));
DFF_save_fm DFF_W3097(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D018));
DFF_save_fm DFF_W3098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D028));
DFF_save_fm DFF_W3099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D108));
DFF_save_fm DFF_W3100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D118));
DFF_save_fm DFF_W3101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D128));
DFF_save_fm DFF_W3102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D208));
DFF_save_fm DFF_W3103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D218));
DFF_save_fm DFF_W3104(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D228));
DFF_save_fm DFF_W3105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D009));
DFF_save_fm DFF_W3106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D019));
DFF_save_fm DFF_W3107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D029));
DFF_save_fm DFF_W3108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D109));
DFF_save_fm DFF_W3109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D119));
DFF_save_fm DFF_W3110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D129));
DFF_save_fm DFF_W3111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D209));
DFF_save_fm DFF_W3112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D219));
DFF_save_fm DFF_W3113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D229));
DFF_save_fm DFF_W3114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D00A));
DFF_save_fm DFF_W3115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D01A));
DFF_save_fm DFF_W3116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D02A));
DFF_save_fm DFF_W3117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D10A));
DFF_save_fm DFF_W3118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D11A));
DFF_save_fm DFF_W3119(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D12A));
DFF_save_fm DFF_W3120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D20A));
DFF_save_fm DFF_W3121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D21A));
DFF_save_fm DFF_W3122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D22A));
DFF_save_fm DFF_W3123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D00B));
DFF_save_fm DFF_W3124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D01B));
DFF_save_fm DFF_W3125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D02B));
DFF_save_fm DFF_W3126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D10B));
DFF_save_fm DFF_W3127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D11B));
DFF_save_fm DFF_W3128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D12B));
DFF_save_fm DFF_W3129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D20B));
DFF_save_fm DFF_W3130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D21B));
DFF_save_fm DFF_W3131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D22B));
DFF_save_fm DFF_W3132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D00C));
DFF_save_fm DFF_W3133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D01C));
DFF_save_fm DFF_W3134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D02C));
DFF_save_fm DFF_W3135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D10C));
DFF_save_fm DFF_W3136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D11C));
DFF_save_fm DFF_W3137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D12C));
DFF_save_fm DFF_W3138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D20C));
DFF_save_fm DFF_W3139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D21C));
DFF_save_fm DFF_W3140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D22C));
DFF_save_fm DFF_W3141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D00D));
DFF_save_fm DFF_W3142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D01D));
DFF_save_fm DFF_W3143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D02D));
DFF_save_fm DFF_W3144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D10D));
DFF_save_fm DFF_W3145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D11D));
DFF_save_fm DFF_W3146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D12D));
DFF_save_fm DFF_W3147(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D20D));
DFF_save_fm DFF_W3148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D21D));
DFF_save_fm DFF_W3149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D22D));
DFF_save_fm DFF_W3150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D00E));
DFF_save_fm DFF_W3151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D01E));
DFF_save_fm DFF_W3152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D02E));
DFF_save_fm DFF_W3153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D10E));
DFF_save_fm DFF_W3154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D11E));
DFF_save_fm DFF_W3155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D12E));
DFF_save_fm DFF_W3156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D20E));
DFF_save_fm DFF_W3157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D21E));
DFF_save_fm DFF_W3158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D22E));
DFF_save_fm DFF_W3159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D00F));
DFF_save_fm DFF_W3160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D01F));
DFF_save_fm DFF_W3161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D02F));
DFF_save_fm DFF_W3162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D10F));
DFF_save_fm DFF_W3163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3D11F));
DFF_save_fm DFF_W3164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D12F));
DFF_save_fm DFF_W3165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D20F));
DFF_save_fm DFF_W3166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D21F));
DFF_save_fm DFF_W3167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3D22F));
DFF_save_fm DFF_W3168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E000));
DFF_save_fm DFF_W3169(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E010));
DFF_save_fm DFF_W3170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E020));
DFF_save_fm DFF_W3171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E100));
DFF_save_fm DFF_W3172(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E110));
DFF_save_fm DFF_W3173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E120));
DFF_save_fm DFF_W3174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E200));
DFF_save_fm DFF_W3175(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E210));
DFF_save_fm DFF_W3176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E220));
DFF_save_fm DFF_W3177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E001));
DFF_save_fm DFF_W3178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E011));
DFF_save_fm DFF_W3179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E021));
DFF_save_fm DFF_W3180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E101));
DFF_save_fm DFF_W3181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E111));
DFF_save_fm DFF_W3182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E121));
DFF_save_fm DFF_W3183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E201));
DFF_save_fm DFF_W3184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E211));
DFF_save_fm DFF_W3185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E221));
DFF_save_fm DFF_W3186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E002));
DFF_save_fm DFF_W3187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E012));
DFF_save_fm DFF_W3188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E022));
DFF_save_fm DFF_W3189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E102));
DFF_save_fm DFF_W3190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E112));
DFF_save_fm DFF_W3191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E122));
DFF_save_fm DFF_W3192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E202));
DFF_save_fm DFF_W3193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E212));
DFF_save_fm DFF_W3194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E222));
DFF_save_fm DFF_W3195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E003));
DFF_save_fm DFF_W3196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E013));
DFF_save_fm DFF_W3197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E023));
DFF_save_fm DFF_W3198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E103));
DFF_save_fm DFF_W3199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E113));
DFF_save_fm DFF_W3200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E123));
DFF_save_fm DFF_W3201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E203));
DFF_save_fm DFF_W3202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E213));
DFF_save_fm DFF_W3203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E223));
DFF_save_fm DFF_W3204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E004));
DFF_save_fm DFF_W3205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E014));
DFF_save_fm DFF_W3206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E024));
DFF_save_fm DFF_W3207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E104));
DFF_save_fm DFF_W3208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E114));
DFF_save_fm DFF_W3209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E124));
DFF_save_fm DFF_W3210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E204));
DFF_save_fm DFF_W3211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E214));
DFF_save_fm DFF_W3212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E224));
DFF_save_fm DFF_W3213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E005));
DFF_save_fm DFF_W3214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E015));
DFF_save_fm DFF_W3215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E025));
DFF_save_fm DFF_W3216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E105));
DFF_save_fm DFF_W3217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E115));
DFF_save_fm DFF_W3218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E125));
DFF_save_fm DFF_W3219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E205));
DFF_save_fm DFF_W3220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E215));
DFF_save_fm DFF_W3221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E225));
DFF_save_fm DFF_W3222(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E006));
DFF_save_fm DFF_W3223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E016));
DFF_save_fm DFF_W3224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E026));
DFF_save_fm DFF_W3225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E106));
DFF_save_fm DFF_W3226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E116));
DFF_save_fm DFF_W3227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E126));
DFF_save_fm DFF_W3228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E206));
DFF_save_fm DFF_W3229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E216));
DFF_save_fm DFF_W3230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E226));
DFF_save_fm DFF_W3231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E007));
DFF_save_fm DFF_W3232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E017));
DFF_save_fm DFF_W3233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E027));
DFF_save_fm DFF_W3234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E107));
DFF_save_fm DFF_W3235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E117));
DFF_save_fm DFF_W3236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E127));
DFF_save_fm DFF_W3237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E207));
DFF_save_fm DFF_W3238(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E217));
DFF_save_fm DFF_W3239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E227));
DFF_save_fm DFF_W3240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E008));
DFF_save_fm DFF_W3241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E018));
DFF_save_fm DFF_W3242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E028));
DFF_save_fm DFF_W3243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E108));
DFF_save_fm DFF_W3244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E118));
DFF_save_fm DFF_W3245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E128));
DFF_save_fm DFF_W3246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E208));
DFF_save_fm DFF_W3247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E218));
DFF_save_fm DFF_W3248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E228));
DFF_save_fm DFF_W3249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E009));
DFF_save_fm DFF_W3250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E019));
DFF_save_fm DFF_W3251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E029));
DFF_save_fm DFF_W3252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E109));
DFF_save_fm DFF_W3253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E119));
DFF_save_fm DFF_W3254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E129));
DFF_save_fm DFF_W3255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E209));
DFF_save_fm DFF_W3256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E219));
DFF_save_fm DFF_W3257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E229));
DFF_save_fm DFF_W3258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E00A));
DFF_save_fm DFF_W3259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E01A));
DFF_save_fm DFF_W3260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E02A));
DFF_save_fm DFF_W3261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E10A));
DFF_save_fm DFF_W3262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E11A));
DFF_save_fm DFF_W3263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E12A));
DFF_save_fm DFF_W3264(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E20A));
DFF_save_fm DFF_W3265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E21A));
DFF_save_fm DFF_W3266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E22A));
DFF_save_fm DFF_W3267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E00B));
DFF_save_fm DFF_W3268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E01B));
DFF_save_fm DFF_W3269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E02B));
DFF_save_fm DFF_W3270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E10B));
DFF_save_fm DFF_W3271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E11B));
DFF_save_fm DFF_W3272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E12B));
DFF_save_fm DFF_W3273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E20B));
DFF_save_fm DFF_W3274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E21B));
DFF_save_fm DFF_W3275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E22B));
DFF_save_fm DFF_W3276(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E00C));
DFF_save_fm DFF_W3277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E01C));
DFF_save_fm DFF_W3278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E02C));
DFF_save_fm DFF_W3279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E10C));
DFF_save_fm DFF_W3280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E11C));
DFF_save_fm DFF_W3281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E12C));
DFF_save_fm DFF_W3282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E20C));
DFF_save_fm DFF_W3283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E21C));
DFF_save_fm DFF_W3284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E22C));
DFF_save_fm DFF_W3285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E00D));
DFF_save_fm DFF_W3286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E01D));
DFF_save_fm DFF_W3287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E02D));
DFF_save_fm DFF_W3288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E10D));
DFF_save_fm DFF_W3289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E11D));
DFF_save_fm DFF_W3290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E12D));
DFF_save_fm DFF_W3291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E20D));
DFF_save_fm DFF_W3292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E21D));
DFF_save_fm DFF_W3293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E22D));
DFF_save_fm DFF_W3294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E00E));
DFF_save_fm DFF_W3295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E01E));
DFF_save_fm DFF_W3296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E02E));
DFF_save_fm DFF_W3297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E10E));
DFF_save_fm DFF_W3298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E11E));
DFF_save_fm DFF_W3299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E12E));
DFF_save_fm DFF_W3300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E20E));
DFF_save_fm DFF_W3301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E21E));
DFF_save_fm DFF_W3302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E22E));
DFF_save_fm DFF_W3303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E00F));
DFF_save_fm DFF_W3304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E01F));
DFF_save_fm DFF_W3305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E02F));
DFF_save_fm DFF_W3306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E10F));
DFF_save_fm DFF_W3307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E11F));
DFF_save_fm DFF_W3308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E12F));
DFF_save_fm DFF_W3309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E20F));
DFF_save_fm DFF_W3310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3E21F));
DFF_save_fm DFF_W3311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3E22F));
DFF_save_fm DFF_W3312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F000));
DFF_save_fm DFF_W3313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F010));
DFF_save_fm DFF_W3314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F020));
DFF_save_fm DFF_W3315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F100));
DFF_save_fm DFF_W3316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F110));
DFF_save_fm DFF_W3317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F120));
DFF_save_fm DFF_W3318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F200));
DFF_save_fm DFF_W3319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F210));
DFF_save_fm DFF_W3320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F220));
DFF_save_fm DFF_W3321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F001));
DFF_save_fm DFF_W3322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F011));
DFF_save_fm DFF_W3323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F021));
DFF_save_fm DFF_W3324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F101));
DFF_save_fm DFF_W3325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F111));
DFF_save_fm DFF_W3326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F121));
DFF_save_fm DFF_W3327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F201));
DFF_save_fm DFF_W3328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F211));
DFF_save_fm DFF_W3329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F221));
DFF_save_fm DFF_W3330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F002));
DFF_save_fm DFF_W3331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F012));
DFF_save_fm DFF_W3332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F022));
DFF_save_fm DFF_W3333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F102));
DFF_save_fm DFF_W3334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F112));
DFF_save_fm DFF_W3335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F122));
DFF_save_fm DFF_W3336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F202));
DFF_save_fm DFF_W3337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F212));
DFF_save_fm DFF_W3338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F222));
DFF_save_fm DFF_W3339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F003));
DFF_save_fm DFF_W3340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F013));
DFF_save_fm DFF_W3341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F023));
DFF_save_fm DFF_W3342(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F103));
DFF_save_fm DFF_W3343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F113));
DFF_save_fm DFF_W3344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F123));
DFF_save_fm DFF_W3345(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F203));
DFF_save_fm DFF_W3346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F213));
DFF_save_fm DFF_W3347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F223));
DFF_save_fm DFF_W3348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F004));
DFF_save_fm DFF_W3349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F014));
DFF_save_fm DFF_W3350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F024));
DFF_save_fm DFF_W3351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F104));
DFF_save_fm DFF_W3352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F114));
DFF_save_fm DFF_W3353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F124));
DFF_save_fm DFF_W3354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F204));
DFF_save_fm DFF_W3355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F214));
DFF_save_fm DFF_W3356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F224));
DFF_save_fm DFF_W3357(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F005));
DFF_save_fm DFF_W3358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F015));
DFF_save_fm DFF_W3359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F025));
DFF_save_fm DFF_W3360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F105));
DFF_save_fm DFF_W3361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F115));
DFF_save_fm DFF_W3362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F125));
DFF_save_fm DFF_W3363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F205));
DFF_save_fm DFF_W3364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F215));
DFF_save_fm DFF_W3365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F225));
DFF_save_fm DFF_W3366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F006));
DFF_save_fm DFF_W3367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F016));
DFF_save_fm DFF_W3368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F026));
DFF_save_fm DFF_W3369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F106));
DFF_save_fm DFF_W3370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F116));
DFF_save_fm DFF_W3371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F126));
DFF_save_fm DFF_W3372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F206));
DFF_save_fm DFF_W3373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F216));
DFF_save_fm DFF_W3374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F226));
DFF_save_fm DFF_W3375(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F007));
DFF_save_fm DFF_W3376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F017));
DFF_save_fm DFF_W3377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F027));
DFF_save_fm DFF_W3378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F107));
DFF_save_fm DFF_W3379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F117));
DFF_save_fm DFF_W3380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F127));
DFF_save_fm DFF_W3381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F207));
DFF_save_fm DFF_W3382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F217));
DFF_save_fm DFF_W3383(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F227));
DFF_save_fm DFF_W3384(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F008));
DFF_save_fm DFF_W3385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F018));
DFF_save_fm DFF_W3386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F028));
DFF_save_fm DFF_W3387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F108));
DFF_save_fm DFF_W3388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F118));
DFF_save_fm DFF_W3389(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F128));
DFF_save_fm DFF_W3390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F208));
DFF_save_fm DFF_W3391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F218));
DFF_save_fm DFF_W3392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F228));
DFF_save_fm DFF_W3393(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F009));
DFF_save_fm DFF_W3394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F019));
DFF_save_fm DFF_W3395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F029));
DFF_save_fm DFF_W3396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F109));
DFF_save_fm DFF_W3397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F119));
DFF_save_fm DFF_W3398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F129));
DFF_save_fm DFF_W3399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F209));
DFF_save_fm DFF_W3400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F219));
DFF_save_fm DFF_W3401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F229));
DFF_save_fm DFF_W3402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F00A));
DFF_save_fm DFF_W3403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F01A));
DFF_save_fm DFF_W3404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F02A));
DFF_save_fm DFF_W3405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F10A));
DFF_save_fm DFF_W3406(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F11A));
DFF_save_fm DFF_W3407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F12A));
DFF_save_fm DFF_W3408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F20A));
DFF_save_fm DFF_W3409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F21A));
DFF_save_fm DFF_W3410(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F22A));
DFF_save_fm DFF_W3411(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F00B));
DFF_save_fm DFF_W3412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F01B));
DFF_save_fm DFF_W3413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F02B));
DFF_save_fm DFF_W3414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F10B));
DFF_save_fm DFF_W3415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F11B));
DFF_save_fm DFF_W3416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F12B));
DFF_save_fm DFF_W3417(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F20B));
DFF_save_fm DFF_W3418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F21B));
DFF_save_fm DFF_W3419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F22B));
DFF_save_fm DFF_W3420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F00C));
DFF_save_fm DFF_W3421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F01C));
DFF_save_fm DFF_W3422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F02C));
DFF_save_fm DFF_W3423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F10C));
DFF_save_fm DFF_W3424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F11C));
DFF_save_fm DFF_W3425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F12C));
DFF_save_fm DFF_W3426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F20C));
DFF_save_fm DFF_W3427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F21C));
DFF_save_fm DFF_W3428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F22C));
DFF_save_fm DFF_W3429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F00D));
DFF_save_fm DFF_W3430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F01D));
DFF_save_fm DFF_W3431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F02D));
DFF_save_fm DFF_W3432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F10D));
DFF_save_fm DFF_W3433(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F11D));
DFF_save_fm DFF_W3434(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F12D));
DFF_save_fm DFF_W3435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F20D));
DFF_save_fm DFF_W3436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F21D));
DFF_save_fm DFF_W3437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F22D));
DFF_save_fm DFF_W3438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F00E));
DFF_save_fm DFF_W3439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F01E));
DFF_save_fm DFF_W3440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F02E));
DFF_save_fm DFF_W3441(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F10E));
DFF_save_fm DFF_W3442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F11E));
DFF_save_fm DFF_W3443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F12E));
DFF_save_fm DFF_W3444(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F20E));
DFF_save_fm DFF_W3445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F21E));
DFF_save_fm DFF_W3446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F22E));
DFF_save_fm DFF_W3447(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F00F));
DFF_save_fm DFF_W3448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F01F));
DFF_save_fm DFF_W3449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F02F));
DFF_save_fm DFF_W3450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F10F));
DFF_save_fm DFF_W3451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F11F));
DFF_save_fm DFF_W3452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F12F));
DFF_save_fm DFF_W3453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F20F));
DFF_save_fm DFF_W3454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3F21F));
DFF_save_fm DFF_W3455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3F22F));
DFF_save_fm DFF_W3456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G000));
DFF_save_fm DFF_W3457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G010));
DFF_save_fm DFF_W3458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G020));
DFF_save_fm DFF_W3459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G100));
DFF_save_fm DFF_W3460(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G110));
DFF_save_fm DFF_W3461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G120));
DFF_save_fm DFF_W3462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G200));
DFF_save_fm DFF_W3463(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G210));
DFF_save_fm DFF_W3464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G220));
DFF_save_fm DFF_W3465(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G001));
DFF_save_fm DFF_W3466(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G011));
DFF_save_fm DFF_W3467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G021));
DFF_save_fm DFF_W3468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G101));
DFF_save_fm DFF_W3469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G111));
DFF_save_fm DFF_W3470(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G121));
DFF_save_fm DFF_W3471(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G201));
DFF_save_fm DFF_W3472(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G211));
DFF_save_fm DFF_W3473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G221));
DFF_save_fm DFF_W3474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G002));
DFF_save_fm DFF_W3475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G012));
DFF_save_fm DFF_W3476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G022));
DFF_save_fm DFF_W3477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G102));
DFF_save_fm DFF_W3478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G112));
DFF_save_fm DFF_W3479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G122));
DFF_save_fm DFF_W3480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G202));
DFF_save_fm DFF_W3481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G212));
DFF_save_fm DFF_W3482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G222));
DFF_save_fm DFF_W3483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G003));
DFF_save_fm DFF_W3484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G013));
DFF_save_fm DFF_W3485(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G023));
DFF_save_fm DFF_W3486(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G103));
DFF_save_fm DFF_W3487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G113));
DFF_save_fm DFF_W3488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G123));
DFF_save_fm DFF_W3489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G203));
DFF_save_fm DFF_W3490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G213));
DFF_save_fm DFF_W3491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G223));
DFF_save_fm DFF_W3492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G004));
DFF_save_fm DFF_W3493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G014));
DFF_save_fm DFF_W3494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G024));
DFF_save_fm DFF_W3495(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G104));
DFF_save_fm DFF_W3496(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G114));
DFF_save_fm DFF_W3497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G124));
DFF_save_fm DFF_W3498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G204));
DFF_save_fm DFF_W3499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G214));
DFF_save_fm DFF_W3500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G224));
DFF_save_fm DFF_W3501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G005));
DFF_save_fm DFF_W3502(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G015));
DFF_save_fm DFF_W3503(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G025));
DFF_save_fm DFF_W3504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G105));
DFF_save_fm DFF_W3505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G115));
DFF_save_fm DFF_W3506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G125));
DFF_save_fm DFF_W3507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G205));
DFF_save_fm DFF_W3508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G215));
DFF_save_fm DFF_W3509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G225));
DFF_save_fm DFF_W3510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G006));
DFF_save_fm DFF_W3511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G016));
DFF_save_fm DFF_W3512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G026));
DFF_save_fm DFF_W3513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G106));
DFF_save_fm DFF_W3514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G116));
DFF_save_fm DFF_W3515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G126));
DFF_save_fm DFF_W3516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G206));
DFF_save_fm DFF_W3517(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G216));
DFF_save_fm DFF_W3518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G226));
DFF_save_fm DFF_W3519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G007));
DFF_save_fm DFF_W3520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G017));
DFF_save_fm DFF_W3521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G027));
DFF_save_fm DFF_W3522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G107));
DFF_save_fm DFF_W3523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G117));
DFF_save_fm DFF_W3524(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G127));
DFF_save_fm DFF_W3525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G207));
DFF_save_fm DFF_W3526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G217));
DFF_save_fm DFF_W3527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G227));
DFF_save_fm DFF_W3528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G008));
DFF_save_fm DFF_W3529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G018));
DFF_save_fm DFF_W3530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G028));
DFF_save_fm DFF_W3531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G108));
DFF_save_fm DFF_W3532(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G118));
DFF_save_fm DFF_W3533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G128));
DFF_save_fm DFF_W3534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G208));
DFF_save_fm DFF_W3535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G218));
DFF_save_fm DFF_W3536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G228));
DFF_save_fm DFF_W3537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G009));
DFF_save_fm DFF_W3538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G019));
DFF_save_fm DFF_W3539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G029));
DFF_save_fm DFF_W3540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G109));
DFF_save_fm DFF_W3541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G119));
DFF_save_fm DFF_W3542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G129));
DFF_save_fm DFF_W3543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G209));
DFF_save_fm DFF_W3544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G219));
DFF_save_fm DFF_W3545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G229));
DFF_save_fm DFF_W3546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G00A));
DFF_save_fm DFF_W3547(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G01A));
DFF_save_fm DFF_W3548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G02A));
DFF_save_fm DFF_W3549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G10A));
DFF_save_fm DFF_W3550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G11A));
DFF_save_fm DFF_W3551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G12A));
DFF_save_fm DFF_W3552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G20A));
DFF_save_fm DFF_W3553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G21A));
DFF_save_fm DFF_W3554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G22A));
DFF_save_fm DFF_W3555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G00B));
DFF_save_fm DFF_W3556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G01B));
DFF_save_fm DFF_W3557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G02B));
DFF_save_fm DFF_W3558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G10B));
DFF_save_fm DFF_W3559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G11B));
DFF_save_fm DFF_W3560(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G12B));
DFF_save_fm DFF_W3561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G20B));
DFF_save_fm DFF_W3562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G21B));
DFF_save_fm DFF_W3563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G22B));
DFF_save_fm DFF_W3564(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G00C));
DFF_save_fm DFF_W3565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G01C));
DFF_save_fm DFF_W3566(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G02C));
DFF_save_fm DFF_W3567(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G10C));
DFF_save_fm DFF_W3568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G11C));
DFF_save_fm DFF_W3569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G12C));
DFF_save_fm DFF_W3570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G20C));
DFF_save_fm DFF_W3571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G21C));
DFF_save_fm DFF_W3572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G22C));
DFF_save_fm DFF_W3573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G00D));
DFF_save_fm DFF_W3574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G01D));
DFF_save_fm DFF_W3575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G02D));
DFF_save_fm DFF_W3576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G10D));
DFF_save_fm DFF_W3577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G11D));
DFF_save_fm DFF_W3578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G12D));
DFF_save_fm DFF_W3579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G20D));
DFF_save_fm DFF_W3580(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G21D));
DFF_save_fm DFF_W3581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G22D));
DFF_save_fm DFF_W3582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G00E));
DFF_save_fm DFF_W3583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G01E));
DFF_save_fm DFF_W3584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G02E));
DFF_save_fm DFF_W3585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G10E));
DFF_save_fm DFF_W3586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G11E));
DFF_save_fm DFF_W3587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G12E));
DFF_save_fm DFF_W3588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G20E));
DFF_save_fm DFF_W3589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G21E));
DFF_save_fm DFF_W3590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G22E));
DFF_save_fm DFF_W3591(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G00F));
DFF_save_fm DFF_W3592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G01F));
DFF_save_fm DFF_W3593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G02F));
DFF_save_fm DFF_W3594(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G10F));
DFF_save_fm DFF_W3595(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G11F));
DFF_save_fm DFF_W3596(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G12F));
DFF_save_fm DFF_W3597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G20F));
DFF_save_fm DFF_W3598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3G21F));
DFF_save_fm DFF_W3599(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3G22F));
DFF_save_fm DFF_W3600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H000));
DFF_save_fm DFF_W3601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H010));
DFF_save_fm DFF_W3602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H020));
DFF_save_fm DFF_W3603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H100));
DFF_save_fm DFF_W3604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H110));
DFF_save_fm DFF_W3605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H120));
DFF_save_fm DFF_W3606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H200));
DFF_save_fm DFF_W3607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H210));
DFF_save_fm DFF_W3608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H220));
DFF_save_fm DFF_W3609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H001));
DFF_save_fm DFF_W3610(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H011));
DFF_save_fm DFF_W3611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H021));
DFF_save_fm DFF_W3612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H101));
DFF_save_fm DFF_W3613(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H111));
DFF_save_fm DFF_W3614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H121));
DFF_save_fm DFF_W3615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H201));
DFF_save_fm DFF_W3616(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H211));
DFF_save_fm DFF_W3617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H221));
DFF_save_fm DFF_W3618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H002));
DFF_save_fm DFF_W3619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H012));
DFF_save_fm DFF_W3620(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H022));
DFF_save_fm DFF_W3621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H102));
DFF_save_fm DFF_W3622(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H112));
DFF_save_fm DFF_W3623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H122));
DFF_save_fm DFF_W3624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H202));
DFF_save_fm DFF_W3625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H212));
DFF_save_fm DFF_W3626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H222));
DFF_save_fm DFF_W3627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H003));
DFF_save_fm DFF_W3628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H013));
DFF_save_fm DFF_W3629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H023));
DFF_save_fm DFF_W3630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H103));
DFF_save_fm DFF_W3631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H113));
DFF_save_fm DFF_W3632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H123));
DFF_save_fm DFF_W3633(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H203));
DFF_save_fm DFF_W3634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H213));
DFF_save_fm DFF_W3635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H223));
DFF_save_fm DFF_W3636(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H004));
DFF_save_fm DFF_W3637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H014));
DFF_save_fm DFF_W3638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H024));
DFF_save_fm DFF_W3639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H104));
DFF_save_fm DFF_W3640(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H114));
DFF_save_fm DFF_W3641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H124));
DFF_save_fm DFF_W3642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H204));
DFF_save_fm DFF_W3643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H214));
DFF_save_fm DFF_W3644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H224));
DFF_save_fm DFF_W3645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H005));
DFF_save_fm DFF_W3646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H015));
DFF_save_fm DFF_W3647(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H025));
DFF_save_fm DFF_W3648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H105));
DFF_save_fm DFF_W3649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H115));
DFF_save_fm DFF_W3650(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H125));
DFF_save_fm DFF_W3651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H205));
DFF_save_fm DFF_W3652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H215));
DFF_save_fm DFF_W3653(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H225));
DFF_save_fm DFF_W3654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H006));
DFF_save_fm DFF_W3655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H016));
DFF_save_fm DFF_W3656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H026));
DFF_save_fm DFF_W3657(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H106));
DFF_save_fm DFF_W3658(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H116));
DFF_save_fm DFF_W3659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H126));
DFF_save_fm DFF_W3660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H206));
DFF_save_fm DFF_W3661(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H216));
DFF_save_fm DFF_W3662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H226));
DFF_save_fm DFF_W3663(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H007));
DFF_save_fm DFF_W3664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H017));
DFF_save_fm DFF_W3665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H027));
DFF_save_fm DFF_W3666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H107));
DFF_save_fm DFF_W3667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H117));
DFF_save_fm DFF_W3668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H127));
DFF_save_fm DFF_W3669(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H207));
DFF_save_fm DFF_W3670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H217));
DFF_save_fm DFF_W3671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H227));
DFF_save_fm DFF_W3672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H008));
DFF_save_fm DFF_W3673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H018));
DFF_save_fm DFF_W3674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H028));
DFF_save_fm DFF_W3675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H108));
DFF_save_fm DFF_W3676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H118));
DFF_save_fm DFF_W3677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H128));
DFF_save_fm DFF_W3678(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H208));
DFF_save_fm DFF_W3679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H218));
DFF_save_fm DFF_W3680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H228));
DFF_save_fm DFF_W3681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H009));
DFF_save_fm DFF_W3682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H019));
DFF_save_fm DFF_W3683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H029));
DFF_save_fm DFF_W3684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H109));
DFF_save_fm DFF_W3685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H119));
DFF_save_fm DFF_W3686(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H129));
DFF_save_fm DFF_W3687(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H209));
DFF_save_fm DFF_W3688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H219));
DFF_save_fm DFF_W3689(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H229));
DFF_save_fm DFF_W3690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H00A));
DFF_save_fm DFF_W3691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H01A));
DFF_save_fm DFF_W3692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H02A));
DFF_save_fm DFF_W3693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H10A));
DFF_save_fm DFF_W3694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H11A));
DFF_save_fm DFF_W3695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H12A));
DFF_save_fm DFF_W3696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H20A));
DFF_save_fm DFF_W3697(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H21A));
DFF_save_fm DFF_W3698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H22A));
DFF_save_fm DFF_W3699(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H00B));
DFF_save_fm DFF_W3700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H01B));
DFF_save_fm DFF_W3701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H02B));
DFF_save_fm DFF_W3702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H10B));
DFF_save_fm DFF_W3703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H11B));
DFF_save_fm DFF_W3704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H12B));
DFF_save_fm DFF_W3705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H20B));
DFF_save_fm DFF_W3706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H21B));
DFF_save_fm DFF_W3707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H22B));
DFF_save_fm DFF_W3708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H00C));
DFF_save_fm DFF_W3709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H01C));
DFF_save_fm DFF_W3710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H02C));
DFF_save_fm DFF_W3711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H10C));
DFF_save_fm DFF_W3712(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H11C));
DFF_save_fm DFF_W3713(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H12C));
DFF_save_fm DFF_W3714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H20C));
DFF_save_fm DFF_W3715(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H21C));
DFF_save_fm DFF_W3716(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H22C));
DFF_save_fm DFF_W3717(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H00D));
DFF_save_fm DFF_W3718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H01D));
DFF_save_fm DFF_W3719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H02D));
DFF_save_fm DFF_W3720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H10D));
DFF_save_fm DFF_W3721(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H11D));
DFF_save_fm DFF_W3722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H12D));
DFF_save_fm DFF_W3723(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H20D));
DFF_save_fm DFF_W3724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H21D));
DFF_save_fm DFF_W3725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H22D));
DFF_save_fm DFF_W3726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H00E));
DFF_save_fm DFF_W3727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H01E));
DFF_save_fm DFF_W3728(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H02E));
DFF_save_fm DFF_W3729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H10E));
DFF_save_fm DFF_W3730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H11E));
DFF_save_fm DFF_W3731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H12E));
DFF_save_fm DFF_W3732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H20E));
DFF_save_fm DFF_W3733(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H21E));
DFF_save_fm DFF_W3734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H22E));
DFF_save_fm DFF_W3735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H00F));
DFF_save_fm DFF_W3736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H01F));
DFF_save_fm DFF_W3737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H02F));
DFF_save_fm DFF_W3738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H10F));
DFF_save_fm DFF_W3739(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H11F));
DFF_save_fm DFF_W3740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H12F));
DFF_save_fm DFF_W3741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H20F));
DFF_save_fm DFF_W3742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3H21F));
DFF_save_fm DFF_W3743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3H22F));
DFF_save_fm DFF_W3744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I000));
DFF_save_fm DFF_W3745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I010));
DFF_save_fm DFF_W3746(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I020));
DFF_save_fm DFF_W3747(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I100));
DFF_save_fm DFF_W3748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I110));
DFF_save_fm DFF_W3749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I120));
DFF_save_fm DFF_W3750(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I200));
DFF_save_fm DFF_W3751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I210));
DFF_save_fm DFF_W3752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I220));
DFF_save_fm DFF_W3753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I001));
DFF_save_fm DFF_W3754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I011));
DFF_save_fm DFF_W3755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I021));
DFF_save_fm DFF_W3756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I101));
DFF_save_fm DFF_W3757(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I111));
DFF_save_fm DFF_W3758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I121));
DFF_save_fm DFF_W3759(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I201));
DFF_save_fm DFF_W3760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I211));
DFF_save_fm DFF_W3761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I221));
DFF_save_fm DFF_W3762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I002));
DFF_save_fm DFF_W3763(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I012));
DFF_save_fm DFF_W3764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I022));
DFF_save_fm DFF_W3765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I102));
DFF_save_fm DFF_W3766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I112));
DFF_save_fm DFF_W3767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I122));
DFF_save_fm DFF_W3768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I202));
DFF_save_fm DFF_W3769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I212));
DFF_save_fm DFF_W3770(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I222));
DFF_save_fm DFF_W3771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I003));
DFF_save_fm DFF_W3772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I013));
DFF_save_fm DFF_W3773(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I023));
DFF_save_fm DFF_W3774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I103));
DFF_save_fm DFF_W3775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I113));
DFF_save_fm DFF_W3776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I123));
DFF_save_fm DFF_W3777(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I203));
DFF_save_fm DFF_W3778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I213));
DFF_save_fm DFF_W3779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I223));
DFF_save_fm DFF_W3780(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I004));
DFF_save_fm DFF_W3781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I014));
DFF_save_fm DFF_W3782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I024));
DFF_save_fm DFF_W3783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I104));
DFF_save_fm DFF_W3784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I114));
DFF_save_fm DFF_W3785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I124));
DFF_save_fm DFF_W3786(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I204));
DFF_save_fm DFF_W3787(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I214));
DFF_save_fm DFF_W3788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I224));
DFF_save_fm DFF_W3789(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I005));
DFF_save_fm DFF_W3790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I015));
DFF_save_fm DFF_W3791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I025));
DFF_save_fm DFF_W3792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I105));
DFF_save_fm DFF_W3793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I115));
DFF_save_fm DFF_W3794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I125));
DFF_save_fm DFF_W3795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I205));
DFF_save_fm DFF_W3796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I215));
DFF_save_fm DFF_W3797(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I225));
DFF_save_fm DFF_W3798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I006));
DFF_save_fm DFF_W3799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I016));
DFF_save_fm DFF_W3800(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I026));
DFF_save_fm DFF_W3801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I106));
DFF_save_fm DFF_W3802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I116));
DFF_save_fm DFF_W3803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I126));
DFF_save_fm DFF_W3804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I206));
DFF_save_fm DFF_W3805(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I216));
DFF_save_fm DFF_W3806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I226));
DFF_save_fm DFF_W3807(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I007));
DFF_save_fm DFF_W3808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I017));
DFF_save_fm DFF_W3809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I027));
DFF_save_fm DFF_W3810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I107));
DFF_save_fm DFF_W3811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I117));
DFF_save_fm DFF_W3812(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I127));
DFF_save_fm DFF_W3813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I207));
DFF_save_fm DFF_W3814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I217));
DFF_save_fm DFF_W3815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I227));
DFF_save_fm DFF_W3816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I008));
DFF_save_fm DFF_W3817(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I018));
DFF_save_fm DFF_W3818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I028));
DFF_save_fm DFF_W3819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I108));
DFF_save_fm DFF_W3820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I118));
DFF_save_fm DFF_W3821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I128));
DFF_save_fm DFF_W3822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I208));
DFF_save_fm DFF_W3823(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I218));
DFF_save_fm DFF_W3824(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I228));
DFF_save_fm DFF_W3825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I009));
DFF_save_fm DFF_W3826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I019));
DFF_save_fm DFF_W3827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I029));
DFF_save_fm DFF_W3828(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I109));
DFF_save_fm DFF_W3829(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I119));
DFF_save_fm DFF_W3830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I129));
DFF_save_fm DFF_W3831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I209));
DFF_save_fm DFF_W3832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I219));
DFF_save_fm DFF_W3833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I229));
DFF_save_fm DFF_W3834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I00A));
DFF_save_fm DFF_W3835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I01A));
DFF_save_fm DFF_W3836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I02A));
DFF_save_fm DFF_W3837(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I10A));
DFF_save_fm DFF_W3838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I11A));
DFF_save_fm DFF_W3839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I12A));
DFF_save_fm DFF_W3840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I20A));
DFF_save_fm DFF_W3841(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I21A));
DFF_save_fm DFF_W3842(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I22A));
DFF_save_fm DFF_W3843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I00B));
DFF_save_fm DFF_W3844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I01B));
DFF_save_fm DFF_W3845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I02B));
DFF_save_fm DFF_W3846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I10B));
DFF_save_fm DFF_W3847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I11B));
DFF_save_fm DFF_W3848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I12B));
DFF_save_fm DFF_W3849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I20B));
DFF_save_fm DFF_W3850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I21B));
DFF_save_fm DFF_W3851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I22B));
DFF_save_fm DFF_W3852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I00C));
DFF_save_fm DFF_W3853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I01C));
DFF_save_fm DFF_W3854(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I02C));
DFF_save_fm DFF_W3855(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I10C));
DFF_save_fm DFF_W3856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I11C));
DFF_save_fm DFF_W3857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I12C));
DFF_save_fm DFF_W3858(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I20C));
DFF_save_fm DFF_W3859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I21C));
DFF_save_fm DFF_W3860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I22C));
DFF_save_fm DFF_W3861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I00D));
DFF_save_fm DFF_W3862(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I01D));
DFF_save_fm DFF_W3863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I02D));
DFF_save_fm DFF_W3864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I10D));
DFF_save_fm DFF_W3865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I11D));
DFF_save_fm DFF_W3866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I12D));
DFF_save_fm DFF_W3867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I20D));
DFF_save_fm DFF_W3868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I21D));
DFF_save_fm DFF_W3869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I22D));
DFF_save_fm DFF_W3870(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I00E));
DFF_save_fm DFF_W3871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I01E));
DFF_save_fm DFF_W3872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I02E));
DFF_save_fm DFF_W3873(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I10E));
DFF_save_fm DFF_W3874(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I11E));
DFF_save_fm DFF_W3875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I12E));
DFF_save_fm DFF_W3876(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I20E));
DFF_save_fm DFF_W3877(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I21E));
DFF_save_fm DFF_W3878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I22E));
DFF_save_fm DFF_W3879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I00F));
DFF_save_fm DFF_W3880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I01F));
DFF_save_fm DFF_W3881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I02F));
DFF_save_fm DFF_W3882(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I10F));
DFF_save_fm DFF_W3883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I11F));
DFF_save_fm DFF_W3884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I12F));
DFF_save_fm DFF_W3885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I20F));
DFF_save_fm DFF_W3886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3I21F));
DFF_save_fm DFF_W3887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3I22F));
DFF_save_fm DFF_W3888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J000));
DFF_save_fm DFF_W3889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J010));
DFF_save_fm DFF_W3890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J020));
DFF_save_fm DFF_W3891(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J100));
DFF_save_fm DFF_W3892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J110));
DFF_save_fm DFF_W3893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J120));
DFF_save_fm DFF_W3894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J200));
DFF_save_fm DFF_W3895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J210));
DFF_save_fm DFF_W3896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J220));
DFF_save_fm DFF_W3897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J001));
DFF_save_fm DFF_W3898(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J011));
DFF_save_fm DFF_W3899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J021));
DFF_save_fm DFF_W3900(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J101));
DFF_save_fm DFF_W3901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J111));
DFF_save_fm DFF_W3902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J121));
DFF_save_fm DFF_W3903(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J201));
DFF_save_fm DFF_W3904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J211));
DFF_save_fm DFF_W3905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J221));
DFF_save_fm DFF_W3906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J002));
DFF_save_fm DFF_W3907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J012));
DFF_save_fm DFF_W3908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J022));
DFF_save_fm DFF_W3909(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J102));
DFF_save_fm DFF_W3910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J112));
DFF_save_fm DFF_W3911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J122));
DFF_save_fm DFF_W3912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J202));
DFF_save_fm DFF_W3913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J212));
DFF_save_fm DFF_W3914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J222));
DFF_save_fm DFF_W3915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J003));
DFF_save_fm DFF_W3916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J013));
DFF_save_fm DFF_W3917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J023));
DFF_save_fm DFF_W3918(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J103));
DFF_save_fm DFF_W3919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J113));
DFF_save_fm DFF_W3920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J123));
DFF_save_fm DFF_W3921(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J203));
DFF_save_fm DFF_W3922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J213));
DFF_save_fm DFF_W3923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J223));
DFF_save_fm DFF_W3924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J004));
DFF_save_fm DFF_W3925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J014));
DFF_save_fm DFF_W3926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J024));
DFF_save_fm DFF_W3927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J104));
DFF_save_fm DFF_W3928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J114));
DFF_save_fm DFF_W3929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J124));
DFF_save_fm DFF_W3930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J204));
DFF_save_fm DFF_W3931(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J214));
DFF_save_fm DFF_W3932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J224));
DFF_save_fm DFF_W3933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J005));
DFF_save_fm DFF_W3934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J015));
DFF_save_fm DFF_W3935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J025));
DFF_save_fm DFF_W3936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J105));
DFF_save_fm DFF_W3937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J115));
DFF_save_fm DFF_W3938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J125));
DFF_save_fm DFF_W3939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J205));
DFF_save_fm DFF_W3940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J215));
DFF_save_fm DFF_W3941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J225));
DFF_save_fm DFF_W3942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J006));
DFF_save_fm DFF_W3943(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J016));
DFF_save_fm DFF_W3944(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J026));
DFF_save_fm DFF_W3945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J106));
DFF_save_fm DFF_W3946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J116));
DFF_save_fm DFF_W3947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J126));
DFF_save_fm DFF_W3948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J206));
DFF_save_fm DFF_W3949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J216));
DFF_save_fm DFF_W3950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J226));
DFF_save_fm DFF_W3951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J007));
DFF_save_fm DFF_W3952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J017));
DFF_save_fm DFF_W3953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J027));
DFF_save_fm DFF_W3954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J107));
DFF_save_fm DFF_W3955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J117));
DFF_save_fm DFF_W3956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J127));
DFF_save_fm DFF_W3957(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J207));
DFF_save_fm DFF_W3958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J217));
DFF_save_fm DFF_W3959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J227));
DFF_save_fm DFF_W3960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J008));
DFF_save_fm DFF_W3961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J018));
DFF_save_fm DFF_W3962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J028));
DFF_save_fm DFF_W3963(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J108));
DFF_save_fm DFF_W3964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J118));
DFF_save_fm DFF_W3965(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J128));
DFF_save_fm DFF_W3966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J208));
DFF_save_fm DFF_W3967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J218));
DFF_save_fm DFF_W3968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J228));
DFF_save_fm DFF_W3969(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J009));
DFF_save_fm DFF_W3970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J019));
DFF_save_fm DFF_W3971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J029));
DFF_save_fm DFF_W3972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J109));
DFF_save_fm DFF_W3973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J119));
DFF_save_fm DFF_W3974(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J129));
DFF_save_fm DFF_W3975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J209));
DFF_save_fm DFF_W3976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J219));
DFF_save_fm DFF_W3977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J229));
DFF_save_fm DFF_W3978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J00A));
DFF_save_fm DFF_W3979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J01A));
DFF_save_fm DFF_W3980(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J02A));
DFF_save_fm DFF_W3981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J10A));
DFF_save_fm DFF_W3982(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J11A));
DFF_save_fm DFF_W3983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J12A));
DFF_save_fm DFF_W3984(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J20A));
DFF_save_fm DFF_W3985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J21A));
DFF_save_fm DFF_W3986(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J22A));
DFF_save_fm DFF_W3987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J00B));
DFF_save_fm DFF_W3988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J01B));
DFF_save_fm DFF_W3989(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J02B));
DFF_save_fm DFF_W3990(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J10B));
DFF_save_fm DFF_W3991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J11B));
DFF_save_fm DFF_W3992(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J12B));
DFF_save_fm DFF_W3993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J20B));
DFF_save_fm DFF_W3994(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J21B));
DFF_save_fm DFF_W3995(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J22B));
DFF_save_fm DFF_W3996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J00C));
DFF_save_fm DFF_W3997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J01C));
DFF_save_fm DFF_W3998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J02C));
DFF_save_fm DFF_W3999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J10C));
DFF_save_fm DFF_W4000(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J11C));
DFF_save_fm DFF_W4001(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J12C));
DFF_save_fm DFF_W4002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J20C));
DFF_save_fm DFF_W4003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J21C));
DFF_save_fm DFF_W4004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J22C));
DFF_save_fm DFF_W4005(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J00D));
DFF_save_fm DFF_W4006(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J01D));
DFF_save_fm DFF_W4007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J02D));
DFF_save_fm DFF_W4008(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J10D));
DFF_save_fm DFF_W4009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J11D));
DFF_save_fm DFF_W4010(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J12D));
DFF_save_fm DFF_W4011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J20D));
DFF_save_fm DFF_W4012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J21D));
DFF_save_fm DFF_W4013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J22D));
DFF_save_fm DFF_W4014(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J00E));
DFF_save_fm DFF_W4015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J01E));
DFF_save_fm DFF_W4016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J02E));
DFF_save_fm DFF_W4017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J10E));
DFF_save_fm DFF_W4018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J11E));
DFF_save_fm DFF_W4019(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J12E));
DFF_save_fm DFF_W4020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J20E));
DFF_save_fm DFF_W4021(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J21E));
DFF_save_fm DFF_W4022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J22E));
DFF_save_fm DFF_W4023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J00F));
DFF_save_fm DFF_W4024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J01F));
DFF_save_fm DFF_W4025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J02F));
DFF_save_fm DFF_W4026(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J10F));
DFF_save_fm DFF_W4027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J11F));
DFF_save_fm DFF_W4028(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3J12F));
DFF_save_fm DFF_W4029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J20F));
DFF_save_fm DFF_W4030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J21F));
DFF_save_fm DFF_W4031(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3J22F));
DFF_save_fm DFF_W4032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K000));
DFF_save_fm DFF_W4033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K010));
DFF_save_fm DFF_W4034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K020));
DFF_save_fm DFF_W4035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K100));
DFF_save_fm DFF_W4036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K110));
DFF_save_fm DFF_W4037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K120));
DFF_save_fm DFF_W4038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K200));
DFF_save_fm DFF_W4039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K210));
DFF_save_fm DFF_W4040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K220));
DFF_save_fm DFF_W4041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K001));
DFF_save_fm DFF_W4042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K011));
DFF_save_fm DFF_W4043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K021));
DFF_save_fm DFF_W4044(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K101));
DFF_save_fm DFF_W4045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K111));
DFF_save_fm DFF_W4046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K121));
DFF_save_fm DFF_W4047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K201));
DFF_save_fm DFF_W4048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K211));
DFF_save_fm DFF_W4049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K221));
DFF_save_fm DFF_W4050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K002));
DFF_save_fm DFF_W4051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K012));
DFF_save_fm DFF_W4052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K022));
DFF_save_fm DFF_W4053(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K102));
DFF_save_fm DFF_W4054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K112));
DFF_save_fm DFF_W4055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K122));
DFF_save_fm DFF_W4056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K202));
DFF_save_fm DFF_W4057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K212));
DFF_save_fm DFF_W4058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K222));
DFF_save_fm DFF_W4059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K003));
DFF_save_fm DFF_W4060(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K013));
DFF_save_fm DFF_W4061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K023));
DFF_save_fm DFF_W4062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K103));
DFF_save_fm DFF_W4063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K113));
DFF_save_fm DFF_W4064(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K123));
DFF_save_fm DFF_W4065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K203));
DFF_save_fm DFF_W4066(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K213));
DFF_save_fm DFF_W4067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K223));
DFF_save_fm DFF_W4068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K004));
DFF_save_fm DFF_W4069(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K014));
DFF_save_fm DFF_W4070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K024));
DFF_save_fm DFF_W4071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K104));
DFF_save_fm DFF_W4072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K114));
DFF_save_fm DFF_W4073(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K124));
DFF_save_fm DFF_W4074(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K204));
DFF_save_fm DFF_W4075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K214));
DFF_save_fm DFF_W4076(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K224));
DFF_save_fm DFF_W4077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K005));
DFF_save_fm DFF_W4078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K015));
DFF_save_fm DFF_W4079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K025));
DFF_save_fm DFF_W4080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K105));
DFF_save_fm DFF_W4081(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K115));
DFF_save_fm DFF_W4082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K125));
DFF_save_fm DFF_W4083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K205));
DFF_save_fm DFF_W4084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K215));
DFF_save_fm DFF_W4085(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K225));
DFF_save_fm DFF_W4086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K006));
DFF_save_fm DFF_W4087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K016));
DFF_save_fm DFF_W4088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K026));
DFF_save_fm DFF_W4089(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K106));
DFF_save_fm DFF_W4090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K116));
DFF_save_fm DFF_W4091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K126));
DFF_save_fm DFF_W4092(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K206));
DFF_save_fm DFF_W4093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K216));
DFF_save_fm DFF_W4094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K226));
DFF_save_fm DFF_W4095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K007));
DFF_save_fm DFF_W4096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K017));
DFF_save_fm DFF_W4097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K027));
DFF_save_fm DFF_W4098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K107));
DFF_save_fm DFF_W4099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K117));
DFF_save_fm DFF_W4100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K127));
DFF_save_fm DFF_W4101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K207));
DFF_save_fm DFF_W4102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K217));
DFF_save_fm DFF_W4103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K227));
DFF_save_fm DFF_W4104(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K008));
DFF_save_fm DFF_W4105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K018));
DFF_save_fm DFF_W4106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K028));
DFF_save_fm DFF_W4107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K108));
DFF_save_fm DFF_W4108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K118));
DFF_save_fm DFF_W4109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K128));
DFF_save_fm DFF_W4110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K208));
DFF_save_fm DFF_W4111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K218));
DFF_save_fm DFF_W4112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K228));
DFF_save_fm DFF_W4113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K009));
DFF_save_fm DFF_W4114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K019));
DFF_save_fm DFF_W4115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K029));
DFF_save_fm DFF_W4116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K109));
DFF_save_fm DFF_W4117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K119));
DFF_save_fm DFF_W4118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K129));
DFF_save_fm DFF_W4119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K209));
DFF_save_fm DFF_W4120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K219));
DFF_save_fm DFF_W4121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K229));
DFF_save_fm DFF_W4122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K00A));
DFF_save_fm DFF_W4123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K01A));
DFF_save_fm DFF_W4124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K02A));
DFF_save_fm DFF_W4125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K10A));
DFF_save_fm DFF_W4126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K11A));
DFF_save_fm DFF_W4127(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K12A));
DFF_save_fm DFF_W4128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K20A));
DFF_save_fm DFF_W4129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K21A));
DFF_save_fm DFF_W4130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K22A));
DFF_save_fm DFF_W4131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K00B));
DFF_save_fm DFF_W4132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K01B));
DFF_save_fm DFF_W4133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K02B));
DFF_save_fm DFF_W4134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K10B));
DFF_save_fm DFF_W4135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K11B));
DFF_save_fm DFF_W4136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K12B));
DFF_save_fm DFF_W4137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K20B));
DFF_save_fm DFF_W4138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K21B));
DFF_save_fm DFF_W4139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K22B));
DFF_save_fm DFF_W4140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K00C));
DFF_save_fm DFF_W4141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K01C));
DFF_save_fm DFF_W4142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K02C));
DFF_save_fm DFF_W4143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K10C));
DFF_save_fm DFF_W4144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K11C));
DFF_save_fm DFF_W4145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K12C));
DFF_save_fm DFF_W4146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K20C));
DFF_save_fm DFF_W4147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K21C));
DFF_save_fm DFF_W4148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K22C));
DFF_save_fm DFF_W4149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K00D));
DFF_save_fm DFF_W4150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K01D));
DFF_save_fm DFF_W4151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K02D));
DFF_save_fm DFF_W4152(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K10D));
DFF_save_fm DFF_W4153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K11D));
DFF_save_fm DFF_W4154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K12D));
DFF_save_fm DFF_W4155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K20D));
DFF_save_fm DFF_W4156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K21D));
DFF_save_fm DFF_W4157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K22D));
DFF_save_fm DFF_W4158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K00E));
DFF_save_fm DFF_W4159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K01E));
DFF_save_fm DFF_W4160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K02E));
DFF_save_fm DFF_W4161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K10E));
DFF_save_fm DFF_W4162(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K11E));
DFF_save_fm DFF_W4163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K12E));
DFF_save_fm DFF_W4164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K20E));
DFF_save_fm DFF_W4165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K21E));
DFF_save_fm DFF_W4166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K22E));
DFF_save_fm DFF_W4167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K00F));
DFF_save_fm DFF_W4168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K01F));
DFF_save_fm DFF_W4169(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K02F));
DFF_save_fm DFF_W4170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K10F));
DFF_save_fm DFF_W4171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K11F));
DFF_save_fm DFF_W4172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3K12F));
DFF_save_fm DFF_W4173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K20F));
DFF_save_fm DFF_W4174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K21F));
DFF_save_fm DFF_W4175(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3K22F));
DFF_save_fm DFF_W4176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L000));
DFF_save_fm DFF_W4177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L010));
DFF_save_fm DFF_W4178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L020));
DFF_save_fm DFF_W4179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L100));
DFF_save_fm DFF_W4180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L110));
DFF_save_fm DFF_W4181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L120));
DFF_save_fm DFF_W4182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L200));
DFF_save_fm DFF_W4183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L210));
DFF_save_fm DFF_W4184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L220));
DFF_save_fm DFF_W4185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L001));
DFF_save_fm DFF_W4186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L011));
DFF_save_fm DFF_W4187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L021));
DFF_save_fm DFF_W4188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L101));
DFF_save_fm DFF_W4189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L111));
DFF_save_fm DFF_W4190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L121));
DFF_save_fm DFF_W4191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L201));
DFF_save_fm DFF_W4192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L211));
DFF_save_fm DFF_W4193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L221));
DFF_save_fm DFF_W4194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L002));
DFF_save_fm DFF_W4195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L012));
DFF_save_fm DFF_W4196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L022));
DFF_save_fm DFF_W4197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L102));
DFF_save_fm DFF_W4198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L112));
DFF_save_fm DFF_W4199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L122));
DFF_save_fm DFF_W4200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L202));
DFF_save_fm DFF_W4201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L212));
DFF_save_fm DFF_W4202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L222));
DFF_save_fm DFF_W4203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L003));
DFF_save_fm DFF_W4204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L013));
DFF_save_fm DFF_W4205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L023));
DFF_save_fm DFF_W4206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L103));
DFF_save_fm DFF_W4207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L113));
DFF_save_fm DFF_W4208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L123));
DFF_save_fm DFF_W4209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L203));
DFF_save_fm DFF_W4210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L213));
DFF_save_fm DFF_W4211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L223));
DFF_save_fm DFF_W4212(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L004));
DFF_save_fm DFF_W4213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L014));
DFF_save_fm DFF_W4214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L024));
DFF_save_fm DFF_W4215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L104));
DFF_save_fm DFF_W4216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L114));
DFF_save_fm DFF_W4217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L124));
DFF_save_fm DFF_W4218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L204));
DFF_save_fm DFF_W4219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L214));
DFF_save_fm DFF_W4220(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L224));
DFF_save_fm DFF_W4221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L005));
DFF_save_fm DFF_W4222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L015));
DFF_save_fm DFF_W4223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L025));
DFF_save_fm DFF_W4224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L105));
DFF_save_fm DFF_W4225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L115));
DFF_save_fm DFF_W4226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L125));
DFF_save_fm DFF_W4227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L205));
DFF_save_fm DFF_W4228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L215));
DFF_save_fm DFF_W4229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L225));
DFF_save_fm DFF_W4230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L006));
DFF_save_fm DFF_W4231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L016));
DFF_save_fm DFF_W4232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L026));
DFF_save_fm DFF_W4233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L106));
DFF_save_fm DFF_W4234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L116));
DFF_save_fm DFF_W4235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L126));
DFF_save_fm DFF_W4236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L206));
DFF_save_fm DFF_W4237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L216));
DFF_save_fm DFF_W4238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L226));
DFF_save_fm DFF_W4239(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L007));
DFF_save_fm DFF_W4240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L017));
DFF_save_fm DFF_W4241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L027));
DFF_save_fm DFF_W4242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L107));
DFF_save_fm DFF_W4243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L117));
DFF_save_fm DFF_W4244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L127));
DFF_save_fm DFF_W4245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L207));
DFF_save_fm DFF_W4246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L217));
DFF_save_fm DFF_W4247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L227));
DFF_save_fm DFF_W4248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L008));
DFF_save_fm DFF_W4249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L018));
DFF_save_fm DFF_W4250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L028));
DFF_save_fm DFF_W4251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L108));
DFF_save_fm DFF_W4252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L118));
DFF_save_fm DFF_W4253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L128));
DFF_save_fm DFF_W4254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L208));
DFF_save_fm DFF_W4255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L218));
DFF_save_fm DFF_W4256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L228));
DFF_save_fm DFF_W4257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L009));
DFF_save_fm DFF_W4258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L019));
DFF_save_fm DFF_W4259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L029));
DFF_save_fm DFF_W4260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L109));
DFF_save_fm DFF_W4261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L119));
DFF_save_fm DFF_W4262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L129));
DFF_save_fm DFF_W4263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L209));
DFF_save_fm DFF_W4264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L219));
DFF_save_fm DFF_W4265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L229));
DFF_save_fm DFF_W4266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L00A));
DFF_save_fm DFF_W4267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L01A));
DFF_save_fm DFF_W4268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L02A));
DFF_save_fm DFF_W4269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L10A));
DFF_save_fm DFF_W4270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L11A));
DFF_save_fm DFF_W4271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L12A));
DFF_save_fm DFF_W4272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L20A));
DFF_save_fm DFF_W4273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L21A));
DFF_save_fm DFF_W4274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L22A));
DFF_save_fm DFF_W4275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L00B));
DFF_save_fm DFF_W4276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L01B));
DFF_save_fm DFF_W4277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L02B));
DFF_save_fm DFF_W4278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L10B));
DFF_save_fm DFF_W4279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L11B));
DFF_save_fm DFF_W4280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L12B));
DFF_save_fm DFF_W4281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L20B));
DFF_save_fm DFF_W4282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L21B));
DFF_save_fm DFF_W4283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L22B));
DFF_save_fm DFF_W4284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L00C));
DFF_save_fm DFF_W4285(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L01C));
DFF_save_fm DFF_W4286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L02C));
DFF_save_fm DFF_W4287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L10C));
DFF_save_fm DFF_W4288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L11C));
DFF_save_fm DFF_W4289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L12C));
DFF_save_fm DFF_W4290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L20C));
DFF_save_fm DFF_W4291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L21C));
DFF_save_fm DFF_W4292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L22C));
DFF_save_fm DFF_W4293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L00D));
DFF_save_fm DFF_W4294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L01D));
DFF_save_fm DFF_W4295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L02D));
DFF_save_fm DFF_W4296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L10D));
DFF_save_fm DFF_W4297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L11D));
DFF_save_fm DFF_W4298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L12D));
DFF_save_fm DFF_W4299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L20D));
DFF_save_fm DFF_W4300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L21D));
DFF_save_fm DFF_W4301(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L22D));
DFF_save_fm DFF_W4302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L00E));
DFF_save_fm DFF_W4303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L01E));
DFF_save_fm DFF_W4304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L02E));
DFF_save_fm DFF_W4305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L10E));
DFF_save_fm DFF_W4306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L11E));
DFF_save_fm DFF_W4307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L12E));
DFF_save_fm DFF_W4308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L20E));
DFF_save_fm DFF_W4309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L21E));
DFF_save_fm DFF_W4310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L22E));
DFF_save_fm DFF_W4311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L00F));
DFF_save_fm DFF_W4312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L01F));
DFF_save_fm DFF_W4313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L02F));
DFF_save_fm DFF_W4314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L10F));
DFF_save_fm DFF_W4315(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L11F));
DFF_save_fm DFF_W4316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3L12F));
DFF_save_fm DFF_W4317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L20F));
DFF_save_fm DFF_W4318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L21F));
DFF_save_fm DFF_W4319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3L22F));
DFF_save_fm DFF_W4320(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M000));
DFF_save_fm DFF_W4321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M010));
DFF_save_fm DFF_W4322(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M020));
DFF_save_fm DFF_W4323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M100));
DFF_save_fm DFF_W4324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M110));
DFF_save_fm DFF_W4325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M120));
DFF_save_fm DFF_W4326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M200));
DFF_save_fm DFF_W4327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M210));
DFF_save_fm DFF_W4328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M220));
DFF_save_fm DFF_W4329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M001));
DFF_save_fm DFF_W4330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M011));
DFF_save_fm DFF_W4331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M021));
DFF_save_fm DFF_W4332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M101));
DFF_save_fm DFF_W4333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M111));
DFF_save_fm DFF_W4334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M121));
DFF_save_fm DFF_W4335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M201));
DFF_save_fm DFF_W4336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M211));
DFF_save_fm DFF_W4337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M221));
DFF_save_fm DFF_W4338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M002));
DFF_save_fm DFF_W4339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M012));
DFF_save_fm DFF_W4340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M022));
DFF_save_fm DFF_W4341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M102));
DFF_save_fm DFF_W4342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M112));
DFF_save_fm DFF_W4343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M122));
DFF_save_fm DFF_W4344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M202));
DFF_save_fm DFF_W4345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M212));
DFF_save_fm DFF_W4346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M222));
DFF_save_fm DFF_W4347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M003));
DFF_save_fm DFF_W4348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M013));
DFF_save_fm DFF_W4349(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M023));
DFF_save_fm DFF_W4350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M103));
DFF_save_fm DFF_W4351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M113));
DFF_save_fm DFF_W4352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M123));
DFF_save_fm DFF_W4353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M203));
DFF_save_fm DFF_W4354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M213));
DFF_save_fm DFF_W4355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M223));
DFF_save_fm DFF_W4356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M004));
DFF_save_fm DFF_W4357(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M014));
DFF_save_fm DFF_W4358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M024));
DFF_save_fm DFF_W4359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M104));
DFF_save_fm DFF_W4360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M114));
DFF_save_fm DFF_W4361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M124));
DFF_save_fm DFF_W4362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M204));
DFF_save_fm DFF_W4363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M214));
DFF_save_fm DFF_W4364(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M224));
DFF_save_fm DFF_W4365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M005));
DFF_save_fm DFF_W4366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M015));
DFF_save_fm DFF_W4367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M025));
DFF_save_fm DFF_W4368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M105));
DFF_save_fm DFF_W4369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M115));
DFF_save_fm DFF_W4370(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M125));
DFF_save_fm DFF_W4371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M205));
DFF_save_fm DFF_W4372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M215));
DFF_save_fm DFF_W4373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M225));
DFF_save_fm DFF_W4374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M006));
DFF_save_fm DFF_W4375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M016));
DFF_save_fm DFF_W4376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M026));
DFF_save_fm DFF_W4377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M106));
DFF_save_fm DFF_W4378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M116));
DFF_save_fm DFF_W4379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M126));
DFF_save_fm DFF_W4380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M206));
DFF_save_fm DFF_W4381(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M216));
DFF_save_fm DFF_W4382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M226));
DFF_save_fm DFF_W4383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M007));
DFF_save_fm DFF_W4384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M017));
DFF_save_fm DFF_W4385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M027));
DFF_save_fm DFF_W4386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M107));
DFF_save_fm DFF_W4387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M117));
DFF_save_fm DFF_W4388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M127));
DFF_save_fm DFF_W4389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M207));
DFF_save_fm DFF_W4390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M217));
DFF_save_fm DFF_W4391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M227));
DFF_save_fm DFF_W4392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M008));
DFF_save_fm DFF_W4393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M018));
DFF_save_fm DFF_W4394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M028));
DFF_save_fm DFF_W4395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M108));
DFF_save_fm DFF_W4396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M118));
DFF_save_fm DFF_W4397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M128));
DFF_save_fm DFF_W4398(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M208));
DFF_save_fm DFF_W4399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M218));
DFF_save_fm DFF_W4400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M228));
DFF_save_fm DFF_W4401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M009));
DFF_save_fm DFF_W4402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M019));
DFF_save_fm DFF_W4403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M029));
DFF_save_fm DFF_W4404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M109));
DFF_save_fm DFF_W4405(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M119));
DFF_save_fm DFF_W4406(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M129));
DFF_save_fm DFF_W4407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M209));
DFF_save_fm DFF_W4408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M219));
DFF_save_fm DFF_W4409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M229));
DFF_save_fm DFF_W4410(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M00A));
DFF_save_fm DFF_W4411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M01A));
DFF_save_fm DFF_W4412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M02A));
DFF_save_fm DFF_W4413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M10A));
DFF_save_fm DFF_W4414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M11A));
DFF_save_fm DFF_W4415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M12A));
DFF_save_fm DFF_W4416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M20A));
DFF_save_fm DFF_W4417(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M21A));
DFF_save_fm DFF_W4418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M22A));
DFF_save_fm DFF_W4419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M00B));
DFF_save_fm DFF_W4420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M01B));
DFF_save_fm DFF_W4421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M02B));
DFF_save_fm DFF_W4422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M10B));
DFF_save_fm DFF_W4423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M11B));
DFF_save_fm DFF_W4424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M12B));
DFF_save_fm DFF_W4425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M20B));
DFF_save_fm DFF_W4426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M21B));
DFF_save_fm DFF_W4427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M22B));
DFF_save_fm DFF_W4428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M00C));
DFF_save_fm DFF_W4429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M01C));
DFF_save_fm DFF_W4430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M02C));
DFF_save_fm DFF_W4431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M10C));
DFF_save_fm DFF_W4432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M11C));
DFF_save_fm DFF_W4433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M12C));
DFF_save_fm DFF_W4434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M20C));
DFF_save_fm DFF_W4435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M21C));
DFF_save_fm DFF_W4436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M22C));
DFF_save_fm DFF_W4437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M00D));
DFF_save_fm DFF_W4438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M01D));
DFF_save_fm DFF_W4439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M02D));
DFF_save_fm DFF_W4440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M10D));
DFF_save_fm DFF_W4441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M11D));
DFF_save_fm DFF_W4442(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M12D));
DFF_save_fm DFF_W4443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M20D));
DFF_save_fm DFF_W4444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M21D));
DFF_save_fm DFF_W4445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M22D));
DFF_save_fm DFF_W4446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M00E));
DFF_save_fm DFF_W4447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M01E));
DFF_save_fm DFF_W4448(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M02E));
DFF_save_fm DFF_W4449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M10E));
DFF_save_fm DFF_W4450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M11E));
DFF_save_fm DFF_W4451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M12E));
DFF_save_fm DFF_W4452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M20E));
DFF_save_fm DFF_W4453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M21E));
DFF_save_fm DFF_W4454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M22E));
DFF_save_fm DFF_W4455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M00F));
DFF_save_fm DFF_W4456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M01F));
DFF_save_fm DFF_W4457(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M02F));
DFF_save_fm DFF_W4458(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M10F));
DFF_save_fm DFF_W4459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M11F));
DFF_save_fm DFF_W4460(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M12F));
DFF_save_fm DFF_W4461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3M20F));
DFF_save_fm DFF_W4462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M21F));
DFF_save_fm DFF_W4463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3M22F));
DFF_save_fm DFF_W4464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N000));
DFF_save_fm DFF_W4465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N010));
DFF_save_fm DFF_W4466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N020));
DFF_save_fm DFF_W4467(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N100));
DFF_save_fm DFF_W4468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N110));
DFF_save_fm DFF_W4469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N120));
DFF_save_fm DFF_W4470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N200));
DFF_save_fm DFF_W4471(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N210));
DFF_save_fm DFF_W4472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N220));
DFF_save_fm DFF_W4473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N001));
DFF_save_fm DFF_W4474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N011));
DFF_save_fm DFF_W4475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N021));
DFF_save_fm DFF_W4476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N101));
DFF_save_fm DFF_W4477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N111));
DFF_save_fm DFF_W4478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N121));
DFF_save_fm DFF_W4479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N201));
DFF_save_fm DFF_W4480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N211));
DFF_save_fm DFF_W4481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N221));
DFF_save_fm DFF_W4482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N002));
DFF_save_fm DFF_W4483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N012));
DFF_save_fm DFF_W4484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N022));
DFF_save_fm DFF_W4485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N102));
DFF_save_fm DFF_W4486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N112));
DFF_save_fm DFF_W4487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N122));
DFF_save_fm DFF_W4488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N202));
DFF_save_fm DFF_W4489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N212));
DFF_save_fm DFF_W4490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N222));
DFF_save_fm DFF_W4491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N003));
DFF_save_fm DFF_W4492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N013));
DFF_save_fm DFF_W4493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N023));
DFF_save_fm DFF_W4494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N103));
DFF_save_fm DFF_W4495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N113));
DFF_save_fm DFF_W4496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N123));
DFF_save_fm DFF_W4497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N203));
DFF_save_fm DFF_W4498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N213));
DFF_save_fm DFF_W4499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N223));
DFF_save_fm DFF_W4500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N004));
DFF_save_fm DFF_W4501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N014));
DFF_save_fm DFF_W4502(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N024));
DFF_save_fm DFF_W4503(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N104));
DFF_save_fm DFF_W4504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N114));
DFF_save_fm DFF_W4505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N124));
DFF_save_fm DFF_W4506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N204));
DFF_save_fm DFF_W4507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N214));
DFF_save_fm DFF_W4508(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N224));
DFF_save_fm DFF_W4509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N005));
DFF_save_fm DFF_W4510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N015));
DFF_save_fm DFF_W4511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N025));
DFF_save_fm DFF_W4512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N105));
DFF_save_fm DFF_W4513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N115));
DFF_save_fm DFF_W4514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N125));
DFF_save_fm DFF_W4515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N205));
DFF_save_fm DFF_W4516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N215));
DFF_save_fm DFF_W4517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N225));
DFF_save_fm DFF_W4518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N006));
DFF_save_fm DFF_W4519(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N016));
DFF_save_fm DFF_W4520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N026));
DFF_save_fm DFF_W4521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N106));
DFF_save_fm DFF_W4522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N116));
DFF_save_fm DFF_W4523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N126));
DFF_save_fm DFF_W4524(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N206));
DFF_save_fm DFF_W4525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N216));
DFF_save_fm DFF_W4526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N226));
DFF_save_fm DFF_W4527(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N007));
DFF_save_fm DFF_W4528(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N017));
DFF_save_fm DFF_W4529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N027));
DFF_save_fm DFF_W4530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N107));
DFF_save_fm DFF_W4531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N117));
DFF_save_fm DFF_W4532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N127));
DFF_save_fm DFF_W4533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N207));
DFF_save_fm DFF_W4534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N217));
DFF_save_fm DFF_W4535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N227));
DFF_save_fm DFF_W4536(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N008));
DFF_save_fm DFF_W4537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N018));
DFF_save_fm DFF_W4538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N028));
DFF_save_fm DFF_W4539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N108));
DFF_save_fm DFF_W4540(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N118));
DFF_save_fm DFF_W4541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N128));
DFF_save_fm DFF_W4542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N208));
DFF_save_fm DFF_W4543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N218));
DFF_save_fm DFF_W4544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N228));
DFF_save_fm DFF_W4545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N009));
DFF_save_fm DFF_W4546(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N019));
DFF_save_fm DFF_W4547(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N029));
DFF_save_fm DFF_W4548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N109));
DFF_save_fm DFF_W4549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N119));
DFF_save_fm DFF_W4550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N129));
DFF_save_fm DFF_W4551(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N209));
DFF_save_fm DFF_W4552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N219));
DFF_save_fm DFF_W4553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N229));
DFF_save_fm DFF_W4554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N00A));
DFF_save_fm DFF_W4555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N01A));
DFF_save_fm DFF_W4556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N02A));
DFF_save_fm DFF_W4557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N10A));
DFF_save_fm DFF_W4558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N11A));
DFF_save_fm DFF_W4559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N12A));
DFF_save_fm DFF_W4560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N20A));
DFF_save_fm DFF_W4561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N21A));
DFF_save_fm DFF_W4562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N22A));
DFF_save_fm DFF_W4563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N00B));
DFF_save_fm DFF_W4564(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N01B));
DFF_save_fm DFF_W4565(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N02B));
DFF_save_fm DFF_W4566(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N10B));
DFF_save_fm DFF_W4567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N11B));
DFF_save_fm DFF_W4568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N12B));
DFF_save_fm DFF_W4569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N20B));
DFF_save_fm DFF_W4570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N21B));
DFF_save_fm DFF_W4571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N22B));
DFF_save_fm DFF_W4572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N00C));
DFF_save_fm DFF_W4573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N01C));
DFF_save_fm DFF_W4574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N02C));
DFF_save_fm DFF_W4575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N10C));
DFF_save_fm DFF_W4576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N11C));
DFF_save_fm DFF_W4577(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N12C));
DFF_save_fm DFF_W4578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N20C));
DFF_save_fm DFF_W4579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N21C));
DFF_save_fm DFF_W4580(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N22C));
DFF_save_fm DFF_W4581(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N00D));
DFF_save_fm DFF_W4582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N01D));
DFF_save_fm DFF_W4583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N02D));
DFF_save_fm DFF_W4584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N10D));
DFF_save_fm DFF_W4585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N11D));
DFF_save_fm DFF_W4586(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N12D));
DFF_save_fm DFF_W4587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N20D));
DFF_save_fm DFF_W4588(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N21D));
DFF_save_fm DFF_W4589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N22D));
DFF_save_fm DFF_W4590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N00E));
DFF_save_fm DFF_W4591(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N01E));
DFF_save_fm DFF_W4592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N02E));
DFF_save_fm DFF_W4593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N10E));
DFF_save_fm DFF_W4594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N11E));
DFF_save_fm DFF_W4595(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N12E));
DFF_save_fm DFF_W4596(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N20E));
DFF_save_fm DFF_W4597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N21E));
DFF_save_fm DFF_W4598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N22E));
DFF_save_fm DFF_W4599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N00F));
DFF_save_fm DFF_W4600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N01F));
DFF_save_fm DFF_W4601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N02F));
DFF_save_fm DFF_W4602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N10F));
DFF_save_fm DFF_W4603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N11F));
DFF_save_fm DFF_W4604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N12F));
DFF_save_fm DFF_W4605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3N20F));
DFF_save_fm DFF_W4606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N21F));
DFF_save_fm DFF_W4607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3N22F));
DFF_save_fm DFF_W4608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O000));
DFF_save_fm DFF_W4609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O010));
DFF_save_fm DFF_W4610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O020));
DFF_save_fm DFF_W4611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O100));
DFF_save_fm DFF_W4612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O110));
DFF_save_fm DFF_W4613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O120));
DFF_save_fm DFF_W4614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O200));
DFF_save_fm DFF_W4615(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O210));
DFF_save_fm DFF_W4616(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O220));
DFF_save_fm DFF_W4617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O001));
DFF_save_fm DFF_W4618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O011));
DFF_save_fm DFF_W4619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O021));
DFF_save_fm DFF_W4620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O101));
DFF_save_fm DFF_W4621(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O111));
DFF_save_fm DFF_W4622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O121));
DFF_save_fm DFF_W4623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O201));
DFF_save_fm DFF_W4624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O211));
DFF_save_fm DFF_W4625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O221));
DFF_save_fm DFF_W4626(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O002));
DFF_save_fm DFF_W4627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O012));
DFF_save_fm DFF_W4628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O022));
DFF_save_fm DFF_W4629(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O102));
DFF_save_fm DFF_W4630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O112));
DFF_save_fm DFF_W4631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O122));
DFF_save_fm DFF_W4632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O202));
DFF_save_fm DFF_W4633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O212));
DFF_save_fm DFF_W4634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O222));
DFF_save_fm DFF_W4635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O003));
DFF_save_fm DFF_W4636(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O013));
DFF_save_fm DFF_W4637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O023));
DFF_save_fm DFF_W4638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O103));
DFF_save_fm DFF_W4639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O113));
DFF_save_fm DFF_W4640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O123));
DFF_save_fm DFF_W4641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O203));
DFF_save_fm DFF_W4642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O213));
DFF_save_fm DFF_W4643(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O223));
DFF_save_fm DFF_W4644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O004));
DFF_save_fm DFF_W4645(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O014));
DFF_save_fm DFF_W4646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O024));
DFF_save_fm DFF_W4647(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O104));
DFF_save_fm DFF_W4648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O114));
DFF_save_fm DFF_W4649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O124));
DFF_save_fm DFF_W4650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O204));
DFF_save_fm DFF_W4651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O214));
DFF_save_fm DFF_W4652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O224));
DFF_save_fm DFF_W4653(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O005));
DFF_save_fm DFF_W4654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O015));
DFF_save_fm DFF_W4655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O025));
DFF_save_fm DFF_W4656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O105));
DFF_save_fm DFF_W4657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O115));
DFF_save_fm DFF_W4658(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O125));
DFF_save_fm DFF_W4659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O205));
DFF_save_fm DFF_W4660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O215));
DFF_save_fm DFF_W4661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O225));
DFF_save_fm DFF_W4662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O006));
DFF_save_fm DFF_W4663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O016));
DFF_save_fm DFF_W4664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O026));
DFF_save_fm DFF_W4665(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O106));
DFF_save_fm DFF_W4666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O116));
DFF_save_fm DFF_W4667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O126));
DFF_save_fm DFF_W4668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O206));
DFF_save_fm DFF_W4669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O216));
DFF_save_fm DFF_W4670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O226));
DFF_save_fm DFF_W4671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O007));
DFF_save_fm DFF_W4672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O017));
DFF_save_fm DFF_W4673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O027));
DFF_save_fm DFF_W4674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O107));
DFF_save_fm DFF_W4675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O117));
DFF_save_fm DFF_W4676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O127));
DFF_save_fm DFF_W4677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O207));
DFF_save_fm DFF_W4678(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O217));
DFF_save_fm DFF_W4679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O227));
DFF_save_fm DFF_W4680(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O008));
DFF_save_fm DFF_W4681(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O018));
DFF_save_fm DFF_W4682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O028));
DFF_save_fm DFF_W4683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O108));
DFF_save_fm DFF_W4684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O118));
DFF_save_fm DFF_W4685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O128));
DFF_save_fm DFF_W4686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O208));
DFF_save_fm DFF_W4687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O218));
DFF_save_fm DFF_W4688(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O228));
DFF_save_fm DFF_W4689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O009));
DFF_save_fm DFF_W4690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O019));
DFF_save_fm DFF_W4691(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O029));
DFF_save_fm DFF_W4692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O109));
DFF_save_fm DFF_W4693(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O119));
DFF_save_fm DFF_W4694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O129));
DFF_save_fm DFF_W4695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O209));
DFF_save_fm DFF_W4696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O219));
DFF_save_fm DFF_W4697(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O229));
DFF_save_fm DFF_W4698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O00A));
DFF_save_fm DFF_W4699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O01A));
DFF_save_fm DFF_W4700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O02A));
DFF_save_fm DFF_W4701(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O10A));
DFF_save_fm DFF_W4702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O11A));
DFF_save_fm DFF_W4703(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O12A));
DFF_save_fm DFF_W4704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O20A));
DFF_save_fm DFF_W4705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O21A));
DFF_save_fm DFF_W4706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O22A));
DFF_save_fm DFF_W4707(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O00B));
DFF_save_fm DFF_W4708(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O01B));
DFF_save_fm DFF_W4709(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O02B));
DFF_save_fm DFF_W4710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O10B));
DFF_save_fm DFF_W4711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O11B));
DFF_save_fm DFF_W4712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O12B));
DFF_save_fm DFF_W4713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O20B));
DFF_save_fm DFF_W4714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O21B));
DFF_save_fm DFF_W4715(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O22B));
DFF_save_fm DFF_W4716(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O00C));
DFF_save_fm DFF_W4717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O01C));
DFF_save_fm DFF_W4718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O02C));
DFF_save_fm DFF_W4719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O10C));
DFF_save_fm DFF_W4720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O11C));
DFF_save_fm DFF_W4721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O12C));
DFF_save_fm DFF_W4722(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O20C));
DFF_save_fm DFF_W4723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O21C));
DFF_save_fm DFF_W4724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O22C));
DFF_save_fm DFF_W4725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O00D));
DFF_save_fm DFF_W4726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O01D));
DFF_save_fm DFF_W4727(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O02D));
DFF_save_fm DFF_W4728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O10D));
DFF_save_fm DFF_W4729(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O11D));
DFF_save_fm DFF_W4730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O12D));
DFF_save_fm DFF_W4731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O20D));
DFF_save_fm DFF_W4732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O21D));
DFF_save_fm DFF_W4733(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O22D));
DFF_save_fm DFF_W4734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O00E));
DFF_save_fm DFF_W4735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O01E));
DFF_save_fm DFF_W4736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O02E));
DFF_save_fm DFF_W4737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O10E));
DFF_save_fm DFF_W4738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O11E));
DFF_save_fm DFF_W4739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O12E));
DFF_save_fm DFF_W4740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O20E));
DFF_save_fm DFF_W4741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O21E));
DFF_save_fm DFF_W4742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O22E));
DFF_save_fm DFF_W4743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O00F));
DFF_save_fm DFF_W4744(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O01F));
DFF_save_fm DFF_W4745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O02F));
DFF_save_fm DFF_W4746(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O10F));
DFF_save_fm DFF_W4747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O11F));
DFF_save_fm DFF_W4748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O12F));
DFF_save_fm DFF_W4749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3O20F));
DFF_save_fm DFF_W4750(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O21F));
DFF_save_fm DFF_W4751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3O22F));
DFF_save_fm DFF_W4752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P000));
DFF_save_fm DFF_W4753(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P010));
DFF_save_fm DFF_W4754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P020));
DFF_save_fm DFF_W4755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P100));
DFF_save_fm DFF_W4756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P110));
DFF_save_fm DFF_W4757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P120));
DFF_save_fm DFF_W4758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P200));
DFF_save_fm DFF_W4759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P210));
DFF_save_fm DFF_W4760(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P220));
DFF_save_fm DFF_W4761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P001));
DFF_save_fm DFF_W4762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P011));
DFF_save_fm DFF_W4763(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P021));
DFF_save_fm DFF_W4764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P101));
DFF_save_fm DFF_W4765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P111));
DFF_save_fm DFF_W4766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P121));
DFF_save_fm DFF_W4767(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P201));
DFF_save_fm DFF_W4768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P211));
DFF_save_fm DFF_W4769(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P221));
DFF_save_fm DFF_W4770(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P002));
DFF_save_fm DFF_W4771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P012));
DFF_save_fm DFF_W4772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P022));
DFF_save_fm DFF_W4773(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P102));
DFF_save_fm DFF_W4774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P112));
DFF_save_fm DFF_W4775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P122));
DFF_save_fm DFF_W4776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P202));
DFF_save_fm DFF_W4777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P212));
DFF_save_fm DFF_W4778(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P222));
DFF_save_fm DFF_W4779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P003));
DFF_save_fm DFF_W4780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P013));
DFF_save_fm DFF_W4781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P023));
DFF_save_fm DFF_W4782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P103));
DFF_save_fm DFF_W4783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P113));
DFF_save_fm DFF_W4784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P123));
DFF_save_fm DFF_W4785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P203));
DFF_save_fm DFF_W4786(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P213));
DFF_save_fm DFF_W4787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P223));
DFF_save_fm DFF_W4788(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P004));
DFF_save_fm DFF_W4789(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P014));
DFF_save_fm DFF_W4790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P024));
DFF_save_fm DFF_W4791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P104));
DFF_save_fm DFF_W4792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P114));
DFF_save_fm DFF_W4793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P124));
DFF_save_fm DFF_W4794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P204));
DFF_save_fm DFF_W4795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P214));
DFF_save_fm DFF_W4796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P224));
DFF_save_fm DFF_W4797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P005));
DFF_save_fm DFF_W4798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P015));
DFF_save_fm DFF_W4799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P025));
DFF_save_fm DFF_W4800(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P105));
DFF_save_fm DFF_W4801(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P115));
DFF_save_fm DFF_W4802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P125));
DFF_save_fm DFF_W4803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P205));
DFF_save_fm DFF_W4804(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P215));
DFF_save_fm DFF_W4805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P225));
DFF_save_fm DFF_W4806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P006));
DFF_save_fm DFF_W4807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P016));
DFF_save_fm DFF_W4808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P026));
DFF_save_fm DFF_W4809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P106));
DFF_save_fm DFF_W4810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P116));
DFF_save_fm DFF_W4811(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P126));
DFF_save_fm DFF_W4812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P206));
DFF_save_fm DFF_W4813(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P216));
DFF_save_fm DFF_W4814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P226));
DFF_save_fm DFF_W4815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P007));
DFF_save_fm DFF_W4816(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P017));
DFF_save_fm DFF_W4817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P027));
DFF_save_fm DFF_W4818(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P107));
DFF_save_fm DFF_W4819(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P117));
DFF_save_fm DFF_W4820(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P127));
DFF_save_fm DFF_W4821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P207));
DFF_save_fm DFF_W4822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P217));
DFF_save_fm DFF_W4823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P227));
DFF_save_fm DFF_W4824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P008));
DFF_save_fm DFF_W4825(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P018));
DFF_save_fm DFF_W4826(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P028));
DFF_save_fm DFF_W4827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P108));
DFF_save_fm DFF_W4828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P118));
DFF_save_fm DFF_W4829(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P128));
DFF_save_fm DFF_W4830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P208));
DFF_save_fm DFF_W4831(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P218));
DFF_save_fm DFF_W4832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P228));
DFF_save_fm DFF_W4833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P009));
DFF_save_fm DFF_W4834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P019));
DFF_save_fm DFF_W4835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P029));
DFF_save_fm DFF_W4836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P109));
DFF_save_fm DFF_W4837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P119));
DFF_save_fm DFF_W4838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P129));
DFF_save_fm DFF_W4839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P209));
DFF_save_fm DFF_W4840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P219));
DFF_save_fm DFF_W4841(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P229));
DFF_save_fm DFF_W4842(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P00A));
DFF_save_fm DFF_W4843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P01A));
DFF_save_fm DFF_W4844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P02A));
DFF_save_fm DFF_W4845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P10A));
DFF_save_fm DFF_W4846(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P11A));
DFF_save_fm DFF_W4847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P12A));
DFF_save_fm DFF_W4848(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P20A));
DFF_save_fm DFF_W4849(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P21A));
DFF_save_fm DFF_W4850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P22A));
DFF_save_fm DFF_W4851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P00B));
DFF_save_fm DFF_W4852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P01B));
DFF_save_fm DFF_W4853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P02B));
DFF_save_fm DFF_W4854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P10B));
DFF_save_fm DFF_W4855(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P11B));
DFF_save_fm DFF_W4856(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P12B));
DFF_save_fm DFF_W4857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P20B));
DFF_save_fm DFF_W4858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P21B));
DFF_save_fm DFF_W4859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P22B));
DFF_save_fm DFF_W4860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P00C));
DFF_save_fm DFF_W4861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P01C));
DFF_save_fm DFF_W4862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P02C));
DFF_save_fm DFF_W4863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P10C));
DFF_save_fm DFF_W4864(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P11C));
DFF_save_fm DFF_W4865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P12C));
DFF_save_fm DFF_W4866(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P20C));
DFF_save_fm DFF_W4867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P21C));
DFF_save_fm DFF_W4868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P22C));
DFF_save_fm DFF_W4869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P00D));
DFF_save_fm DFF_W4870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P01D));
DFF_save_fm DFF_W4871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P02D));
DFF_save_fm DFF_W4872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P10D));
DFF_save_fm DFF_W4873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P11D));
DFF_save_fm DFF_W4874(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P12D));
DFF_save_fm DFF_W4875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P20D));
DFF_save_fm DFF_W4876(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P21D));
DFF_save_fm DFF_W4877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P22D));
DFF_save_fm DFF_W4878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P00E));
DFF_save_fm DFF_W4879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P01E));
DFF_save_fm DFF_W4880(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P02E));
DFF_save_fm DFF_W4881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P10E));
DFF_save_fm DFF_W4882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P11E));
DFF_save_fm DFF_W4883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P12E));
DFF_save_fm DFF_W4884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P20E));
DFF_save_fm DFF_W4885(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P21E));
DFF_save_fm DFF_W4886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P22E));
DFF_save_fm DFF_W4887(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P00F));
DFF_save_fm DFF_W4888(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P01F));
DFF_save_fm DFF_W4889(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P02F));
DFF_save_fm DFF_W4890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P10F));
DFF_save_fm DFF_W4891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P11F));
DFF_save_fm DFF_W4892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3P12F));
DFF_save_fm DFF_W4893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P20F));
DFF_save_fm DFF_W4894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P21F));
DFF_save_fm DFF_W4895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3P22F));
DFF_save_fm DFF_W4896(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q000));
DFF_save_fm DFF_W4897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q010));
DFF_save_fm DFF_W4898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q020));
DFF_save_fm DFF_W4899(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q100));
DFF_save_fm DFF_W4900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q110));
DFF_save_fm DFF_W4901(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q120));
DFF_save_fm DFF_W4902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q200));
DFF_save_fm DFF_W4903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q210));
DFF_save_fm DFF_W4904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q220));
DFF_save_fm DFF_W4905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q001));
DFF_save_fm DFF_W4906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q011));
DFF_save_fm DFF_W4907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q021));
DFF_save_fm DFF_W4908(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q101));
DFF_save_fm DFF_W4909(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q111));
DFF_save_fm DFF_W4910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q121));
DFF_save_fm DFF_W4911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q201));
DFF_save_fm DFF_W4912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q211));
DFF_save_fm DFF_W4913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q221));
DFF_save_fm DFF_W4914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q002));
DFF_save_fm DFF_W4915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q012));
DFF_save_fm DFF_W4916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q022));
DFF_save_fm DFF_W4917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q102));
DFF_save_fm DFF_W4918(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q112));
DFF_save_fm DFF_W4919(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q122));
DFF_save_fm DFF_W4920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q202));
DFF_save_fm DFF_W4921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q212));
DFF_save_fm DFF_W4922(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q222));
DFF_save_fm DFF_W4923(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q003));
DFF_save_fm DFF_W4924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q013));
DFF_save_fm DFF_W4925(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q023));
DFF_save_fm DFF_W4926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q103));
DFF_save_fm DFF_W4927(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q113));
DFF_save_fm DFF_W4928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q123));
DFF_save_fm DFF_W4929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q203));
DFF_save_fm DFF_W4930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q213));
DFF_save_fm DFF_W4931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q223));
DFF_save_fm DFF_W4932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q004));
DFF_save_fm DFF_W4933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q014));
DFF_save_fm DFF_W4934(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q024));
DFF_save_fm DFF_W4935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q104));
DFF_save_fm DFF_W4936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q114));
DFF_save_fm DFF_W4937(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q124));
DFF_save_fm DFF_W4938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q204));
DFF_save_fm DFF_W4939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q214));
DFF_save_fm DFF_W4940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q224));
DFF_save_fm DFF_W4941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q005));
DFF_save_fm DFF_W4942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q015));
DFF_save_fm DFF_W4943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q025));
DFF_save_fm DFF_W4944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q105));
DFF_save_fm DFF_W4945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q115));
DFF_save_fm DFF_W4946(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q125));
DFF_save_fm DFF_W4947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q205));
DFF_save_fm DFF_W4948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q215));
DFF_save_fm DFF_W4949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q225));
DFF_save_fm DFF_W4950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q006));
DFF_save_fm DFF_W4951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q016));
DFF_save_fm DFF_W4952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q026));
DFF_save_fm DFF_W4953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q106));
DFF_save_fm DFF_W4954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q116));
DFF_save_fm DFF_W4955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q126));
DFF_save_fm DFF_W4956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q206));
DFF_save_fm DFF_W4957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q216));
DFF_save_fm DFF_W4958(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q226));
DFF_save_fm DFF_W4959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q007));
DFF_save_fm DFF_W4960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q017));
DFF_save_fm DFF_W4961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q027));
DFF_save_fm DFF_W4962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q107));
DFF_save_fm DFF_W4963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q117));
DFF_save_fm DFF_W4964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q127));
DFF_save_fm DFF_W4965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q207));
DFF_save_fm DFF_W4966(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q217));
DFF_save_fm DFF_W4967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q227));
DFF_save_fm DFF_W4968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q008));
DFF_save_fm DFF_W4969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q018));
DFF_save_fm DFF_W4970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q028));
DFF_save_fm DFF_W4971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q108));
DFF_save_fm DFF_W4972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q118));
DFF_save_fm DFF_W4973(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q128));
DFF_save_fm DFF_W4974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q208));
DFF_save_fm DFF_W4975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q218));
DFF_save_fm DFF_W4976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q228));
DFF_save_fm DFF_W4977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q009));
DFF_save_fm DFF_W4978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q019));
DFF_save_fm DFF_W4979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q029));
DFF_save_fm DFF_W4980(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q109));
DFF_save_fm DFF_W4981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q119));
DFF_save_fm DFF_W4982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q129));
DFF_save_fm DFF_W4983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q209));
DFF_save_fm DFF_W4984(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q219));
DFF_save_fm DFF_W4985(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q229));
DFF_save_fm DFF_W4986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q00A));
DFF_save_fm DFF_W4987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q01A));
DFF_save_fm DFF_W4988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q02A));
DFF_save_fm DFF_W4989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q10A));
DFF_save_fm DFF_W4990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q11A));
DFF_save_fm DFF_W4991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q12A));
DFF_save_fm DFF_W4992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q20A));
DFF_save_fm DFF_W4993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q21A));
DFF_save_fm DFF_W4994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q22A));
DFF_save_fm DFF_W4995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q00B));
DFF_save_fm DFF_W4996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q01B));
DFF_save_fm DFF_W4997(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q02B));
DFF_save_fm DFF_W4998(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q10B));
DFF_save_fm DFF_W4999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q11B));
DFF_save_fm DFF_W5000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q12B));
DFF_save_fm DFF_W5001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q20B));
DFF_save_fm DFF_W5002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q21B));
DFF_save_fm DFF_W5003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q22B));
DFF_save_fm DFF_W5004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q00C));
DFF_save_fm DFF_W5005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q01C));
DFF_save_fm DFF_W5006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q02C));
DFF_save_fm DFF_W5007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q10C));
DFF_save_fm DFF_W5008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q11C));
DFF_save_fm DFF_W5009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q12C));
DFF_save_fm DFF_W5010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q20C));
DFF_save_fm DFF_W5011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q21C));
DFF_save_fm DFF_W5012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q22C));
DFF_save_fm DFF_W5013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q00D));
DFF_save_fm DFF_W5014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q01D));
DFF_save_fm DFF_W5015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q02D));
DFF_save_fm DFF_W5016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q10D));
DFF_save_fm DFF_W5017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q11D));
DFF_save_fm DFF_W5018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q12D));
DFF_save_fm DFF_W5019(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q20D));
DFF_save_fm DFF_W5020(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q21D));
DFF_save_fm DFF_W5021(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q22D));
DFF_save_fm DFF_W5022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q00E));
DFF_save_fm DFF_W5023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q01E));
DFF_save_fm DFF_W5024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q02E));
DFF_save_fm DFF_W5025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q10E));
DFF_save_fm DFF_W5026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q11E));
DFF_save_fm DFF_W5027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q12E));
DFF_save_fm DFF_W5028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q20E));
DFF_save_fm DFF_W5029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q21E));
DFF_save_fm DFF_W5030(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q22E));
DFF_save_fm DFF_W5031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q00F));
DFF_save_fm DFF_W5032(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q01F));
DFF_save_fm DFF_W5033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q02F));
DFF_save_fm DFF_W5034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q10F));
DFF_save_fm DFF_W5035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3Q11F));
DFF_save_fm DFF_W5036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q12F));
DFF_save_fm DFF_W5037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q20F));
DFF_save_fm DFF_W5038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q21F));
DFF_save_fm DFF_W5039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3Q22F));
DFF_save_fm DFF_W5040(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R000));
DFF_save_fm DFF_W5041(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R010));
DFF_save_fm DFF_W5042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R020));
DFF_save_fm DFF_W5043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R100));
DFF_save_fm DFF_W5044(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R110));
DFF_save_fm DFF_W5045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R120));
DFF_save_fm DFF_W5046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R200));
DFF_save_fm DFF_W5047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R210));
DFF_save_fm DFF_W5048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R220));
DFF_save_fm DFF_W5049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R001));
DFF_save_fm DFF_W5050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R011));
DFF_save_fm DFF_W5051(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R021));
DFF_save_fm DFF_W5052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R101));
DFF_save_fm DFF_W5053(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R111));
DFF_save_fm DFF_W5054(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R121));
DFF_save_fm DFF_W5055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R201));
DFF_save_fm DFF_W5056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R211));
DFF_save_fm DFF_W5057(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R221));
DFF_save_fm DFF_W5058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R002));
DFF_save_fm DFF_W5059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R012));
DFF_save_fm DFF_W5060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R022));
DFF_save_fm DFF_W5061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R102));
DFF_save_fm DFF_W5062(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R112));
DFF_save_fm DFF_W5063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R122));
DFF_save_fm DFF_W5064(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R202));
DFF_save_fm DFF_W5065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R212));
DFF_save_fm DFF_W5066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R222));
DFF_save_fm DFF_W5067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R003));
DFF_save_fm DFF_W5068(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R013));
DFF_save_fm DFF_W5069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R023));
DFF_save_fm DFF_W5070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R103));
DFF_save_fm DFF_W5071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R113));
DFF_save_fm DFF_W5072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R123));
DFF_save_fm DFF_W5073(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R203));
DFF_save_fm DFF_W5074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R213));
DFF_save_fm DFF_W5075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R223));
DFF_save_fm DFF_W5076(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R004));
DFF_save_fm DFF_W5077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R014));
DFF_save_fm DFF_W5078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R024));
DFF_save_fm DFF_W5079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R104));
DFF_save_fm DFF_W5080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R114));
DFF_save_fm DFF_W5081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R124));
DFF_save_fm DFF_W5082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R204));
DFF_save_fm DFF_W5083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R214));
DFF_save_fm DFF_W5084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R224));
DFF_save_fm DFF_W5085(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R005));
DFF_save_fm DFF_W5086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R015));
DFF_save_fm DFF_W5087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R025));
DFF_save_fm DFF_W5088(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R105));
DFF_save_fm DFF_W5089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R115));
DFF_save_fm DFF_W5090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R125));
DFF_save_fm DFF_W5091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R205));
DFF_save_fm DFF_W5092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R215));
DFF_save_fm DFF_W5093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R225));
DFF_save_fm DFF_W5094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R006));
DFF_save_fm DFF_W5095(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R016));
DFF_save_fm DFF_W5096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R026));
DFF_save_fm DFF_W5097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R106));
DFF_save_fm DFF_W5098(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R116));
DFF_save_fm DFF_W5099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R126));
DFF_save_fm DFF_W5100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R206));
DFF_save_fm DFF_W5101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R216));
DFF_save_fm DFF_W5102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R226));
DFF_save_fm DFF_W5103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R007));
DFF_save_fm DFF_W5104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R017));
DFF_save_fm DFF_W5105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R027));
DFF_save_fm DFF_W5106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R107));
DFF_save_fm DFF_W5107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R117));
DFF_save_fm DFF_W5108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R127));
DFF_save_fm DFF_W5109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R207));
DFF_save_fm DFF_W5110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R217));
DFF_save_fm DFF_W5111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R227));
DFF_save_fm DFF_W5112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R008));
DFF_save_fm DFF_W5113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R018));
DFF_save_fm DFF_W5114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R028));
DFF_save_fm DFF_W5115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R108));
DFF_save_fm DFF_W5116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R118));
DFF_save_fm DFF_W5117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R128));
DFF_save_fm DFF_W5118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R208));
DFF_save_fm DFF_W5119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R218));
DFF_save_fm DFF_W5120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R228));
DFF_save_fm DFF_W5121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R009));
DFF_save_fm DFF_W5122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R019));
DFF_save_fm DFF_W5123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R029));
DFF_save_fm DFF_W5124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R109));
DFF_save_fm DFF_W5125(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R119));
DFF_save_fm DFF_W5126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R129));
DFF_save_fm DFF_W5127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R209));
DFF_save_fm DFF_W5128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R219));
DFF_save_fm DFF_W5129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R229));
DFF_save_fm DFF_W5130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R00A));
DFF_save_fm DFF_W5131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R01A));
DFF_save_fm DFF_W5132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R02A));
DFF_save_fm DFF_W5133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R10A));
DFF_save_fm DFF_W5134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R11A));
DFF_save_fm DFF_W5135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R12A));
DFF_save_fm DFF_W5136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R20A));
DFF_save_fm DFF_W5137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R21A));
DFF_save_fm DFF_W5138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R22A));
DFF_save_fm DFF_W5139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R00B));
DFF_save_fm DFF_W5140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R01B));
DFF_save_fm DFF_W5141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R02B));
DFF_save_fm DFF_W5142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R10B));
DFF_save_fm DFF_W5143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R11B));
DFF_save_fm DFF_W5144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R12B));
DFF_save_fm DFF_W5145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R20B));
DFF_save_fm DFF_W5146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R21B));
DFF_save_fm DFF_W5147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R22B));
DFF_save_fm DFF_W5148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R00C));
DFF_save_fm DFF_W5149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R01C));
DFF_save_fm DFF_W5150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R02C));
DFF_save_fm DFF_W5151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R10C));
DFF_save_fm DFF_W5152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R11C));
DFF_save_fm DFF_W5153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R12C));
DFF_save_fm DFF_W5154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R20C));
DFF_save_fm DFF_W5155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R21C));
DFF_save_fm DFF_W5156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R22C));
DFF_save_fm DFF_W5157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R00D));
DFF_save_fm DFF_W5158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R01D));
DFF_save_fm DFF_W5159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R02D));
DFF_save_fm DFF_W5160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R10D));
DFF_save_fm DFF_W5161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R11D));
DFF_save_fm DFF_W5162(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R12D));
DFF_save_fm DFF_W5163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R20D));
DFF_save_fm DFF_W5164(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R21D));
DFF_save_fm DFF_W5165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R22D));
DFF_save_fm DFF_W5166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R00E));
DFF_save_fm DFF_W5167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R01E));
DFF_save_fm DFF_W5168(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R02E));
DFF_save_fm DFF_W5169(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R10E));
DFF_save_fm DFF_W5170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R11E));
DFF_save_fm DFF_W5171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R12E));
DFF_save_fm DFF_W5172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R20E));
DFF_save_fm DFF_W5173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R21E));
DFF_save_fm DFF_W5174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R22E));
DFF_save_fm DFF_W5175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R00F));
DFF_save_fm DFF_W5176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R01F));
DFF_save_fm DFF_W5177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R02F));
DFF_save_fm DFF_W5178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R10F));
DFF_save_fm DFF_W5179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R11F));
DFF_save_fm DFF_W5180(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R12F));
DFF_save_fm DFF_W5181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R20F));
DFF_save_fm DFF_W5182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3R21F));
DFF_save_fm DFF_W5183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3R22F));
DFF_save_fm DFF_W5184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S000));
DFF_save_fm DFF_W5185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S010));
DFF_save_fm DFF_W5186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S020));
DFF_save_fm DFF_W5187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S100));
DFF_save_fm DFF_W5188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S110));
DFF_save_fm DFF_W5189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S120));
DFF_save_fm DFF_W5190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S200));
DFF_save_fm DFF_W5191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S210));
DFF_save_fm DFF_W5192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S220));
DFF_save_fm DFF_W5193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S001));
DFF_save_fm DFF_W5194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S011));
DFF_save_fm DFF_W5195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S021));
DFF_save_fm DFF_W5196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S101));
DFF_save_fm DFF_W5197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S111));
DFF_save_fm DFF_W5198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S121));
DFF_save_fm DFF_W5199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S201));
DFF_save_fm DFF_W5200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S211));
DFF_save_fm DFF_W5201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S221));
DFF_save_fm DFF_W5202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S002));
DFF_save_fm DFF_W5203(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S012));
DFF_save_fm DFF_W5204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S022));
DFF_save_fm DFF_W5205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S102));
DFF_save_fm DFF_W5206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S112));
DFF_save_fm DFF_W5207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S122));
DFF_save_fm DFF_W5208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S202));
DFF_save_fm DFF_W5209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S212));
DFF_save_fm DFF_W5210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S222));
DFF_save_fm DFF_W5211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S003));
DFF_save_fm DFF_W5212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S013));
DFF_save_fm DFF_W5213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S023));
DFF_save_fm DFF_W5214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S103));
DFF_save_fm DFF_W5215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S113));
DFF_save_fm DFF_W5216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S123));
DFF_save_fm DFF_W5217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S203));
DFF_save_fm DFF_W5218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S213));
DFF_save_fm DFF_W5219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S223));
DFF_save_fm DFF_W5220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S004));
DFF_save_fm DFF_W5221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S014));
DFF_save_fm DFF_W5222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S024));
DFF_save_fm DFF_W5223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S104));
DFF_save_fm DFF_W5224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S114));
DFF_save_fm DFF_W5225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S124));
DFF_save_fm DFF_W5226(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S204));
DFF_save_fm DFF_W5227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S214));
DFF_save_fm DFF_W5228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S224));
DFF_save_fm DFF_W5229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S005));
DFF_save_fm DFF_W5230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S015));
DFF_save_fm DFF_W5231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S025));
DFF_save_fm DFF_W5232(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S105));
DFF_save_fm DFF_W5233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S115));
DFF_save_fm DFF_W5234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S125));
DFF_save_fm DFF_W5235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S205));
DFF_save_fm DFF_W5236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S215));
DFF_save_fm DFF_W5237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S225));
DFF_save_fm DFF_W5238(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S006));
DFF_save_fm DFF_W5239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S016));
DFF_save_fm DFF_W5240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S026));
DFF_save_fm DFF_W5241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S106));
DFF_save_fm DFF_W5242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S116));
DFF_save_fm DFF_W5243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S126));
DFF_save_fm DFF_W5244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S206));
DFF_save_fm DFF_W5245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S216));
DFF_save_fm DFF_W5246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S226));
DFF_save_fm DFF_W5247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S007));
DFF_save_fm DFF_W5248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S017));
DFF_save_fm DFF_W5249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S027));
DFF_save_fm DFF_W5250(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S107));
DFF_save_fm DFF_W5251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S117));
DFF_save_fm DFF_W5252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S127));
DFF_save_fm DFF_W5253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S207));
DFF_save_fm DFF_W5254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S217));
DFF_save_fm DFF_W5255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S227));
DFF_save_fm DFF_W5256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S008));
DFF_save_fm DFF_W5257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S018));
DFF_save_fm DFF_W5258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S028));
DFF_save_fm DFF_W5259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S108));
DFF_save_fm DFF_W5260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S118));
DFF_save_fm DFF_W5261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S128));
DFF_save_fm DFF_W5262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S208));
DFF_save_fm DFF_W5263(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S218));
DFF_save_fm DFF_W5264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S228));
DFF_save_fm DFF_W5265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S009));
DFF_save_fm DFF_W5266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S019));
DFF_save_fm DFF_W5267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S029));
DFF_save_fm DFF_W5268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S109));
DFF_save_fm DFF_W5269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S119));
DFF_save_fm DFF_W5270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S129));
DFF_save_fm DFF_W5271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S209));
DFF_save_fm DFF_W5272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S219));
DFF_save_fm DFF_W5273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S229));
DFF_save_fm DFF_W5274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S00A));
DFF_save_fm DFF_W5275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S01A));
DFF_save_fm DFF_W5276(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S02A));
DFF_save_fm DFF_W5277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S10A));
DFF_save_fm DFF_W5278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S11A));
DFF_save_fm DFF_W5279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S12A));
DFF_save_fm DFF_W5280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S20A));
DFF_save_fm DFF_W5281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S21A));
DFF_save_fm DFF_W5282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S22A));
DFF_save_fm DFF_W5283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S00B));
DFF_save_fm DFF_W5284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S01B));
DFF_save_fm DFF_W5285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S02B));
DFF_save_fm DFF_W5286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S10B));
DFF_save_fm DFF_W5287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S11B));
DFF_save_fm DFF_W5288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S12B));
DFF_save_fm DFF_W5289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S20B));
DFF_save_fm DFF_W5290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S21B));
DFF_save_fm DFF_W5291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S22B));
DFF_save_fm DFF_W5292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S00C));
DFF_save_fm DFF_W5293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S01C));
DFF_save_fm DFF_W5294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S02C));
DFF_save_fm DFF_W5295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S10C));
DFF_save_fm DFF_W5296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S11C));
DFF_save_fm DFF_W5297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S12C));
DFF_save_fm DFF_W5298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S20C));
DFF_save_fm DFF_W5299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S21C));
DFF_save_fm DFF_W5300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S22C));
DFF_save_fm DFF_W5301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S00D));
DFF_save_fm DFF_W5302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S01D));
DFF_save_fm DFF_W5303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S02D));
DFF_save_fm DFF_W5304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S10D));
DFF_save_fm DFF_W5305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S11D));
DFF_save_fm DFF_W5306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S12D));
DFF_save_fm DFF_W5307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S20D));
DFF_save_fm DFF_W5308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S21D));
DFF_save_fm DFF_W5309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S22D));
DFF_save_fm DFF_W5310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S00E));
DFF_save_fm DFF_W5311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S01E));
DFF_save_fm DFF_W5312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S02E));
DFF_save_fm DFF_W5313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S10E));
DFF_save_fm DFF_W5314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S11E));
DFF_save_fm DFF_W5315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S12E));
DFF_save_fm DFF_W5316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S20E));
DFF_save_fm DFF_W5317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S21E));
DFF_save_fm DFF_W5318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S22E));
DFF_save_fm DFF_W5319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S00F));
DFF_save_fm DFF_W5320(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S01F));
DFF_save_fm DFF_W5321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S02F));
DFF_save_fm DFF_W5322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3S10F));
DFF_save_fm DFF_W5323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S11F));
DFF_save_fm DFF_W5324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S12F));
DFF_save_fm DFF_W5325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S20F));
DFF_save_fm DFF_W5326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S21F));
DFF_save_fm DFF_W5327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3S22F));
DFF_save_fm DFF_W5328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T000));
DFF_save_fm DFF_W5329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T010));
DFF_save_fm DFF_W5330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T020));
DFF_save_fm DFF_W5331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T100));
DFF_save_fm DFF_W5332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T110));
DFF_save_fm DFF_W5333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T120));
DFF_save_fm DFF_W5334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T200));
DFF_save_fm DFF_W5335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T210));
DFF_save_fm DFF_W5336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T220));
DFF_save_fm DFF_W5337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T001));
DFF_save_fm DFF_W5338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T011));
DFF_save_fm DFF_W5339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T021));
DFF_save_fm DFF_W5340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T101));
DFF_save_fm DFF_W5341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T111));
DFF_save_fm DFF_W5342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T121));
DFF_save_fm DFF_W5343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T201));
DFF_save_fm DFF_W5344(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T211));
DFF_save_fm DFF_W5345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T221));
DFF_save_fm DFF_W5346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T002));
DFF_save_fm DFF_W5347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T012));
DFF_save_fm DFF_W5348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T022));
DFF_save_fm DFF_W5349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T102));
DFF_save_fm DFF_W5350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T112));
DFF_save_fm DFF_W5351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T122));
DFF_save_fm DFF_W5352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T202));
DFF_save_fm DFF_W5353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T212));
DFF_save_fm DFF_W5354(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T222));
DFF_save_fm DFF_W5355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T003));
DFF_save_fm DFF_W5356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T013));
DFF_save_fm DFF_W5357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T023));
DFF_save_fm DFF_W5358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T103));
DFF_save_fm DFF_W5359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T113));
DFF_save_fm DFF_W5360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T123));
DFF_save_fm DFF_W5361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T203));
DFF_save_fm DFF_W5362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T213));
DFF_save_fm DFF_W5363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T223));
DFF_save_fm DFF_W5364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T004));
DFF_save_fm DFF_W5365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T014));
DFF_save_fm DFF_W5366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T024));
DFF_save_fm DFF_W5367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T104));
DFF_save_fm DFF_W5368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T114));
DFF_save_fm DFF_W5369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T124));
DFF_save_fm DFF_W5370(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T204));
DFF_save_fm DFF_W5371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T214));
DFF_save_fm DFF_W5372(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T224));
DFF_save_fm DFF_W5373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T005));
DFF_save_fm DFF_W5374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T015));
DFF_save_fm DFF_W5375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T025));
DFF_save_fm DFF_W5376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T105));
DFF_save_fm DFF_W5377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T115));
DFF_save_fm DFF_W5378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T125));
DFF_save_fm DFF_W5379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T205));
DFF_save_fm DFF_W5380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T215));
DFF_save_fm DFF_W5381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T225));
DFF_save_fm DFF_W5382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T006));
DFF_save_fm DFF_W5383(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T016));
DFF_save_fm DFF_W5384(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T026));
DFF_save_fm DFF_W5385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T106));
DFF_save_fm DFF_W5386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T116));
DFF_save_fm DFF_W5387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T126));
DFF_save_fm DFF_W5388(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T206));
DFF_save_fm DFF_W5389(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T216));
DFF_save_fm DFF_W5390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T226));
DFF_save_fm DFF_W5391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T007));
DFF_save_fm DFF_W5392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T017));
DFF_save_fm DFF_W5393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T027));
DFF_save_fm DFF_W5394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T107));
DFF_save_fm DFF_W5395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T117));
DFF_save_fm DFF_W5396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T127));
DFF_save_fm DFF_W5397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T207));
DFF_save_fm DFF_W5398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T217));
DFF_save_fm DFF_W5399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T227));
DFF_save_fm DFF_W5400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T008));
DFF_save_fm DFF_W5401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T018));
DFF_save_fm DFF_W5402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T028));
DFF_save_fm DFF_W5403(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T108));
DFF_save_fm DFF_W5404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T118));
DFF_save_fm DFF_W5405(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T128));
DFF_save_fm DFF_W5406(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T208));
DFF_save_fm DFF_W5407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T218));
DFF_save_fm DFF_W5408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T228));
DFF_save_fm DFF_W5409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T009));
DFF_save_fm DFF_W5410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T019));
DFF_save_fm DFF_W5411(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T029));
DFF_save_fm DFF_W5412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T109));
DFF_save_fm DFF_W5413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T119));
DFF_save_fm DFF_W5414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T129));
DFF_save_fm DFF_W5415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T209));
DFF_save_fm DFF_W5416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T219));
DFF_save_fm DFF_W5417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T229));
DFF_save_fm DFF_W5418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T00A));
DFF_save_fm DFF_W5419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T01A));
DFF_save_fm DFF_W5420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T02A));
DFF_save_fm DFF_W5421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T10A));
DFF_save_fm DFF_W5422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T11A));
DFF_save_fm DFF_W5423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T12A));
DFF_save_fm DFF_W5424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T20A));
DFF_save_fm DFF_W5425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T21A));
DFF_save_fm DFF_W5426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T22A));
DFF_save_fm DFF_W5427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T00B));
DFF_save_fm DFF_W5428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T01B));
DFF_save_fm DFF_W5429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T02B));
DFF_save_fm DFF_W5430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T10B));
DFF_save_fm DFF_W5431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T11B));
DFF_save_fm DFF_W5432(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T12B));
DFF_save_fm DFF_W5433(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T20B));
DFF_save_fm DFF_W5434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T21B));
DFF_save_fm DFF_W5435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T22B));
DFF_save_fm DFF_W5436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T00C));
DFF_save_fm DFF_W5437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T01C));
DFF_save_fm DFF_W5438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T02C));
DFF_save_fm DFF_W5439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T10C));
DFF_save_fm DFF_W5440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T11C));
DFF_save_fm DFF_W5441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T12C));
DFF_save_fm DFF_W5442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T20C));
DFF_save_fm DFF_W5443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T21C));
DFF_save_fm DFF_W5444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T22C));
DFF_save_fm DFF_W5445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T00D));
DFF_save_fm DFF_W5446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T01D));
DFF_save_fm DFF_W5447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T02D));
DFF_save_fm DFF_W5448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T10D));
DFF_save_fm DFF_W5449(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T11D));
DFF_save_fm DFF_W5450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T12D));
DFF_save_fm DFF_W5451(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T20D));
DFF_save_fm DFF_W5452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T21D));
DFF_save_fm DFF_W5453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T22D));
DFF_save_fm DFF_W5454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T00E));
DFF_save_fm DFF_W5455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T01E));
DFF_save_fm DFF_W5456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T02E));
DFF_save_fm DFF_W5457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T10E));
DFF_save_fm DFF_W5458(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T11E));
DFF_save_fm DFF_W5459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T12E));
DFF_save_fm DFF_W5460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T20E));
DFF_save_fm DFF_W5461(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T21E));
DFF_save_fm DFF_W5462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T22E));
DFF_save_fm DFF_W5463(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T00F));
DFF_save_fm DFF_W5464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T01F));
DFF_save_fm DFF_W5465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T02F));
DFF_save_fm DFF_W5466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T10F));
DFF_save_fm DFF_W5467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T11F));
DFF_save_fm DFF_W5468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T12F));
DFF_save_fm DFF_W5469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T20F));
DFF_save_fm DFF_W5470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3T21F));
DFF_save_fm DFF_W5471(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3T22F));
DFF_save_fm DFF_W5472(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U000));
DFF_save_fm DFF_W5473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U010));
DFF_save_fm DFF_W5474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U020));
DFF_save_fm DFF_W5475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U100));
DFF_save_fm DFF_W5476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U110));
DFF_save_fm DFF_W5477(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U120));
DFF_save_fm DFF_W5478(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U200));
DFF_save_fm DFF_W5479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U210));
DFF_save_fm DFF_W5480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U220));
DFF_save_fm DFF_W5481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U001));
DFF_save_fm DFF_W5482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U011));
DFF_save_fm DFF_W5483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U021));
DFF_save_fm DFF_W5484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U101));
DFF_save_fm DFF_W5485(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U111));
DFF_save_fm DFF_W5486(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U121));
DFF_save_fm DFF_W5487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U201));
DFF_save_fm DFF_W5488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U211));
DFF_save_fm DFF_W5489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U221));
DFF_save_fm DFF_W5490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U002));
DFF_save_fm DFF_W5491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U012));
DFF_save_fm DFF_W5492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U022));
DFF_save_fm DFF_W5493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U102));
DFF_save_fm DFF_W5494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U112));
DFF_save_fm DFF_W5495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U122));
DFF_save_fm DFF_W5496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U202));
DFF_save_fm DFF_W5497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U212));
DFF_save_fm DFF_W5498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U222));
DFF_save_fm DFF_W5499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U003));
DFF_save_fm DFF_W5500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U013));
DFF_save_fm DFF_W5501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U023));
DFF_save_fm DFF_W5502(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U103));
DFF_save_fm DFF_W5503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U113));
DFF_save_fm DFF_W5504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U123));
DFF_save_fm DFF_W5505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U203));
DFF_save_fm DFF_W5506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U213));
DFF_save_fm DFF_W5507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U223));
DFF_save_fm DFF_W5508(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U004));
DFF_save_fm DFF_W5509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U014));
DFF_save_fm DFF_W5510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U024));
DFF_save_fm DFF_W5511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U104));
DFF_save_fm DFF_W5512(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U114));
DFF_save_fm DFF_W5513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U124));
DFF_save_fm DFF_W5514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U204));
DFF_save_fm DFF_W5515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U214));
DFF_save_fm DFF_W5516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U224));
DFF_save_fm DFF_W5517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U005));
DFF_save_fm DFF_W5518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U015));
DFF_save_fm DFF_W5519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U025));
DFF_save_fm DFF_W5520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U105));
DFF_save_fm DFF_W5521(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U115));
DFF_save_fm DFF_W5522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U125));
DFF_save_fm DFF_W5523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U205));
DFF_save_fm DFF_W5524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U215));
DFF_save_fm DFF_W5525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U225));
DFF_save_fm DFF_W5526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U006));
DFF_save_fm DFF_W5527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U016));
DFF_save_fm DFF_W5528(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U026));
DFF_save_fm DFF_W5529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U106));
DFF_save_fm DFF_W5530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U116));
DFF_save_fm DFF_W5531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U126));
DFF_save_fm DFF_W5532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U206));
DFF_save_fm DFF_W5533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U216));
DFF_save_fm DFF_W5534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U226));
DFF_save_fm DFF_W5535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U007));
DFF_save_fm DFF_W5536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U017));
DFF_save_fm DFF_W5537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U027));
DFF_save_fm DFF_W5538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U107));
DFF_save_fm DFF_W5539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U117));
DFF_save_fm DFF_W5540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U127));
DFF_save_fm DFF_W5541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U207));
DFF_save_fm DFF_W5542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U217));
DFF_save_fm DFF_W5543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U227));
DFF_save_fm DFF_W5544(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U008));
DFF_save_fm DFF_W5545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U018));
DFF_save_fm DFF_W5546(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U028));
DFF_save_fm DFF_W5547(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U108));
DFF_save_fm DFF_W5548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U118));
DFF_save_fm DFF_W5549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U128));
DFF_save_fm DFF_W5550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U208));
DFF_save_fm DFF_W5551(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U218));
DFF_save_fm DFF_W5552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U228));
DFF_save_fm DFF_W5553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U009));
DFF_save_fm DFF_W5554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U019));
DFF_save_fm DFF_W5555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U029));
DFF_save_fm DFF_W5556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U109));
DFF_save_fm DFF_W5557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U119));
DFF_save_fm DFF_W5558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U129));
DFF_save_fm DFF_W5559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U209));
DFF_save_fm DFF_W5560(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U219));
DFF_save_fm DFF_W5561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U229));
DFF_save_fm DFF_W5562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U00A));
DFF_save_fm DFF_W5563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U01A));
DFF_save_fm DFF_W5564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U02A));
DFF_save_fm DFF_W5565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U10A));
DFF_save_fm DFF_W5566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U11A));
DFF_save_fm DFF_W5567(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U12A));
DFF_save_fm DFF_W5568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U20A));
DFF_save_fm DFF_W5569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U21A));
DFF_save_fm DFF_W5570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U22A));
DFF_save_fm DFF_W5571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U00B));
DFF_save_fm DFF_W5572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U01B));
DFF_save_fm DFF_W5573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U02B));
DFF_save_fm DFF_W5574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U10B));
DFF_save_fm DFF_W5575(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U11B));
DFF_save_fm DFF_W5576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U12B));
DFF_save_fm DFF_W5577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U20B));
DFF_save_fm DFF_W5578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U21B));
DFF_save_fm DFF_W5579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U22B));
DFF_save_fm DFF_W5580(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U00C));
DFF_save_fm DFF_W5581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U01C));
DFF_save_fm DFF_W5582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U02C));
DFF_save_fm DFF_W5583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U10C));
DFF_save_fm DFF_W5584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U11C));
DFF_save_fm DFF_W5585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U12C));
DFF_save_fm DFF_W5586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U20C));
DFF_save_fm DFF_W5587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U21C));
DFF_save_fm DFF_W5588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U22C));
DFF_save_fm DFF_W5589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U00D));
DFF_save_fm DFF_W5590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U01D));
DFF_save_fm DFF_W5591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U02D));
DFF_save_fm DFF_W5592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U10D));
DFF_save_fm DFF_W5593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U11D));
DFF_save_fm DFF_W5594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U12D));
DFF_save_fm DFF_W5595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U20D));
DFF_save_fm DFF_W5596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U21D));
DFF_save_fm DFF_W5597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U22D));
DFF_save_fm DFF_W5598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U00E));
DFF_save_fm DFF_W5599(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U01E));
DFF_save_fm DFF_W5600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U02E));
DFF_save_fm DFF_W5601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U10E));
DFF_save_fm DFF_W5602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U11E));
DFF_save_fm DFF_W5603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U12E));
DFF_save_fm DFF_W5604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U20E));
DFF_save_fm DFF_W5605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U21E));
DFF_save_fm DFF_W5606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U22E));
DFF_save_fm DFF_W5607(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U00F));
DFF_save_fm DFF_W5608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U01F));
DFF_save_fm DFF_W5609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U02F));
DFF_save_fm DFF_W5610(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U10F));
DFF_save_fm DFF_W5611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U11F));
DFF_save_fm DFF_W5612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U12F));
DFF_save_fm DFF_W5613(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U20F));
DFF_save_fm DFF_W5614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3U21F));
DFF_save_fm DFF_W5615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3U22F));
DFF_save_fm DFF_W5616(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V000));
DFF_save_fm DFF_W5617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V010));
DFF_save_fm DFF_W5618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V020));
DFF_save_fm DFF_W5619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V100));
DFF_save_fm DFF_W5620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V110));
DFF_save_fm DFF_W5621(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V120));
DFF_save_fm DFF_W5622(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V200));
DFF_save_fm DFF_W5623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V210));
DFF_save_fm DFF_W5624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V220));
DFF_save_fm DFF_W5625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V001));
DFF_save_fm DFF_W5626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V011));
DFF_save_fm DFF_W5627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V021));
DFF_save_fm DFF_W5628(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V101));
DFF_save_fm DFF_W5629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V111));
DFF_save_fm DFF_W5630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V121));
DFF_save_fm DFF_W5631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V201));
DFF_save_fm DFF_W5632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V211));
DFF_save_fm DFF_W5633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V221));
DFF_save_fm DFF_W5634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V002));
DFF_save_fm DFF_W5635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V012));
DFF_save_fm DFF_W5636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V022));
DFF_save_fm DFF_W5637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V102));
DFF_save_fm DFF_W5638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V112));
DFF_save_fm DFF_W5639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V122));
DFF_save_fm DFF_W5640(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V202));
DFF_save_fm DFF_W5641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V212));
DFF_save_fm DFF_W5642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V222));
DFF_save_fm DFF_W5643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V003));
DFF_save_fm DFF_W5644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V013));
DFF_save_fm DFF_W5645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V023));
DFF_save_fm DFF_W5646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V103));
DFF_save_fm DFF_W5647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V113));
DFF_save_fm DFF_W5648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V123));
DFF_save_fm DFF_W5649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V203));
DFF_save_fm DFF_W5650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V213));
DFF_save_fm DFF_W5651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V223));
DFF_save_fm DFF_W5652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V004));
DFF_save_fm DFF_W5653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V014));
DFF_save_fm DFF_W5654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V024));
DFF_save_fm DFF_W5655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V104));
DFF_save_fm DFF_W5656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V114));
DFF_save_fm DFF_W5657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V124));
DFF_save_fm DFF_W5658(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V204));
DFF_save_fm DFF_W5659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V214));
DFF_save_fm DFF_W5660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V224));
DFF_save_fm DFF_W5661(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V005));
DFF_save_fm DFF_W5662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V015));
DFF_save_fm DFF_W5663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V025));
DFF_save_fm DFF_W5664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V105));
DFF_save_fm DFF_W5665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V115));
DFF_save_fm DFF_W5666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V125));
DFF_save_fm DFF_W5667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V205));
DFF_save_fm DFF_W5668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V215));
DFF_save_fm DFF_W5669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V225));
DFF_save_fm DFF_W5670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V006));
DFF_save_fm DFF_W5671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V016));
DFF_save_fm DFF_W5672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V026));
DFF_save_fm DFF_W5673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V106));
DFF_save_fm DFF_W5674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V116));
DFF_save_fm DFF_W5675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V126));
DFF_save_fm DFF_W5676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V206));
DFF_save_fm DFF_W5677(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V216));
DFF_save_fm DFF_W5678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V226));
DFF_save_fm DFF_W5679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V007));
DFF_save_fm DFF_W5680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V017));
DFF_save_fm DFF_W5681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V027));
DFF_save_fm DFF_W5682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V107));
DFF_save_fm DFF_W5683(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V117));
DFF_save_fm DFF_W5684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V127));
DFF_save_fm DFF_W5685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V207));
DFF_save_fm DFF_W5686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V217));
DFF_save_fm DFF_W5687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V227));
DFF_save_fm DFF_W5688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V008));
DFF_save_fm DFF_W5689(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V018));
DFF_save_fm DFF_W5690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V028));
DFF_save_fm DFF_W5691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V108));
DFF_save_fm DFF_W5692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V118));
DFF_save_fm DFF_W5693(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V128));
DFF_save_fm DFF_W5694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V208));
DFF_save_fm DFF_W5695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V218));
DFF_save_fm DFF_W5696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V228));
DFF_save_fm DFF_W5697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V009));
DFF_save_fm DFF_W5698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V019));
DFF_save_fm DFF_W5699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V029));
DFF_save_fm DFF_W5700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V109));
DFF_save_fm DFF_W5701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V119));
DFF_save_fm DFF_W5702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V129));
DFF_save_fm DFF_W5703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V209));
DFF_save_fm DFF_W5704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V219));
DFF_save_fm DFF_W5705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V229));
DFF_save_fm DFF_W5706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V00A));
DFF_save_fm DFF_W5707(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V01A));
DFF_save_fm DFF_W5708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V02A));
DFF_save_fm DFF_W5709(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V10A));
DFF_save_fm DFF_W5710(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V11A));
DFF_save_fm DFF_W5711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V12A));
DFF_save_fm DFF_W5712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V20A));
DFF_save_fm DFF_W5713(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V21A));
DFF_save_fm DFF_W5714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V22A));
DFF_save_fm DFF_W5715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V00B));
DFF_save_fm DFF_W5716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V01B));
DFF_save_fm DFF_W5717(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V02B));
DFF_save_fm DFF_W5718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V10B));
DFF_save_fm DFF_W5719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V11B));
DFF_save_fm DFF_W5720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V12B));
DFF_save_fm DFF_W5721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V20B));
DFF_save_fm DFF_W5722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V21B));
DFF_save_fm DFF_W5723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V22B));
DFF_save_fm DFF_W5724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V00C));
DFF_save_fm DFF_W5725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V01C));
DFF_save_fm DFF_W5726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V02C));
DFF_save_fm DFF_W5727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V10C));
DFF_save_fm DFF_W5728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V11C));
DFF_save_fm DFF_W5729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V12C));
DFF_save_fm DFF_W5730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V20C));
DFF_save_fm DFF_W5731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V21C));
DFF_save_fm DFF_W5732(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V22C));
DFF_save_fm DFF_W5733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V00D));
DFF_save_fm DFF_W5734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V01D));
DFF_save_fm DFF_W5735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V02D));
DFF_save_fm DFF_W5736(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V10D));
DFF_save_fm DFF_W5737(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V11D));
DFF_save_fm DFF_W5738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V12D));
DFF_save_fm DFF_W5739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V20D));
DFF_save_fm DFF_W5740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V21D));
DFF_save_fm DFF_W5741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V22D));
DFF_save_fm DFF_W5742(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V00E));
DFF_save_fm DFF_W5743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V01E));
DFF_save_fm DFF_W5744(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V02E));
DFF_save_fm DFF_W5745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V10E));
DFF_save_fm DFF_W5746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V11E));
DFF_save_fm DFF_W5747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V12E));
DFF_save_fm DFF_W5748(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V20E));
DFF_save_fm DFF_W5749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V21E));
DFF_save_fm DFF_W5750(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V22E));
DFF_save_fm DFF_W5751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V00F));
DFF_save_fm DFF_W5752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V01F));
DFF_save_fm DFF_W5753(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V02F));
DFF_save_fm DFF_W5754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V10F));
DFF_save_fm DFF_W5755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V11F));
DFF_save_fm DFF_W5756(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V12F));
DFF_save_fm DFF_W5757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V20F));
DFF_save_fm DFF_W5758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3V21F));
DFF_save_fm DFF_W5759(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3V22F));
ninexnine_unit ninexnine_unit_3200(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30000)
);

ninexnine_unit ninexnine_unit_3201(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31000)
);

ninexnine_unit ninexnine_unit_3202(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32000)
);

ninexnine_unit ninexnine_unit_3203(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33000)
);

ninexnine_unit ninexnine_unit_3204(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34000)
);

ninexnine_unit ninexnine_unit_3205(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35000)
);

ninexnine_unit ninexnine_unit_3206(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36000)
);

ninexnine_unit ninexnine_unit_3207(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37000)
);

ninexnine_unit ninexnine_unit_3208(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38000)
);

ninexnine_unit ninexnine_unit_3209(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39000)
);

ninexnine_unit ninexnine_unit_3210(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A000)
);

ninexnine_unit ninexnine_unit_3211(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B000)
);

ninexnine_unit ninexnine_unit_3212(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C000)
);

ninexnine_unit ninexnine_unit_3213(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D000)
);

ninexnine_unit ninexnine_unit_3214(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E000)
);

ninexnine_unit ninexnine_unit_3215(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F000)
);

assign C3000=c30000+c31000+c32000+c33000+c34000+c35000+c36000+c37000+c38000+c39000+c3A000+c3B000+c3C000+c3D000+c3E000+c3F000;
assign A3000=(C3000>=0)?1:0;

assign P4000=A3000;

ninexnine_unit ninexnine_unit_3216(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30010)
);

ninexnine_unit ninexnine_unit_3217(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31010)
);

ninexnine_unit ninexnine_unit_3218(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32010)
);

ninexnine_unit ninexnine_unit_3219(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33010)
);

ninexnine_unit ninexnine_unit_3220(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34010)
);

ninexnine_unit ninexnine_unit_3221(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35010)
);

ninexnine_unit ninexnine_unit_3222(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36010)
);

ninexnine_unit ninexnine_unit_3223(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37010)
);

ninexnine_unit ninexnine_unit_3224(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38010)
);

ninexnine_unit ninexnine_unit_3225(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39010)
);

ninexnine_unit ninexnine_unit_3226(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A010)
);

ninexnine_unit ninexnine_unit_3227(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B010)
);

ninexnine_unit ninexnine_unit_3228(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C010)
);

ninexnine_unit ninexnine_unit_3229(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D010)
);

ninexnine_unit ninexnine_unit_3230(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E010)
);

ninexnine_unit ninexnine_unit_3231(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F010)
);

assign C3010=c30010+c31010+c32010+c33010+c34010+c35010+c36010+c37010+c38010+c39010+c3A010+c3B010+c3C010+c3D010+c3E010+c3F010;
assign A3010=(C3010>=0)?1:0;

assign P4010=A3010;

ninexnine_unit ninexnine_unit_3232(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30020)
);

ninexnine_unit ninexnine_unit_3233(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31020)
);

ninexnine_unit ninexnine_unit_3234(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32020)
);

ninexnine_unit ninexnine_unit_3235(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33020)
);

ninexnine_unit ninexnine_unit_3236(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34020)
);

ninexnine_unit ninexnine_unit_3237(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35020)
);

ninexnine_unit ninexnine_unit_3238(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36020)
);

ninexnine_unit ninexnine_unit_3239(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37020)
);

ninexnine_unit ninexnine_unit_3240(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38020)
);

ninexnine_unit ninexnine_unit_3241(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39020)
);

ninexnine_unit ninexnine_unit_3242(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A020)
);

ninexnine_unit ninexnine_unit_3243(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B020)
);

ninexnine_unit ninexnine_unit_3244(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C020)
);

ninexnine_unit ninexnine_unit_3245(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D020)
);

ninexnine_unit ninexnine_unit_3246(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E020)
);

ninexnine_unit ninexnine_unit_3247(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F020)
);

assign C3020=c30020+c31020+c32020+c33020+c34020+c35020+c36020+c37020+c38020+c39020+c3A020+c3B020+c3C020+c3D020+c3E020+c3F020;
assign A3020=(C3020>=0)?1:0;

assign P4020=A3020;

ninexnine_unit ninexnine_unit_3248(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30100)
);

ninexnine_unit ninexnine_unit_3249(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31100)
);

ninexnine_unit ninexnine_unit_3250(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32100)
);

ninexnine_unit ninexnine_unit_3251(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33100)
);

ninexnine_unit ninexnine_unit_3252(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34100)
);

ninexnine_unit ninexnine_unit_3253(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35100)
);

ninexnine_unit ninexnine_unit_3254(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36100)
);

ninexnine_unit ninexnine_unit_3255(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37100)
);

ninexnine_unit ninexnine_unit_3256(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38100)
);

ninexnine_unit ninexnine_unit_3257(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39100)
);

ninexnine_unit ninexnine_unit_3258(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A100)
);

ninexnine_unit ninexnine_unit_3259(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B100)
);

ninexnine_unit ninexnine_unit_3260(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C100)
);

ninexnine_unit ninexnine_unit_3261(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D100)
);

ninexnine_unit ninexnine_unit_3262(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E100)
);

ninexnine_unit ninexnine_unit_3263(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F100)
);

assign C3100=c30100+c31100+c32100+c33100+c34100+c35100+c36100+c37100+c38100+c39100+c3A100+c3B100+c3C100+c3D100+c3E100+c3F100;
assign A3100=(C3100>=0)?1:0;

assign P4100=A3100;

ninexnine_unit ninexnine_unit_3264(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30110)
);

ninexnine_unit ninexnine_unit_3265(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31110)
);

ninexnine_unit ninexnine_unit_3266(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32110)
);

ninexnine_unit ninexnine_unit_3267(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33110)
);

ninexnine_unit ninexnine_unit_3268(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34110)
);

ninexnine_unit ninexnine_unit_3269(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35110)
);

ninexnine_unit ninexnine_unit_3270(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36110)
);

ninexnine_unit ninexnine_unit_3271(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37110)
);

ninexnine_unit ninexnine_unit_3272(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38110)
);

ninexnine_unit ninexnine_unit_3273(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39110)
);

ninexnine_unit ninexnine_unit_3274(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A110)
);

ninexnine_unit ninexnine_unit_3275(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B110)
);

ninexnine_unit ninexnine_unit_3276(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C110)
);

ninexnine_unit ninexnine_unit_3277(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D110)
);

ninexnine_unit ninexnine_unit_3278(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E110)
);

ninexnine_unit ninexnine_unit_3279(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F110)
);

assign C3110=c30110+c31110+c32110+c33110+c34110+c35110+c36110+c37110+c38110+c39110+c3A110+c3B110+c3C110+c3D110+c3E110+c3F110;
assign A3110=(C3110>=0)?1:0;

assign P4110=A3110;

ninexnine_unit ninexnine_unit_3280(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30120)
);

ninexnine_unit ninexnine_unit_3281(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31120)
);

ninexnine_unit ninexnine_unit_3282(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32120)
);

ninexnine_unit ninexnine_unit_3283(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33120)
);

ninexnine_unit ninexnine_unit_3284(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34120)
);

ninexnine_unit ninexnine_unit_3285(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35120)
);

ninexnine_unit ninexnine_unit_3286(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36120)
);

ninexnine_unit ninexnine_unit_3287(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37120)
);

ninexnine_unit ninexnine_unit_3288(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38120)
);

ninexnine_unit ninexnine_unit_3289(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39120)
);

ninexnine_unit ninexnine_unit_3290(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A120)
);

ninexnine_unit ninexnine_unit_3291(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B120)
);

ninexnine_unit ninexnine_unit_3292(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C120)
);

ninexnine_unit ninexnine_unit_3293(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D120)
);

ninexnine_unit ninexnine_unit_3294(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E120)
);

ninexnine_unit ninexnine_unit_3295(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F120)
);

assign C3120=c30120+c31120+c32120+c33120+c34120+c35120+c36120+c37120+c38120+c39120+c3A120+c3B120+c3C120+c3D120+c3E120+c3F120;
assign A3120=(C3120>=0)?1:0;

assign P4120=A3120;

ninexnine_unit ninexnine_unit_3296(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30200)
);

ninexnine_unit ninexnine_unit_3297(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31200)
);

ninexnine_unit ninexnine_unit_3298(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32200)
);

ninexnine_unit ninexnine_unit_3299(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33200)
);

ninexnine_unit ninexnine_unit_3300(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34200)
);

ninexnine_unit ninexnine_unit_3301(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35200)
);

ninexnine_unit ninexnine_unit_3302(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36200)
);

ninexnine_unit ninexnine_unit_3303(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37200)
);

ninexnine_unit ninexnine_unit_3304(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38200)
);

ninexnine_unit ninexnine_unit_3305(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39200)
);

ninexnine_unit ninexnine_unit_3306(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A200)
);

ninexnine_unit ninexnine_unit_3307(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B200)
);

ninexnine_unit ninexnine_unit_3308(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C200)
);

ninexnine_unit ninexnine_unit_3309(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D200)
);

ninexnine_unit ninexnine_unit_3310(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E200)
);

ninexnine_unit ninexnine_unit_3311(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F200)
);

assign C3200=c30200+c31200+c32200+c33200+c34200+c35200+c36200+c37200+c38200+c39200+c3A200+c3B200+c3C200+c3D200+c3E200+c3F200;
assign A3200=(C3200>=0)?1:0;

assign P4200=A3200;

ninexnine_unit ninexnine_unit_3312(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30210)
);

ninexnine_unit ninexnine_unit_3313(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31210)
);

ninexnine_unit ninexnine_unit_3314(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32210)
);

ninexnine_unit ninexnine_unit_3315(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33210)
);

ninexnine_unit ninexnine_unit_3316(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34210)
);

ninexnine_unit ninexnine_unit_3317(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35210)
);

ninexnine_unit ninexnine_unit_3318(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36210)
);

ninexnine_unit ninexnine_unit_3319(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37210)
);

ninexnine_unit ninexnine_unit_3320(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38210)
);

ninexnine_unit ninexnine_unit_3321(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39210)
);

ninexnine_unit ninexnine_unit_3322(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A210)
);

ninexnine_unit ninexnine_unit_3323(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B210)
);

ninexnine_unit ninexnine_unit_3324(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C210)
);

ninexnine_unit ninexnine_unit_3325(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D210)
);

ninexnine_unit ninexnine_unit_3326(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E210)
);

ninexnine_unit ninexnine_unit_3327(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F210)
);

assign C3210=c30210+c31210+c32210+c33210+c34210+c35210+c36210+c37210+c38210+c39210+c3A210+c3B210+c3C210+c3D210+c3E210+c3F210;
assign A3210=(C3210>=0)?1:0;

assign P4210=A3210;

ninexnine_unit ninexnine_unit_3328(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30220)
);

ninexnine_unit ninexnine_unit_3329(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31220)
);

ninexnine_unit ninexnine_unit_3330(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32220)
);

ninexnine_unit ninexnine_unit_3331(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33220)
);

ninexnine_unit ninexnine_unit_3332(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34220)
);

ninexnine_unit ninexnine_unit_3333(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35220)
);

ninexnine_unit ninexnine_unit_3334(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36220)
);

ninexnine_unit ninexnine_unit_3335(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37220)
);

ninexnine_unit ninexnine_unit_3336(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38220)
);

ninexnine_unit ninexnine_unit_3337(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39220)
);

ninexnine_unit ninexnine_unit_3338(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A220)
);

ninexnine_unit ninexnine_unit_3339(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B220)
);

ninexnine_unit ninexnine_unit_3340(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C220)
);

ninexnine_unit ninexnine_unit_3341(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D220)
);

ninexnine_unit ninexnine_unit_3342(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E220)
);

ninexnine_unit ninexnine_unit_3343(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F220)
);

assign C3220=c30220+c31220+c32220+c33220+c34220+c35220+c36220+c37220+c38220+c39220+c3A220+c3B220+c3C220+c3D220+c3E220+c3F220;
assign A3220=(C3220>=0)?1:0;

assign P4220=A3220;

ninexnine_unit ninexnine_unit_3344(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30001)
);

ninexnine_unit ninexnine_unit_3345(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31001)
);

ninexnine_unit ninexnine_unit_3346(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32001)
);

ninexnine_unit ninexnine_unit_3347(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33001)
);

ninexnine_unit ninexnine_unit_3348(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34001)
);

ninexnine_unit ninexnine_unit_3349(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35001)
);

ninexnine_unit ninexnine_unit_3350(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36001)
);

ninexnine_unit ninexnine_unit_3351(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37001)
);

ninexnine_unit ninexnine_unit_3352(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38001)
);

ninexnine_unit ninexnine_unit_3353(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39001)
);

ninexnine_unit ninexnine_unit_3354(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A001)
);

ninexnine_unit ninexnine_unit_3355(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B001)
);

ninexnine_unit ninexnine_unit_3356(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C001)
);

ninexnine_unit ninexnine_unit_3357(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D001)
);

ninexnine_unit ninexnine_unit_3358(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E001)
);

ninexnine_unit ninexnine_unit_3359(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F001)
);

assign C3001=c30001+c31001+c32001+c33001+c34001+c35001+c36001+c37001+c38001+c39001+c3A001+c3B001+c3C001+c3D001+c3E001+c3F001;
assign A3001=(C3001>=0)?1:0;

assign P4001=A3001;

ninexnine_unit ninexnine_unit_3360(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30011)
);

ninexnine_unit ninexnine_unit_3361(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31011)
);

ninexnine_unit ninexnine_unit_3362(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32011)
);

ninexnine_unit ninexnine_unit_3363(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33011)
);

ninexnine_unit ninexnine_unit_3364(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34011)
);

ninexnine_unit ninexnine_unit_3365(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35011)
);

ninexnine_unit ninexnine_unit_3366(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36011)
);

ninexnine_unit ninexnine_unit_3367(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37011)
);

ninexnine_unit ninexnine_unit_3368(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38011)
);

ninexnine_unit ninexnine_unit_3369(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39011)
);

ninexnine_unit ninexnine_unit_3370(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A011)
);

ninexnine_unit ninexnine_unit_3371(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B011)
);

ninexnine_unit ninexnine_unit_3372(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C011)
);

ninexnine_unit ninexnine_unit_3373(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D011)
);

ninexnine_unit ninexnine_unit_3374(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E011)
);

ninexnine_unit ninexnine_unit_3375(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F011)
);

assign C3011=c30011+c31011+c32011+c33011+c34011+c35011+c36011+c37011+c38011+c39011+c3A011+c3B011+c3C011+c3D011+c3E011+c3F011;
assign A3011=(C3011>=0)?1:0;

assign P4011=A3011;

ninexnine_unit ninexnine_unit_3376(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30021)
);

ninexnine_unit ninexnine_unit_3377(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31021)
);

ninexnine_unit ninexnine_unit_3378(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32021)
);

ninexnine_unit ninexnine_unit_3379(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33021)
);

ninexnine_unit ninexnine_unit_3380(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34021)
);

ninexnine_unit ninexnine_unit_3381(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35021)
);

ninexnine_unit ninexnine_unit_3382(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36021)
);

ninexnine_unit ninexnine_unit_3383(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37021)
);

ninexnine_unit ninexnine_unit_3384(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38021)
);

ninexnine_unit ninexnine_unit_3385(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39021)
);

ninexnine_unit ninexnine_unit_3386(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A021)
);

ninexnine_unit ninexnine_unit_3387(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B021)
);

ninexnine_unit ninexnine_unit_3388(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C021)
);

ninexnine_unit ninexnine_unit_3389(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D021)
);

ninexnine_unit ninexnine_unit_3390(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E021)
);

ninexnine_unit ninexnine_unit_3391(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F021)
);

assign C3021=c30021+c31021+c32021+c33021+c34021+c35021+c36021+c37021+c38021+c39021+c3A021+c3B021+c3C021+c3D021+c3E021+c3F021;
assign A3021=(C3021>=0)?1:0;

assign P4021=A3021;

ninexnine_unit ninexnine_unit_3392(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30101)
);

ninexnine_unit ninexnine_unit_3393(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31101)
);

ninexnine_unit ninexnine_unit_3394(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32101)
);

ninexnine_unit ninexnine_unit_3395(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33101)
);

ninexnine_unit ninexnine_unit_3396(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34101)
);

ninexnine_unit ninexnine_unit_3397(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35101)
);

ninexnine_unit ninexnine_unit_3398(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36101)
);

ninexnine_unit ninexnine_unit_3399(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37101)
);

ninexnine_unit ninexnine_unit_3400(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38101)
);

ninexnine_unit ninexnine_unit_3401(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39101)
);

ninexnine_unit ninexnine_unit_3402(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A101)
);

ninexnine_unit ninexnine_unit_3403(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B101)
);

ninexnine_unit ninexnine_unit_3404(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C101)
);

ninexnine_unit ninexnine_unit_3405(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D101)
);

ninexnine_unit ninexnine_unit_3406(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E101)
);

ninexnine_unit ninexnine_unit_3407(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F101)
);

assign C3101=c30101+c31101+c32101+c33101+c34101+c35101+c36101+c37101+c38101+c39101+c3A101+c3B101+c3C101+c3D101+c3E101+c3F101;
assign A3101=(C3101>=0)?1:0;

assign P4101=A3101;

ninexnine_unit ninexnine_unit_3408(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30111)
);

ninexnine_unit ninexnine_unit_3409(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31111)
);

ninexnine_unit ninexnine_unit_3410(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32111)
);

ninexnine_unit ninexnine_unit_3411(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33111)
);

ninexnine_unit ninexnine_unit_3412(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34111)
);

ninexnine_unit ninexnine_unit_3413(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35111)
);

ninexnine_unit ninexnine_unit_3414(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36111)
);

ninexnine_unit ninexnine_unit_3415(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37111)
);

ninexnine_unit ninexnine_unit_3416(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38111)
);

ninexnine_unit ninexnine_unit_3417(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39111)
);

ninexnine_unit ninexnine_unit_3418(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A111)
);

ninexnine_unit ninexnine_unit_3419(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B111)
);

ninexnine_unit ninexnine_unit_3420(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C111)
);

ninexnine_unit ninexnine_unit_3421(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D111)
);

ninexnine_unit ninexnine_unit_3422(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E111)
);

ninexnine_unit ninexnine_unit_3423(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F111)
);

assign C3111=c30111+c31111+c32111+c33111+c34111+c35111+c36111+c37111+c38111+c39111+c3A111+c3B111+c3C111+c3D111+c3E111+c3F111;
assign A3111=(C3111>=0)?1:0;

assign P4111=A3111;

ninexnine_unit ninexnine_unit_3424(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30121)
);

ninexnine_unit ninexnine_unit_3425(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31121)
);

ninexnine_unit ninexnine_unit_3426(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32121)
);

ninexnine_unit ninexnine_unit_3427(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33121)
);

ninexnine_unit ninexnine_unit_3428(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34121)
);

ninexnine_unit ninexnine_unit_3429(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35121)
);

ninexnine_unit ninexnine_unit_3430(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36121)
);

ninexnine_unit ninexnine_unit_3431(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37121)
);

ninexnine_unit ninexnine_unit_3432(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38121)
);

ninexnine_unit ninexnine_unit_3433(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39121)
);

ninexnine_unit ninexnine_unit_3434(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A121)
);

ninexnine_unit ninexnine_unit_3435(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B121)
);

ninexnine_unit ninexnine_unit_3436(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C121)
);

ninexnine_unit ninexnine_unit_3437(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D121)
);

ninexnine_unit ninexnine_unit_3438(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E121)
);

ninexnine_unit ninexnine_unit_3439(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F121)
);

assign C3121=c30121+c31121+c32121+c33121+c34121+c35121+c36121+c37121+c38121+c39121+c3A121+c3B121+c3C121+c3D121+c3E121+c3F121;
assign A3121=(C3121>=0)?1:0;

assign P4121=A3121;

ninexnine_unit ninexnine_unit_3440(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30201)
);

ninexnine_unit ninexnine_unit_3441(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31201)
);

ninexnine_unit ninexnine_unit_3442(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32201)
);

ninexnine_unit ninexnine_unit_3443(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33201)
);

ninexnine_unit ninexnine_unit_3444(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34201)
);

ninexnine_unit ninexnine_unit_3445(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35201)
);

ninexnine_unit ninexnine_unit_3446(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36201)
);

ninexnine_unit ninexnine_unit_3447(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37201)
);

ninexnine_unit ninexnine_unit_3448(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38201)
);

ninexnine_unit ninexnine_unit_3449(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39201)
);

ninexnine_unit ninexnine_unit_3450(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A201)
);

ninexnine_unit ninexnine_unit_3451(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B201)
);

ninexnine_unit ninexnine_unit_3452(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C201)
);

ninexnine_unit ninexnine_unit_3453(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D201)
);

ninexnine_unit ninexnine_unit_3454(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E201)
);

ninexnine_unit ninexnine_unit_3455(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F201)
);

assign C3201=c30201+c31201+c32201+c33201+c34201+c35201+c36201+c37201+c38201+c39201+c3A201+c3B201+c3C201+c3D201+c3E201+c3F201;
assign A3201=(C3201>=0)?1:0;

assign P4201=A3201;

ninexnine_unit ninexnine_unit_3456(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30211)
);

ninexnine_unit ninexnine_unit_3457(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31211)
);

ninexnine_unit ninexnine_unit_3458(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32211)
);

ninexnine_unit ninexnine_unit_3459(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33211)
);

ninexnine_unit ninexnine_unit_3460(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34211)
);

ninexnine_unit ninexnine_unit_3461(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35211)
);

ninexnine_unit ninexnine_unit_3462(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36211)
);

ninexnine_unit ninexnine_unit_3463(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37211)
);

ninexnine_unit ninexnine_unit_3464(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38211)
);

ninexnine_unit ninexnine_unit_3465(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39211)
);

ninexnine_unit ninexnine_unit_3466(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A211)
);

ninexnine_unit ninexnine_unit_3467(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B211)
);

ninexnine_unit ninexnine_unit_3468(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C211)
);

ninexnine_unit ninexnine_unit_3469(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D211)
);

ninexnine_unit ninexnine_unit_3470(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E211)
);

ninexnine_unit ninexnine_unit_3471(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F211)
);

assign C3211=c30211+c31211+c32211+c33211+c34211+c35211+c36211+c37211+c38211+c39211+c3A211+c3B211+c3C211+c3D211+c3E211+c3F211;
assign A3211=(C3211>=0)?1:0;

assign P4211=A3211;

ninexnine_unit ninexnine_unit_3472(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30221)
);

ninexnine_unit ninexnine_unit_3473(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31221)
);

ninexnine_unit ninexnine_unit_3474(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32221)
);

ninexnine_unit ninexnine_unit_3475(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33221)
);

ninexnine_unit ninexnine_unit_3476(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34221)
);

ninexnine_unit ninexnine_unit_3477(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35221)
);

ninexnine_unit ninexnine_unit_3478(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36221)
);

ninexnine_unit ninexnine_unit_3479(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37221)
);

ninexnine_unit ninexnine_unit_3480(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38221)
);

ninexnine_unit ninexnine_unit_3481(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39221)
);

ninexnine_unit ninexnine_unit_3482(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A221)
);

ninexnine_unit ninexnine_unit_3483(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B221)
);

ninexnine_unit ninexnine_unit_3484(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C221)
);

ninexnine_unit ninexnine_unit_3485(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D221)
);

ninexnine_unit ninexnine_unit_3486(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E221)
);

ninexnine_unit ninexnine_unit_3487(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F221)
);

assign C3221=c30221+c31221+c32221+c33221+c34221+c35221+c36221+c37221+c38221+c39221+c3A221+c3B221+c3C221+c3D221+c3E221+c3F221;
assign A3221=(C3221>=0)?1:0;

assign P4221=A3221;

ninexnine_unit ninexnine_unit_3488(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30002)
);

ninexnine_unit ninexnine_unit_3489(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31002)
);

ninexnine_unit ninexnine_unit_3490(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32002)
);

ninexnine_unit ninexnine_unit_3491(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33002)
);

ninexnine_unit ninexnine_unit_3492(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34002)
);

ninexnine_unit ninexnine_unit_3493(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35002)
);

ninexnine_unit ninexnine_unit_3494(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36002)
);

ninexnine_unit ninexnine_unit_3495(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37002)
);

ninexnine_unit ninexnine_unit_3496(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38002)
);

ninexnine_unit ninexnine_unit_3497(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39002)
);

ninexnine_unit ninexnine_unit_3498(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A002)
);

ninexnine_unit ninexnine_unit_3499(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B002)
);

ninexnine_unit ninexnine_unit_3500(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C002)
);

ninexnine_unit ninexnine_unit_3501(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D002)
);

ninexnine_unit ninexnine_unit_3502(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E002)
);

ninexnine_unit ninexnine_unit_3503(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F002)
);

assign C3002=c30002+c31002+c32002+c33002+c34002+c35002+c36002+c37002+c38002+c39002+c3A002+c3B002+c3C002+c3D002+c3E002+c3F002;
assign A3002=(C3002>=0)?1:0;

assign P4002=A3002;

ninexnine_unit ninexnine_unit_3504(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30012)
);

ninexnine_unit ninexnine_unit_3505(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31012)
);

ninexnine_unit ninexnine_unit_3506(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32012)
);

ninexnine_unit ninexnine_unit_3507(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33012)
);

ninexnine_unit ninexnine_unit_3508(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34012)
);

ninexnine_unit ninexnine_unit_3509(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35012)
);

ninexnine_unit ninexnine_unit_3510(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36012)
);

ninexnine_unit ninexnine_unit_3511(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37012)
);

ninexnine_unit ninexnine_unit_3512(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38012)
);

ninexnine_unit ninexnine_unit_3513(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39012)
);

ninexnine_unit ninexnine_unit_3514(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A012)
);

ninexnine_unit ninexnine_unit_3515(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B012)
);

ninexnine_unit ninexnine_unit_3516(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C012)
);

ninexnine_unit ninexnine_unit_3517(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D012)
);

ninexnine_unit ninexnine_unit_3518(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E012)
);

ninexnine_unit ninexnine_unit_3519(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F012)
);

assign C3012=c30012+c31012+c32012+c33012+c34012+c35012+c36012+c37012+c38012+c39012+c3A012+c3B012+c3C012+c3D012+c3E012+c3F012;
assign A3012=(C3012>=0)?1:0;

assign P4012=A3012;

ninexnine_unit ninexnine_unit_3520(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30022)
);

ninexnine_unit ninexnine_unit_3521(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31022)
);

ninexnine_unit ninexnine_unit_3522(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32022)
);

ninexnine_unit ninexnine_unit_3523(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33022)
);

ninexnine_unit ninexnine_unit_3524(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34022)
);

ninexnine_unit ninexnine_unit_3525(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35022)
);

ninexnine_unit ninexnine_unit_3526(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36022)
);

ninexnine_unit ninexnine_unit_3527(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37022)
);

ninexnine_unit ninexnine_unit_3528(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38022)
);

ninexnine_unit ninexnine_unit_3529(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39022)
);

ninexnine_unit ninexnine_unit_3530(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A022)
);

ninexnine_unit ninexnine_unit_3531(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B022)
);

ninexnine_unit ninexnine_unit_3532(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C022)
);

ninexnine_unit ninexnine_unit_3533(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D022)
);

ninexnine_unit ninexnine_unit_3534(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E022)
);

ninexnine_unit ninexnine_unit_3535(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F022)
);

assign C3022=c30022+c31022+c32022+c33022+c34022+c35022+c36022+c37022+c38022+c39022+c3A022+c3B022+c3C022+c3D022+c3E022+c3F022;
assign A3022=(C3022>=0)?1:0;

assign P4022=A3022;

ninexnine_unit ninexnine_unit_3536(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30102)
);

ninexnine_unit ninexnine_unit_3537(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31102)
);

ninexnine_unit ninexnine_unit_3538(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32102)
);

ninexnine_unit ninexnine_unit_3539(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33102)
);

ninexnine_unit ninexnine_unit_3540(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34102)
);

ninexnine_unit ninexnine_unit_3541(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35102)
);

ninexnine_unit ninexnine_unit_3542(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36102)
);

ninexnine_unit ninexnine_unit_3543(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37102)
);

ninexnine_unit ninexnine_unit_3544(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38102)
);

ninexnine_unit ninexnine_unit_3545(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39102)
);

ninexnine_unit ninexnine_unit_3546(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A102)
);

ninexnine_unit ninexnine_unit_3547(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B102)
);

ninexnine_unit ninexnine_unit_3548(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C102)
);

ninexnine_unit ninexnine_unit_3549(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D102)
);

ninexnine_unit ninexnine_unit_3550(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E102)
);

ninexnine_unit ninexnine_unit_3551(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F102)
);

assign C3102=c30102+c31102+c32102+c33102+c34102+c35102+c36102+c37102+c38102+c39102+c3A102+c3B102+c3C102+c3D102+c3E102+c3F102;
assign A3102=(C3102>=0)?1:0;

assign P4102=A3102;

ninexnine_unit ninexnine_unit_3552(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30112)
);

ninexnine_unit ninexnine_unit_3553(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31112)
);

ninexnine_unit ninexnine_unit_3554(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32112)
);

ninexnine_unit ninexnine_unit_3555(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33112)
);

ninexnine_unit ninexnine_unit_3556(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34112)
);

ninexnine_unit ninexnine_unit_3557(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35112)
);

ninexnine_unit ninexnine_unit_3558(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36112)
);

ninexnine_unit ninexnine_unit_3559(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37112)
);

ninexnine_unit ninexnine_unit_3560(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38112)
);

ninexnine_unit ninexnine_unit_3561(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39112)
);

ninexnine_unit ninexnine_unit_3562(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A112)
);

ninexnine_unit ninexnine_unit_3563(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B112)
);

ninexnine_unit ninexnine_unit_3564(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C112)
);

ninexnine_unit ninexnine_unit_3565(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D112)
);

ninexnine_unit ninexnine_unit_3566(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E112)
);

ninexnine_unit ninexnine_unit_3567(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F112)
);

assign C3112=c30112+c31112+c32112+c33112+c34112+c35112+c36112+c37112+c38112+c39112+c3A112+c3B112+c3C112+c3D112+c3E112+c3F112;
assign A3112=(C3112>=0)?1:0;

assign P4112=A3112;

ninexnine_unit ninexnine_unit_3568(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30122)
);

ninexnine_unit ninexnine_unit_3569(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31122)
);

ninexnine_unit ninexnine_unit_3570(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32122)
);

ninexnine_unit ninexnine_unit_3571(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33122)
);

ninexnine_unit ninexnine_unit_3572(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34122)
);

ninexnine_unit ninexnine_unit_3573(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35122)
);

ninexnine_unit ninexnine_unit_3574(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36122)
);

ninexnine_unit ninexnine_unit_3575(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37122)
);

ninexnine_unit ninexnine_unit_3576(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38122)
);

ninexnine_unit ninexnine_unit_3577(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39122)
);

ninexnine_unit ninexnine_unit_3578(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A122)
);

ninexnine_unit ninexnine_unit_3579(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B122)
);

ninexnine_unit ninexnine_unit_3580(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C122)
);

ninexnine_unit ninexnine_unit_3581(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D122)
);

ninexnine_unit ninexnine_unit_3582(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E122)
);

ninexnine_unit ninexnine_unit_3583(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F122)
);

assign C3122=c30122+c31122+c32122+c33122+c34122+c35122+c36122+c37122+c38122+c39122+c3A122+c3B122+c3C122+c3D122+c3E122+c3F122;
assign A3122=(C3122>=0)?1:0;

assign P4122=A3122;

ninexnine_unit ninexnine_unit_3584(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30202)
);

ninexnine_unit ninexnine_unit_3585(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31202)
);

ninexnine_unit ninexnine_unit_3586(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32202)
);

ninexnine_unit ninexnine_unit_3587(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33202)
);

ninexnine_unit ninexnine_unit_3588(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34202)
);

ninexnine_unit ninexnine_unit_3589(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35202)
);

ninexnine_unit ninexnine_unit_3590(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36202)
);

ninexnine_unit ninexnine_unit_3591(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37202)
);

ninexnine_unit ninexnine_unit_3592(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38202)
);

ninexnine_unit ninexnine_unit_3593(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39202)
);

ninexnine_unit ninexnine_unit_3594(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A202)
);

ninexnine_unit ninexnine_unit_3595(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B202)
);

ninexnine_unit ninexnine_unit_3596(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C202)
);

ninexnine_unit ninexnine_unit_3597(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D202)
);

ninexnine_unit ninexnine_unit_3598(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E202)
);

ninexnine_unit ninexnine_unit_3599(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F202)
);

assign C3202=c30202+c31202+c32202+c33202+c34202+c35202+c36202+c37202+c38202+c39202+c3A202+c3B202+c3C202+c3D202+c3E202+c3F202;
assign A3202=(C3202>=0)?1:0;

assign P4202=A3202;

ninexnine_unit ninexnine_unit_3600(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30212)
);

ninexnine_unit ninexnine_unit_3601(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31212)
);

ninexnine_unit ninexnine_unit_3602(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32212)
);

ninexnine_unit ninexnine_unit_3603(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33212)
);

ninexnine_unit ninexnine_unit_3604(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34212)
);

ninexnine_unit ninexnine_unit_3605(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35212)
);

ninexnine_unit ninexnine_unit_3606(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36212)
);

ninexnine_unit ninexnine_unit_3607(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37212)
);

ninexnine_unit ninexnine_unit_3608(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38212)
);

ninexnine_unit ninexnine_unit_3609(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39212)
);

ninexnine_unit ninexnine_unit_3610(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A212)
);

ninexnine_unit ninexnine_unit_3611(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B212)
);

ninexnine_unit ninexnine_unit_3612(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C212)
);

ninexnine_unit ninexnine_unit_3613(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D212)
);

ninexnine_unit ninexnine_unit_3614(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E212)
);

ninexnine_unit ninexnine_unit_3615(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F212)
);

assign C3212=c30212+c31212+c32212+c33212+c34212+c35212+c36212+c37212+c38212+c39212+c3A212+c3B212+c3C212+c3D212+c3E212+c3F212;
assign A3212=(C3212>=0)?1:0;

assign P4212=A3212;

ninexnine_unit ninexnine_unit_3616(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W32000),
				.b1(W32010),
				.b2(W32020),
				.b3(W32100),
				.b4(W32110),
				.b5(W32120),
				.b6(W32200),
				.b7(W32210),
				.b8(W32220),
				.c(c30222)
);

ninexnine_unit ninexnine_unit_3617(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W32001),
				.b1(W32011),
				.b2(W32021),
				.b3(W32101),
				.b4(W32111),
				.b5(W32121),
				.b6(W32201),
				.b7(W32211),
				.b8(W32221),
				.c(c31222)
);

ninexnine_unit ninexnine_unit_3618(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W32002),
				.b1(W32012),
				.b2(W32022),
				.b3(W32102),
				.b4(W32112),
				.b5(W32122),
				.b6(W32202),
				.b7(W32212),
				.b8(W32222),
				.c(c32222)
);

ninexnine_unit ninexnine_unit_3619(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W32003),
				.b1(W32013),
				.b2(W32023),
				.b3(W32103),
				.b4(W32113),
				.b5(W32123),
				.b6(W32203),
				.b7(W32213),
				.b8(W32223),
				.c(c33222)
);

ninexnine_unit ninexnine_unit_3620(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W32004),
				.b1(W32014),
				.b2(W32024),
				.b3(W32104),
				.b4(W32114),
				.b5(W32124),
				.b6(W32204),
				.b7(W32214),
				.b8(W32224),
				.c(c34222)
);

ninexnine_unit ninexnine_unit_3621(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W32005),
				.b1(W32015),
				.b2(W32025),
				.b3(W32105),
				.b4(W32115),
				.b5(W32125),
				.b6(W32205),
				.b7(W32215),
				.b8(W32225),
				.c(c35222)
);

ninexnine_unit ninexnine_unit_3622(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W32006),
				.b1(W32016),
				.b2(W32026),
				.b3(W32106),
				.b4(W32116),
				.b5(W32126),
				.b6(W32206),
				.b7(W32216),
				.b8(W32226),
				.c(c36222)
);

ninexnine_unit ninexnine_unit_3623(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W32007),
				.b1(W32017),
				.b2(W32027),
				.b3(W32107),
				.b4(W32117),
				.b5(W32127),
				.b6(W32207),
				.b7(W32217),
				.b8(W32227),
				.c(c37222)
);

ninexnine_unit ninexnine_unit_3624(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W32008),
				.b1(W32018),
				.b2(W32028),
				.b3(W32108),
				.b4(W32118),
				.b5(W32128),
				.b6(W32208),
				.b7(W32218),
				.b8(W32228),
				.c(c38222)
);

ninexnine_unit ninexnine_unit_3625(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W32009),
				.b1(W32019),
				.b2(W32029),
				.b3(W32109),
				.b4(W32119),
				.b5(W32129),
				.b6(W32209),
				.b7(W32219),
				.b8(W32229),
				.c(c39222)
);

ninexnine_unit ninexnine_unit_3626(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3200A),
				.b1(W3201A),
				.b2(W3202A),
				.b3(W3210A),
				.b4(W3211A),
				.b5(W3212A),
				.b6(W3220A),
				.b7(W3221A),
				.b8(W3222A),
				.c(c3A222)
);

ninexnine_unit ninexnine_unit_3627(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3200B),
				.b1(W3201B),
				.b2(W3202B),
				.b3(W3210B),
				.b4(W3211B),
				.b5(W3212B),
				.b6(W3220B),
				.b7(W3221B),
				.b8(W3222B),
				.c(c3B222)
);

ninexnine_unit ninexnine_unit_3628(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3200C),
				.b1(W3201C),
				.b2(W3202C),
				.b3(W3210C),
				.b4(W3211C),
				.b5(W3212C),
				.b6(W3220C),
				.b7(W3221C),
				.b8(W3222C),
				.c(c3C222)
);

ninexnine_unit ninexnine_unit_3629(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3200D),
				.b1(W3201D),
				.b2(W3202D),
				.b3(W3210D),
				.b4(W3211D),
				.b5(W3212D),
				.b6(W3220D),
				.b7(W3221D),
				.b8(W3222D),
				.c(c3D222)
);

ninexnine_unit ninexnine_unit_3630(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3200E),
				.b1(W3201E),
				.b2(W3202E),
				.b3(W3210E),
				.b4(W3211E),
				.b5(W3212E),
				.b6(W3220E),
				.b7(W3221E),
				.b8(W3222E),
				.c(c3E222)
);

ninexnine_unit ninexnine_unit_3631(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3200F),
				.b1(W3201F),
				.b2(W3202F),
				.b3(W3210F),
				.b4(W3211F),
				.b5(W3212F),
				.b6(W3220F),
				.b7(W3221F),
				.b8(W3222F),
				.c(c3F222)
);

assign C3222=c30222+c31222+c32222+c33222+c34222+c35222+c36222+c37222+c38222+c39222+c3A222+c3B222+c3C222+c3D222+c3E222+c3F222;
assign A3222=(C3222>=0)?1:0;

assign P4222=A3222;

ninexnine_unit ninexnine_unit_3632(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30003)
);

ninexnine_unit ninexnine_unit_3633(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31003)
);

ninexnine_unit ninexnine_unit_3634(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32003)
);

ninexnine_unit ninexnine_unit_3635(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33003)
);

ninexnine_unit ninexnine_unit_3636(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34003)
);

ninexnine_unit ninexnine_unit_3637(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35003)
);

ninexnine_unit ninexnine_unit_3638(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36003)
);

ninexnine_unit ninexnine_unit_3639(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37003)
);

ninexnine_unit ninexnine_unit_3640(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38003)
);

ninexnine_unit ninexnine_unit_3641(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39003)
);

ninexnine_unit ninexnine_unit_3642(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A003)
);

ninexnine_unit ninexnine_unit_3643(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B003)
);

ninexnine_unit ninexnine_unit_3644(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C003)
);

ninexnine_unit ninexnine_unit_3645(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D003)
);

ninexnine_unit ninexnine_unit_3646(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E003)
);

ninexnine_unit ninexnine_unit_3647(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F003)
);

assign C3003=c30003+c31003+c32003+c33003+c34003+c35003+c36003+c37003+c38003+c39003+c3A003+c3B003+c3C003+c3D003+c3E003+c3F003;
assign A3003=(C3003>=0)?1:0;

assign P4003=A3003;

ninexnine_unit ninexnine_unit_3648(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30013)
);

ninexnine_unit ninexnine_unit_3649(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31013)
);

ninexnine_unit ninexnine_unit_3650(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32013)
);

ninexnine_unit ninexnine_unit_3651(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33013)
);

ninexnine_unit ninexnine_unit_3652(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34013)
);

ninexnine_unit ninexnine_unit_3653(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35013)
);

ninexnine_unit ninexnine_unit_3654(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36013)
);

ninexnine_unit ninexnine_unit_3655(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37013)
);

ninexnine_unit ninexnine_unit_3656(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38013)
);

ninexnine_unit ninexnine_unit_3657(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39013)
);

ninexnine_unit ninexnine_unit_3658(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A013)
);

ninexnine_unit ninexnine_unit_3659(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B013)
);

ninexnine_unit ninexnine_unit_3660(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C013)
);

ninexnine_unit ninexnine_unit_3661(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D013)
);

ninexnine_unit ninexnine_unit_3662(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E013)
);

ninexnine_unit ninexnine_unit_3663(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F013)
);

assign C3013=c30013+c31013+c32013+c33013+c34013+c35013+c36013+c37013+c38013+c39013+c3A013+c3B013+c3C013+c3D013+c3E013+c3F013;
assign A3013=(C3013>=0)?1:0;

assign P4013=A3013;

ninexnine_unit ninexnine_unit_3664(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30023)
);

ninexnine_unit ninexnine_unit_3665(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31023)
);

ninexnine_unit ninexnine_unit_3666(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32023)
);

ninexnine_unit ninexnine_unit_3667(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33023)
);

ninexnine_unit ninexnine_unit_3668(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34023)
);

ninexnine_unit ninexnine_unit_3669(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35023)
);

ninexnine_unit ninexnine_unit_3670(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36023)
);

ninexnine_unit ninexnine_unit_3671(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37023)
);

ninexnine_unit ninexnine_unit_3672(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38023)
);

ninexnine_unit ninexnine_unit_3673(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39023)
);

ninexnine_unit ninexnine_unit_3674(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A023)
);

ninexnine_unit ninexnine_unit_3675(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B023)
);

ninexnine_unit ninexnine_unit_3676(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C023)
);

ninexnine_unit ninexnine_unit_3677(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D023)
);

ninexnine_unit ninexnine_unit_3678(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E023)
);

ninexnine_unit ninexnine_unit_3679(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F023)
);

assign C3023=c30023+c31023+c32023+c33023+c34023+c35023+c36023+c37023+c38023+c39023+c3A023+c3B023+c3C023+c3D023+c3E023+c3F023;
assign A3023=(C3023>=0)?1:0;

assign P4023=A3023;

ninexnine_unit ninexnine_unit_3680(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30103)
);

ninexnine_unit ninexnine_unit_3681(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31103)
);

ninexnine_unit ninexnine_unit_3682(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32103)
);

ninexnine_unit ninexnine_unit_3683(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33103)
);

ninexnine_unit ninexnine_unit_3684(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34103)
);

ninexnine_unit ninexnine_unit_3685(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35103)
);

ninexnine_unit ninexnine_unit_3686(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36103)
);

ninexnine_unit ninexnine_unit_3687(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37103)
);

ninexnine_unit ninexnine_unit_3688(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38103)
);

ninexnine_unit ninexnine_unit_3689(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39103)
);

ninexnine_unit ninexnine_unit_3690(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A103)
);

ninexnine_unit ninexnine_unit_3691(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B103)
);

ninexnine_unit ninexnine_unit_3692(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C103)
);

ninexnine_unit ninexnine_unit_3693(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D103)
);

ninexnine_unit ninexnine_unit_3694(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E103)
);

ninexnine_unit ninexnine_unit_3695(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F103)
);

assign C3103=c30103+c31103+c32103+c33103+c34103+c35103+c36103+c37103+c38103+c39103+c3A103+c3B103+c3C103+c3D103+c3E103+c3F103;
assign A3103=(C3103>=0)?1:0;

assign P4103=A3103;

ninexnine_unit ninexnine_unit_3696(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30113)
);

ninexnine_unit ninexnine_unit_3697(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31113)
);

ninexnine_unit ninexnine_unit_3698(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32113)
);

ninexnine_unit ninexnine_unit_3699(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33113)
);

ninexnine_unit ninexnine_unit_3700(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34113)
);

ninexnine_unit ninexnine_unit_3701(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35113)
);

ninexnine_unit ninexnine_unit_3702(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36113)
);

ninexnine_unit ninexnine_unit_3703(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37113)
);

ninexnine_unit ninexnine_unit_3704(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38113)
);

ninexnine_unit ninexnine_unit_3705(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39113)
);

ninexnine_unit ninexnine_unit_3706(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A113)
);

ninexnine_unit ninexnine_unit_3707(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B113)
);

ninexnine_unit ninexnine_unit_3708(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C113)
);

ninexnine_unit ninexnine_unit_3709(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D113)
);

ninexnine_unit ninexnine_unit_3710(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E113)
);

ninexnine_unit ninexnine_unit_3711(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F113)
);

assign C3113=c30113+c31113+c32113+c33113+c34113+c35113+c36113+c37113+c38113+c39113+c3A113+c3B113+c3C113+c3D113+c3E113+c3F113;
assign A3113=(C3113>=0)?1:0;

assign P4113=A3113;

ninexnine_unit ninexnine_unit_3712(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30123)
);

ninexnine_unit ninexnine_unit_3713(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31123)
);

ninexnine_unit ninexnine_unit_3714(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32123)
);

ninexnine_unit ninexnine_unit_3715(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33123)
);

ninexnine_unit ninexnine_unit_3716(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34123)
);

ninexnine_unit ninexnine_unit_3717(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35123)
);

ninexnine_unit ninexnine_unit_3718(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36123)
);

ninexnine_unit ninexnine_unit_3719(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37123)
);

ninexnine_unit ninexnine_unit_3720(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38123)
);

ninexnine_unit ninexnine_unit_3721(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39123)
);

ninexnine_unit ninexnine_unit_3722(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A123)
);

ninexnine_unit ninexnine_unit_3723(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B123)
);

ninexnine_unit ninexnine_unit_3724(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C123)
);

ninexnine_unit ninexnine_unit_3725(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D123)
);

ninexnine_unit ninexnine_unit_3726(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E123)
);

ninexnine_unit ninexnine_unit_3727(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F123)
);

assign C3123=c30123+c31123+c32123+c33123+c34123+c35123+c36123+c37123+c38123+c39123+c3A123+c3B123+c3C123+c3D123+c3E123+c3F123;
assign A3123=(C3123>=0)?1:0;

assign P4123=A3123;

ninexnine_unit ninexnine_unit_3728(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30203)
);

ninexnine_unit ninexnine_unit_3729(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31203)
);

ninexnine_unit ninexnine_unit_3730(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32203)
);

ninexnine_unit ninexnine_unit_3731(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33203)
);

ninexnine_unit ninexnine_unit_3732(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34203)
);

ninexnine_unit ninexnine_unit_3733(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35203)
);

ninexnine_unit ninexnine_unit_3734(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36203)
);

ninexnine_unit ninexnine_unit_3735(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37203)
);

ninexnine_unit ninexnine_unit_3736(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38203)
);

ninexnine_unit ninexnine_unit_3737(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39203)
);

ninexnine_unit ninexnine_unit_3738(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A203)
);

ninexnine_unit ninexnine_unit_3739(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B203)
);

ninexnine_unit ninexnine_unit_3740(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C203)
);

ninexnine_unit ninexnine_unit_3741(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D203)
);

ninexnine_unit ninexnine_unit_3742(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E203)
);

ninexnine_unit ninexnine_unit_3743(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F203)
);

assign C3203=c30203+c31203+c32203+c33203+c34203+c35203+c36203+c37203+c38203+c39203+c3A203+c3B203+c3C203+c3D203+c3E203+c3F203;
assign A3203=(C3203>=0)?1:0;

assign P4203=A3203;

ninexnine_unit ninexnine_unit_3744(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30213)
);

ninexnine_unit ninexnine_unit_3745(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31213)
);

ninexnine_unit ninexnine_unit_3746(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32213)
);

ninexnine_unit ninexnine_unit_3747(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33213)
);

ninexnine_unit ninexnine_unit_3748(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34213)
);

ninexnine_unit ninexnine_unit_3749(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35213)
);

ninexnine_unit ninexnine_unit_3750(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36213)
);

ninexnine_unit ninexnine_unit_3751(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37213)
);

ninexnine_unit ninexnine_unit_3752(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38213)
);

ninexnine_unit ninexnine_unit_3753(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39213)
);

ninexnine_unit ninexnine_unit_3754(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A213)
);

ninexnine_unit ninexnine_unit_3755(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B213)
);

ninexnine_unit ninexnine_unit_3756(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C213)
);

ninexnine_unit ninexnine_unit_3757(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D213)
);

ninexnine_unit ninexnine_unit_3758(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E213)
);

ninexnine_unit ninexnine_unit_3759(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F213)
);

assign C3213=c30213+c31213+c32213+c33213+c34213+c35213+c36213+c37213+c38213+c39213+c3A213+c3B213+c3C213+c3D213+c3E213+c3F213;
assign A3213=(C3213>=0)?1:0;

assign P4213=A3213;

ninexnine_unit ninexnine_unit_3760(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W33000),
				.b1(W33010),
				.b2(W33020),
				.b3(W33100),
				.b4(W33110),
				.b5(W33120),
				.b6(W33200),
				.b7(W33210),
				.b8(W33220),
				.c(c30223)
);

ninexnine_unit ninexnine_unit_3761(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W33001),
				.b1(W33011),
				.b2(W33021),
				.b3(W33101),
				.b4(W33111),
				.b5(W33121),
				.b6(W33201),
				.b7(W33211),
				.b8(W33221),
				.c(c31223)
);

ninexnine_unit ninexnine_unit_3762(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W33002),
				.b1(W33012),
				.b2(W33022),
				.b3(W33102),
				.b4(W33112),
				.b5(W33122),
				.b6(W33202),
				.b7(W33212),
				.b8(W33222),
				.c(c32223)
);

ninexnine_unit ninexnine_unit_3763(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W33003),
				.b1(W33013),
				.b2(W33023),
				.b3(W33103),
				.b4(W33113),
				.b5(W33123),
				.b6(W33203),
				.b7(W33213),
				.b8(W33223),
				.c(c33223)
);

ninexnine_unit ninexnine_unit_3764(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W33004),
				.b1(W33014),
				.b2(W33024),
				.b3(W33104),
				.b4(W33114),
				.b5(W33124),
				.b6(W33204),
				.b7(W33214),
				.b8(W33224),
				.c(c34223)
);

ninexnine_unit ninexnine_unit_3765(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W33005),
				.b1(W33015),
				.b2(W33025),
				.b3(W33105),
				.b4(W33115),
				.b5(W33125),
				.b6(W33205),
				.b7(W33215),
				.b8(W33225),
				.c(c35223)
);

ninexnine_unit ninexnine_unit_3766(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W33006),
				.b1(W33016),
				.b2(W33026),
				.b3(W33106),
				.b4(W33116),
				.b5(W33126),
				.b6(W33206),
				.b7(W33216),
				.b8(W33226),
				.c(c36223)
);

ninexnine_unit ninexnine_unit_3767(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W33007),
				.b1(W33017),
				.b2(W33027),
				.b3(W33107),
				.b4(W33117),
				.b5(W33127),
				.b6(W33207),
				.b7(W33217),
				.b8(W33227),
				.c(c37223)
);

ninexnine_unit ninexnine_unit_3768(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W33008),
				.b1(W33018),
				.b2(W33028),
				.b3(W33108),
				.b4(W33118),
				.b5(W33128),
				.b6(W33208),
				.b7(W33218),
				.b8(W33228),
				.c(c38223)
);

ninexnine_unit ninexnine_unit_3769(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W33009),
				.b1(W33019),
				.b2(W33029),
				.b3(W33109),
				.b4(W33119),
				.b5(W33129),
				.b6(W33209),
				.b7(W33219),
				.b8(W33229),
				.c(c39223)
);

ninexnine_unit ninexnine_unit_3770(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3300A),
				.b1(W3301A),
				.b2(W3302A),
				.b3(W3310A),
				.b4(W3311A),
				.b5(W3312A),
				.b6(W3320A),
				.b7(W3321A),
				.b8(W3322A),
				.c(c3A223)
);

ninexnine_unit ninexnine_unit_3771(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3300B),
				.b1(W3301B),
				.b2(W3302B),
				.b3(W3310B),
				.b4(W3311B),
				.b5(W3312B),
				.b6(W3320B),
				.b7(W3321B),
				.b8(W3322B),
				.c(c3B223)
);

ninexnine_unit ninexnine_unit_3772(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3300C),
				.b1(W3301C),
				.b2(W3302C),
				.b3(W3310C),
				.b4(W3311C),
				.b5(W3312C),
				.b6(W3320C),
				.b7(W3321C),
				.b8(W3322C),
				.c(c3C223)
);

ninexnine_unit ninexnine_unit_3773(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3300D),
				.b1(W3301D),
				.b2(W3302D),
				.b3(W3310D),
				.b4(W3311D),
				.b5(W3312D),
				.b6(W3320D),
				.b7(W3321D),
				.b8(W3322D),
				.c(c3D223)
);

ninexnine_unit ninexnine_unit_3774(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3300E),
				.b1(W3301E),
				.b2(W3302E),
				.b3(W3310E),
				.b4(W3311E),
				.b5(W3312E),
				.b6(W3320E),
				.b7(W3321E),
				.b8(W3322E),
				.c(c3E223)
);

ninexnine_unit ninexnine_unit_3775(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3300F),
				.b1(W3301F),
				.b2(W3302F),
				.b3(W3310F),
				.b4(W3311F),
				.b5(W3312F),
				.b6(W3320F),
				.b7(W3321F),
				.b8(W3322F),
				.c(c3F223)
);

assign C3223=c30223+c31223+c32223+c33223+c34223+c35223+c36223+c37223+c38223+c39223+c3A223+c3B223+c3C223+c3D223+c3E223+c3F223;
assign A3223=(C3223>=0)?1:0;

assign P4223=A3223;

ninexnine_unit ninexnine_unit_3776(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30004)
);

ninexnine_unit ninexnine_unit_3777(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31004)
);

ninexnine_unit ninexnine_unit_3778(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32004)
);

ninexnine_unit ninexnine_unit_3779(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33004)
);

ninexnine_unit ninexnine_unit_3780(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34004)
);

ninexnine_unit ninexnine_unit_3781(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35004)
);

ninexnine_unit ninexnine_unit_3782(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36004)
);

ninexnine_unit ninexnine_unit_3783(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37004)
);

ninexnine_unit ninexnine_unit_3784(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38004)
);

ninexnine_unit ninexnine_unit_3785(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39004)
);

ninexnine_unit ninexnine_unit_3786(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A004)
);

ninexnine_unit ninexnine_unit_3787(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B004)
);

ninexnine_unit ninexnine_unit_3788(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C004)
);

ninexnine_unit ninexnine_unit_3789(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D004)
);

ninexnine_unit ninexnine_unit_3790(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E004)
);

ninexnine_unit ninexnine_unit_3791(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F004)
);

assign C3004=c30004+c31004+c32004+c33004+c34004+c35004+c36004+c37004+c38004+c39004+c3A004+c3B004+c3C004+c3D004+c3E004+c3F004;
assign A3004=(C3004>=0)?1:0;

assign P4004=A3004;

ninexnine_unit ninexnine_unit_3792(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30014)
);

ninexnine_unit ninexnine_unit_3793(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31014)
);

ninexnine_unit ninexnine_unit_3794(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32014)
);

ninexnine_unit ninexnine_unit_3795(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33014)
);

ninexnine_unit ninexnine_unit_3796(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34014)
);

ninexnine_unit ninexnine_unit_3797(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35014)
);

ninexnine_unit ninexnine_unit_3798(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36014)
);

ninexnine_unit ninexnine_unit_3799(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37014)
);

ninexnine_unit ninexnine_unit_3800(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38014)
);

ninexnine_unit ninexnine_unit_3801(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39014)
);

ninexnine_unit ninexnine_unit_3802(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A014)
);

ninexnine_unit ninexnine_unit_3803(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B014)
);

ninexnine_unit ninexnine_unit_3804(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C014)
);

ninexnine_unit ninexnine_unit_3805(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D014)
);

ninexnine_unit ninexnine_unit_3806(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E014)
);

ninexnine_unit ninexnine_unit_3807(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F014)
);

assign C3014=c30014+c31014+c32014+c33014+c34014+c35014+c36014+c37014+c38014+c39014+c3A014+c3B014+c3C014+c3D014+c3E014+c3F014;
assign A3014=(C3014>=0)?1:0;

assign P4014=A3014;

ninexnine_unit ninexnine_unit_3808(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30024)
);

ninexnine_unit ninexnine_unit_3809(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31024)
);

ninexnine_unit ninexnine_unit_3810(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32024)
);

ninexnine_unit ninexnine_unit_3811(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33024)
);

ninexnine_unit ninexnine_unit_3812(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34024)
);

ninexnine_unit ninexnine_unit_3813(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35024)
);

ninexnine_unit ninexnine_unit_3814(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36024)
);

ninexnine_unit ninexnine_unit_3815(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37024)
);

ninexnine_unit ninexnine_unit_3816(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38024)
);

ninexnine_unit ninexnine_unit_3817(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39024)
);

ninexnine_unit ninexnine_unit_3818(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A024)
);

ninexnine_unit ninexnine_unit_3819(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B024)
);

ninexnine_unit ninexnine_unit_3820(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C024)
);

ninexnine_unit ninexnine_unit_3821(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D024)
);

ninexnine_unit ninexnine_unit_3822(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E024)
);

ninexnine_unit ninexnine_unit_3823(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F024)
);

assign C3024=c30024+c31024+c32024+c33024+c34024+c35024+c36024+c37024+c38024+c39024+c3A024+c3B024+c3C024+c3D024+c3E024+c3F024;
assign A3024=(C3024>=0)?1:0;

assign P4024=A3024;

ninexnine_unit ninexnine_unit_3824(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30104)
);

ninexnine_unit ninexnine_unit_3825(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31104)
);

ninexnine_unit ninexnine_unit_3826(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32104)
);

ninexnine_unit ninexnine_unit_3827(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33104)
);

ninexnine_unit ninexnine_unit_3828(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34104)
);

ninexnine_unit ninexnine_unit_3829(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35104)
);

ninexnine_unit ninexnine_unit_3830(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36104)
);

ninexnine_unit ninexnine_unit_3831(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37104)
);

ninexnine_unit ninexnine_unit_3832(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38104)
);

ninexnine_unit ninexnine_unit_3833(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39104)
);

ninexnine_unit ninexnine_unit_3834(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A104)
);

ninexnine_unit ninexnine_unit_3835(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B104)
);

ninexnine_unit ninexnine_unit_3836(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C104)
);

ninexnine_unit ninexnine_unit_3837(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D104)
);

ninexnine_unit ninexnine_unit_3838(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E104)
);

ninexnine_unit ninexnine_unit_3839(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F104)
);

assign C3104=c30104+c31104+c32104+c33104+c34104+c35104+c36104+c37104+c38104+c39104+c3A104+c3B104+c3C104+c3D104+c3E104+c3F104;
assign A3104=(C3104>=0)?1:0;

assign P4104=A3104;

ninexnine_unit ninexnine_unit_3840(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30114)
);

ninexnine_unit ninexnine_unit_3841(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31114)
);

ninexnine_unit ninexnine_unit_3842(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32114)
);

ninexnine_unit ninexnine_unit_3843(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33114)
);

ninexnine_unit ninexnine_unit_3844(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34114)
);

ninexnine_unit ninexnine_unit_3845(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35114)
);

ninexnine_unit ninexnine_unit_3846(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36114)
);

ninexnine_unit ninexnine_unit_3847(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37114)
);

ninexnine_unit ninexnine_unit_3848(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38114)
);

ninexnine_unit ninexnine_unit_3849(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39114)
);

ninexnine_unit ninexnine_unit_3850(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A114)
);

ninexnine_unit ninexnine_unit_3851(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B114)
);

ninexnine_unit ninexnine_unit_3852(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C114)
);

ninexnine_unit ninexnine_unit_3853(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D114)
);

ninexnine_unit ninexnine_unit_3854(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E114)
);

ninexnine_unit ninexnine_unit_3855(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F114)
);

assign C3114=c30114+c31114+c32114+c33114+c34114+c35114+c36114+c37114+c38114+c39114+c3A114+c3B114+c3C114+c3D114+c3E114+c3F114;
assign A3114=(C3114>=0)?1:0;

assign P4114=A3114;

ninexnine_unit ninexnine_unit_3856(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30124)
);

ninexnine_unit ninexnine_unit_3857(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31124)
);

ninexnine_unit ninexnine_unit_3858(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32124)
);

ninexnine_unit ninexnine_unit_3859(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33124)
);

ninexnine_unit ninexnine_unit_3860(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34124)
);

ninexnine_unit ninexnine_unit_3861(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35124)
);

ninexnine_unit ninexnine_unit_3862(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36124)
);

ninexnine_unit ninexnine_unit_3863(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37124)
);

ninexnine_unit ninexnine_unit_3864(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38124)
);

ninexnine_unit ninexnine_unit_3865(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39124)
);

ninexnine_unit ninexnine_unit_3866(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A124)
);

ninexnine_unit ninexnine_unit_3867(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B124)
);

ninexnine_unit ninexnine_unit_3868(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C124)
);

ninexnine_unit ninexnine_unit_3869(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D124)
);

ninexnine_unit ninexnine_unit_3870(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E124)
);

ninexnine_unit ninexnine_unit_3871(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F124)
);

assign C3124=c30124+c31124+c32124+c33124+c34124+c35124+c36124+c37124+c38124+c39124+c3A124+c3B124+c3C124+c3D124+c3E124+c3F124;
assign A3124=(C3124>=0)?1:0;

assign P4124=A3124;

ninexnine_unit ninexnine_unit_3872(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30204)
);

ninexnine_unit ninexnine_unit_3873(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31204)
);

ninexnine_unit ninexnine_unit_3874(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32204)
);

ninexnine_unit ninexnine_unit_3875(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33204)
);

ninexnine_unit ninexnine_unit_3876(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34204)
);

ninexnine_unit ninexnine_unit_3877(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35204)
);

ninexnine_unit ninexnine_unit_3878(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36204)
);

ninexnine_unit ninexnine_unit_3879(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37204)
);

ninexnine_unit ninexnine_unit_3880(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38204)
);

ninexnine_unit ninexnine_unit_3881(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39204)
);

ninexnine_unit ninexnine_unit_3882(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A204)
);

ninexnine_unit ninexnine_unit_3883(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B204)
);

ninexnine_unit ninexnine_unit_3884(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C204)
);

ninexnine_unit ninexnine_unit_3885(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D204)
);

ninexnine_unit ninexnine_unit_3886(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E204)
);

ninexnine_unit ninexnine_unit_3887(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F204)
);

assign C3204=c30204+c31204+c32204+c33204+c34204+c35204+c36204+c37204+c38204+c39204+c3A204+c3B204+c3C204+c3D204+c3E204+c3F204;
assign A3204=(C3204>=0)?1:0;

assign P4204=A3204;

ninexnine_unit ninexnine_unit_3888(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30214)
);

ninexnine_unit ninexnine_unit_3889(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31214)
);

ninexnine_unit ninexnine_unit_3890(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32214)
);

ninexnine_unit ninexnine_unit_3891(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33214)
);

ninexnine_unit ninexnine_unit_3892(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34214)
);

ninexnine_unit ninexnine_unit_3893(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35214)
);

ninexnine_unit ninexnine_unit_3894(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36214)
);

ninexnine_unit ninexnine_unit_3895(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37214)
);

ninexnine_unit ninexnine_unit_3896(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38214)
);

ninexnine_unit ninexnine_unit_3897(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39214)
);

ninexnine_unit ninexnine_unit_3898(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A214)
);

ninexnine_unit ninexnine_unit_3899(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B214)
);

ninexnine_unit ninexnine_unit_3900(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C214)
);

ninexnine_unit ninexnine_unit_3901(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D214)
);

ninexnine_unit ninexnine_unit_3902(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E214)
);

ninexnine_unit ninexnine_unit_3903(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F214)
);

assign C3214=c30214+c31214+c32214+c33214+c34214+c35214+c36214+c37214+c38214+c39214+c3A214+c3B214+c3C214+c3D214+c3E214+c3F214;
assign A3214=(C3214>=0)?1:0;

assign P4214=A3214;

ninexnine_unit ninexnine_unit_3904(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W34000),
				.b1(W34010),
				.b2(W34020),
				.b3(W34100),
				.b4(W34110),
				.b5(W34120),
				.b6(W34200),
				.b7(W34210),
				.b8(W34220),
				.c(c30224)
);

ninexnine_unit ninexnine_unit_3905(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W34001),
				.b1(W34011),
				.b2(W34021),
				.b3(W34101),
				.b4(W34111),
				.b5(W34121),
				.b6(W34201),
				.b7(W34211),
				.b8(W34221),
				.c(c31224)
);

ninexnine_unit ninexnine_unit_3906(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W34002),
				.b1(W34012),
				.b2(W34022),
				.b3(W34102),
				.b4(W34112),
				.b5(W34122),
				.b6(W34202),
				.b7(W34212),
				.b8(W34222),
				.c(c32224)
);

ninexnine_unit ninexnine_unit_3907(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W34003),
				.b1(W34013),
				.b2(W34023),
				.b3(W34103),
				.b4(W34113),
				.b5(W34123),
				.b6(W34203),
				.b7(W34213),
				.b8(W34223),
				.c(c33224)
);

ninexnine_unit ninexnine_unit_3908(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W34004),
				.b1(W34014),
				.b2(W34024),
				.b3(W34104),
				.b4(W34114),
				.b5(W34124),
				.b6(W34204),
				.b7(W34214),
				.b8(W34224),
				.c(c34224)
);

ninexnine_unit ninexnine_unit_3909(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W34005),
				.b1(W34015),
				.b2(W34025),
				.b3(W34105),
				.b4(W34115),
				.b5(W34125),
				.b6(W34205),
				.b7(W34215),
				.b8(W34225),
				.c(c35224)
);

ninexnine_unit ninexnine_unit_3910(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W34006),
				.b1(W34016),
				.b2(W34026),
				.b3(W34106),
				.b4(W34116),
				.b5(W34126),
				.b6(W34206),
				.b7(W34216),
				.b8(W34226),
				.c(c36224)
);

ninexnine_unit ninexnine_unit_3911(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W34007),
				.b1(W34017),
				.b2(W34027),
				.b3(W34107),
				.b4(W34117),
				.b5(W34127),
				.b6(W34207),
				.b7(W34217),
				.b8(W34227),
				.c(c37224)
);

ninexnine_unit ninexnine_unit_3912(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W34008),
				.b1(W34018),
				.b2(W34028),
				.b3(W34108),
				.b4(W34118),
				.b5(W34128),
				.b6(W34208),
				.b7(W34218),
				.b8(W34228),
				.c(c38224)
);

ninexnine_unit ninexnine_unit_3913(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W34009),
				.b1(W34019),
				.b2(W34029),
				.b3(W34109),
				.b4(W34119),
				.b5(W34129),
				.b6(W34209),
				.b7(W34219),
				.b8(W34229),
				.c(c39224)
);

ninexnine_unit ninexnine_unit_3914(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3400A),
				.b1(W3401A),
				.b2(W3402A),
				.b3(W3410A),
				.b4(W3411A),
				.b5(W3412A),
				.b6(W3420A),
				.b7(W3421A),
				.b8(W3422A),
				.c(c3A224)
);

ninexnine_unit ninexnine_unit_3915(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3400B),
				.b1(W3401B),
				.b2(W3402B),
				.b3(W3410B),
				.b4(W3411B),
				.b5(W3412B),
				.b6(W3420B),
				.b7(W3421B),
				.b8(W3422B),
				.c(c3B224)
);

ninexnine_unit ninexnine_unit_3916(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3400C),
				.b1(W3401C),
				.b2(W3402C),
				.b3(W3410C),
				.b4(W3411C),
				.b5(W3412C),
				.b6(W3420C),
				.b7(W3421C),
				.b8(W3422C),
				.c(c3C224)
);

ninexnine_unit ninexnine_unit_3917(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3400D),
				.b1(W3401D),
				.b2(W3402D),
				.b3(W3410D),
				.b4(W3411D),
				.b5(W3412D),
				.b6(W3420D),
				.b7(W3421D),
				.b8(W3422D),
				.c(c3D224)
);

ninexnine_unit ninexnine_unit_3918(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3400E),
				.b1(W3401E),
				.b2(W3402E),
				.b3(W3410E),
				.b4(W3411E),
				.b5(W3412E),
				.b6(W3420E),
				.b7(W3421E),
				.b8(W3422E),
				.c(c3E224)
);

ninexnine_unit ninexnine_unit_3919(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3400F),
				.b1(W3401F),
				.b2(W3402F),
				.b3(W3410F),
				.b4(W3411F),
				.b5(W3412F),
				.b6(W3420F),
				.b7(W3421F),
				.b8(W3422F),
				.c(c3F224)
);

assign C3224=c30224+c31224+c32224+c33224+c34224+c35224+c36224+c37224+c38224+c39224+c3A224+c3B224+c3C224+c3D224+c3E224+c3F224;
assign A3224=(C3224>=0)?1:0;

assign P4224=A3224;

ninexnine_unit ninexnine_unit_3920(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30005)
);

ninexnine_unit ninexnine_unit_3921(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31005)
);

ninexnine_unit ninexnine_unit_3922(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32005)
);

ninexnine_unit ninexnine_unit_3923(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33005)
);

ninexnine_unit ninexnine_unit_3924(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34005)
);

ninexnine_unit ninexnine_unit_3925(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35005)
);

ninexnine_unit ninexnine_unit_3926(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36005)
);

ninexnine_unit ninexnine_unit_3927(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37005)
);

ninexnine_unit ninexnine_unit_3928(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38005)
);

ninexnine_unit ninexnine_unit_3929(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39005)
);

ninexnine_unit ninexnine_unit_3930(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A005)
);

ninexnine_unit ninexnine_unit_3931(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B005)
);

ninexnine_unit ninexnine_unit_3932(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C005)
);

ninexnine_unit ninexnine_unit_3933(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D005)
);

ninexnine_unit ninexnine_unit_3934(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E005)
);

ninexnine_unit ninexnine_unit_3935(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F005)
);

assign C3005=c30005+c31005+c32005+c33005+c34005+c35005+c36005+c37005+c38005+c39005+c3A005+c3B005+c3C005+c3D005+c3E005+c3F005;
assign A3005=(C3005>=0)?1:0;

assign P4005=A3005;

ninexnine_unit ninexnine_unit_3936(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30015)
);

ninexnine_unit ninexnine_unit_3937(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31015)
);

ninexnine_unit ninexnine_unit_3938(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32015)
);

ninexnine_unit ninexnine_unit_3939(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33015)
);

ninexnine_unit ninexnine_unit_3940(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34015)
);

ninexnine_unit ninexnine_unit_3941(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35015)
);

ninexnine_unit ninexnine_unit_3942(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36015)
);

ninexnine_unit ninexnine_unit_3943(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37015)
);

ninexnine_unit ninexnine_unit_3944(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38015)
);

ninexnine_unit ninexnine_unit_3945(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39015)
);

ninexnine_unit ninexnine_unit_3946(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A015)
);

ninexnine_unit ninexnine_unit_3947(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B015)
);

ninexnine_unit ninexnine_unit_3948(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C015)
);

ninexnine_unit ninexnine_unit_3949(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D015)
);

ninexnine_unit ninexnine_unit_3950(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E015)
);

ninexnine_unit ninexnine_unit_3951(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F015)
);

assign C3015=c30015+c31015+c32015+c33015+c34015+c35015+c36015+c37015+c38015+c39015+c3A015+c3B015+c3C015+c3D015+c3E015+c3F015;
assign A3015=(C3015>=0)?1:0;

assign P4015=A3015;

ninexnine_unit ninexnine_unit_3952(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30025)
);

ninexnine_unit ninexnine_unit_3953(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31025)
);

ninexnine_unit ninexnine_unit_3954(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32025)
);

ninexnine_unit ninexnine_unit_3955(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33025)
);

ninexnine_unit ninexnine_unit_3956(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34025)
);

ninexnine_unit ninexnine_unit_3957(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35025)
);

ninexnine_unit ninexnine_unit_3958(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36025)
);

ninexnine_unit ninexnine_unit_3959(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37025)
);

ninexnine_unit ninexnine_unit_3960(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38025)
);

ninexnine_unit ninexnine_unit_3961(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39025)
);

ninexnine_unit ninexnine_unit_3962(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A025)
);

ninexnine_unit ninexnine_unit_3963(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B025)
);

ninexnine_unit ninexnine_unit_3964(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C025)
);

ninexnine_unit ninexnine_unit_3965(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D025)
);

ninexnine_unit ninexnine_unit_3966(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E025)
);

ninexnine_unit ninexnine_unit_3967(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F025)
);

assign C3025=c30025+c31025+c32025+c33025+c34025+c35025+c36025+c37025+c38025+c39025+c3A025+c3B025+c3C025+c3D025+c3E025+c3F025;
assign A3025=(C3025>=0)?1:0;

assign P4025=A3025;

ninexnine_unit ninexnine_unit_3968(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30105)
);

ninexnine_unit ninexnine_unit_3969(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31105)
);

ninexnine_unit ninexnine_unit_3970(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32105)
);

ninexnine_unit ninexnine_unit_3971(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33105)
);

ninexnine_unit ninexnine_unit_3972(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34105)
);

ninexnine_unit ninexnine_unit_3973(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35105)
);

ninexnine_unit ninexnine_unit_3974(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36105)
);

ninexnine_unit ninexnine_unit_3975(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37105)
);

ninexnine_unit ninexnine_unit_3976(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38105)
);

ninexnine_unit ninexnine_unit_3977(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39105)
);

ninexnine_unit ninexnine_unit_3978(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A105)
);

ninexnine_unit ninexnine_unit_3979(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B105)
);

ninexnine_unit ninexnine_unit_3980(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C105)
);

ninexnine_unit ninexnine_unit_3981(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D105)
);

ninexnine_unit ninexnine_unit_3982(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E105)
);

ninexnine_unit ninexnine_unit_3983(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F105)
);

assign C3105=c30105+c31105+c32105+c33105+c34105+c35105+c36105+c37105+c38105+c39105+c3A105+c3B105+c3C105+c3D105+c3E105+c3F105;
assign A3105=(C3105>=0)?1:0;

assign P4105=A3105;

ninexnine_unit ninexnine_unit_3984(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30115)
);

ninexnine_unit ninexnine_unit_3985(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31115)
);

ninexnine_unit ninexnine_unit_3986(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32115)
);

ninexnine_unit ninexnine_unit_3987(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33115)
);

ninexnine_unit ninexnine_unit_3988(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34115)
);

ninexnine_unit ninexnine_unit_3989(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35115)
);

ninexnine_unit ninexnine_unit_3990(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36115)
);

ninexnine_unit ninexnine_unit_3991(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37115)
);

ninexnine_unit ninexnine_unit_3992(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38115)
);

ninexnine_unit ninexnine_unit_3993(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39115)
);

ninexnine_unit ninexnine_unit_3994(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A115)
);

ninexnine_unit ninexnine_unit_3995(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B115)
);

ninexnine_unit ninexnine_unit_3996(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C115)
);

ninexnine_unit ninexnine_unit_3997(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D115)
);

ninexnine_unit ninexnine_unit_3998(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E115)
);

ninexnine_unit ninexnine_unit_3999(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F115)
);

assign C3115=c30115+c31115+c32115+c33115+c34115+c35115+c36115+c37115+c38115+c39115+c3A115+c3B115+c3C115+c3D115+c3E115+c3F115;
assign A3115=(C3115>=0)?1:0;

assign P4115=A3115;

ninexnine_unit ninexnine_unit_4000(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30125)
);

ninexnine_unit ninexnine_unit_4001(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31125)
);

ninexnine_unit ninexnine_unit_4002(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32125)
);

ninexnine_unit ninexnine_unit_4003(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33125)
);

ninexnine_unit ninexnine_unit_4004(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34125)
);

ninexnine_unit ninexnine_unit_4005(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35125)
);

ninexnine_unit ninexnine_unit_4006(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36125)
);

ninexnine_unit ninexnine_unit_4007(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37125)
);

ninexnine_unit ninexnine_unit_4008(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38125)
);

ninexnine_unit ninexnine_unit_4009(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39125)
);

ninexnine_unit ninexnine_unit_4010(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A125)
);

ninexnine_unit ninexnine_unit_4011(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B125)
);

ninexnine_unit ninexnine_unit_4012(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C125)
);

ninexnine_unit ninexnine_unit_4013(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D125)
);

ninexnine_unit ninexnine_unit_4014(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E125)
);

ninexnine_unit ninexnine_unit_4015(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F125)
);

assign C3125=c30125+c31125+c32125+c33125+c34125+c35125+c36125+c37125+c38125+c39125+c3A125+c3B125+c3C125+c3D125+c3E125+c3F125;
assign A3125=(C3125>=0)?1:0;

assign P4125=A3125;

ninexnine_unit ninexnine_unit_4016(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30205)
);

ninexnine_unit ninexnine_unit_4017(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31205)
);

ninexnine_unit ninexnine_unit_4018(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32205)
);

ninexnine_unit ninexnine_unit_4019(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33205)
);

ninexnine_unit ninexnine_unit_4020(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34205)
);

ninexnine_unit ninexnine_unit_4021(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35205)
);

ninexnine_unit ninexnine_unit_4022(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36205)
);

ninexnine_unit ninexnine_unit_4023(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37205)
);

ninexnine_unit ninexnine_unit_4024(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38205)
);

ninexnine_unit ninexnine_unit_4025(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39205)
);

ninexnine_unit ninexnine_unit_4026(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A205)
);

ninexnine_unit ninexnine_unit_4027(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B205)
);

ninexnine_unit ninexnine_unit_4028(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C205)
);

ninexnine_unit ninexnine_unit_4029(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D205)
);

ninexnine_unit ninexnine_unit_4030(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E205)
);

ninexnine_unit ninexnine_unit_4031(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F205)
);

assign C3205=c30205+c31205+c32205+c33205+c34205+c35205+c36205+c37205+c38205+c39205+c3A205+c3B205+c3C205+c3D205+c3E205+c3F205;
assign A3205=(C3205>=0)?1:0;

assign P4205=A3205;

ninexnine_unit ninexnine_unit_4032(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30215)
);

ninexnine_unit ninexnine_unit_4033(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31215)
);

ninexnine_unit ninexnine_unit_4034(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32215)
);

ninexnine_unit ninexnine_unit_4035(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33215)
);

ninexnine_unit ninexnine_unit_4036(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34215)
);

ninexnine_unit ninexnine_unit_4037(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35215)
);

ninexnine_unit ninexnine_unit_4038(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36215)
);

ninexnine_unit ninexnine_unit_4039(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37215)
);

ninexnine_unit ninexnine_unit_4040(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38215)
);

ninexnine_unit ninexnine_unit_4041(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39215)
);

ninexnine_unit ninexnine_unit_4042(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A215)
);

ninexnine_unit ninexnine_unit_4043(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B215)
);

ninexnine_unit ninexnine_unit_4044(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C215)
);

ninexnine_unit ninexnine_unit_4045(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D215)
);

ninexnine_unit ninexnine_unit_4046(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E215)
);

ninexnine_unit ninexnine_unit_4047(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F215)
);

assign C3215=c30215+c31215+c32215+c33215+c34215+c35215+c36215+c37215+c38215+c39215+c3A215+c3B215+c3C215+c3D215+c3E215+c3F215;
assign A3215=(C3215>=0)?1:0;

assign P4215=A3215;

ninexnine_unit ninexnine_unit_4048(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W35000),
				.b1(W35010),
				.b2(W35020),
				.b3(W35100),
				.b4(W35110),
				.b5(W35120),
				.b6(W35200),
				.b7(W35210),
				.b8(W35220),
				.c(c30225)
);

ninexnine_unit ninexnine_unit_4049(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W35001),
				.b1(W35011),
				.b2(W35021),
				.b3(W35101),
				.b4(W35111),
				.b5(W35121),
				.b6(W35201),
				.b7(W35211),
				.b8(W35221),
				.c(c31225)
);

ninexnine_unit ninexnine_unit_4050(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W35002),
				.b1(W35012),
				.b2(W35022),
				.b3(W35102),
				.b4(W35112),
				.b5(W35122),
				.b6(W35202),
				.b7(W35212),
				.b8(W35222),
				.c(c32225)
);

ninexnine_unit ninexnine_unit_4051(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W35003),
				.b1(W35013),
				.b2(W35023),
				.b3(W35103),
				.b4(W35113),
				.b5(W35123),
				.b6(W35203),
				.b7(W35213),
				.b8(W35223),
				.c(c33225)
);

ninexnine_unit ninexnine_unit_4052(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W35004),
				.b1(W35014),
				.b2(W35024),
				.b3(W35104),
				.b4(W35114),
				.b5(W35124),
				.b6(W35204),
				.b7(W35214),
				.b8(W35224),
				.c(c34225)
);

ninexnine_unit ninexnine_unit_4053(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W35005),
				.b1(W35015),
				.b2(W35025),
				.b3(W35105),
				.b4(W35115),
				.b5(W35125),
				.b6(W35205),
				.b7(W35215),
				.b8(W35225),
				.c(c35225)
);

ninexnine_unit ninexnine_unit_4054(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W35006),
				.b1(W35016),
				.b2(W35026),
				.b3(W35106),
				.b4(W35116),
				.b5(W35126),
				.b6(W35206),
				.b7(W35216),
				.b8(W35226),
				.c(c36225)
);

ninexnine_unit ninexnine_unit_4055(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W35007),
				.b1(W35017),
				.b2(W35027),
				.b3(W35107),
				.b4(W35117),
				.b5(W35127),
				.b6(W35207),
				.b7(W35217),
				.b8(W35227),
				.c(c37225)
);

ninexnine_unit ninexnine_unit_4056(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W35008),
				.b1(W35018),
				.b2(W35028),
				.b3(W35108),
				.b4(W35118),
				.b5(W35128),
				.b6(W35208),
				.b7(W35218),
				.b8(W35228),
				.c(c38225)
);

ninexnine_unit ninexnine_unit_4057(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W35009),
				.b1(W35019),
				.b2(W35029),
				.b3(W35109),
				.b4(W35119),
				.b5(W35129),
				.b6(W35209),
				.b7(W35219),
				.b8(W35229),
				.c(c39225)
);

ninexnine_unit ninexnine_unit_4058(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3500A),
				.b1(W3501A),
				.b2(W3502A),
				.b3(W3510A),
				.b4(W3511A),
				.b5(W3512A),
				.b6(W3520A),
				.b7(W3521A),
				.b8(W3522A),
				.c(c3A225)
);

ninexnine_unit ninexnine_unit_4059(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3500B),
				.b1(W3501B),
				.b2(W3502B),
				.b3(W3510B),
				.b4(W3511B),
				.b5(W3512B),
				.b6(W3520B),
				.b7(W3521B),
				.b8(W3522B),
				.c(c3B225)
);

ninexnine_unit ninexnine_unit_4060(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3500C),
				.b1(W3501C),
				.b2(W3502C),
				.b3(W3510C),
				.b4(W3511C),
				.b5(W3512C),
				.b6(W3520C),
				.b7(W3521C),
				.b8(W3522C),
				.c(c3C225)
);

ninexnine_unit ninexnine_unit_4061(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3500D),
				.b1(W3501D),
				.b2(W3502D),
				.b3(W3510D),
				.b4(W3511D),
				.b5(W3512D),
				.b6(W3520D),
				.b7(W3521D),
				.b8(W3522D),
				.c(c3D225)
);

ninexnine_unit ninexnine_unit_4062(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3500E),
				.b1(W3501E),
				.b2(W3502E),
				.b3(W3510E),
				.b4(W3511E),
				.b5(W3512E),
				.b6(W3520E),
				.b7(W3521E),
				.b8(W3522E),
				.c(c3E225)
);

ninexnine_unit ninexnine_unit_4063(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3500F),
				.b1(W3501F),
				.b2(W3502F),
				.b3(W3510F),
				.b4(W3511F),
				.b5(W3512F),
				.b6(W3520F),
				.b7(W3521F),
				.b8(W3522F),
				.c(c3F225)
);

assign C3225=c30225+c31225+c32225+c33225+c34225+c35225+c36225+c37225+c38225+c39225+c3A225+c3B225+c3C225+c3D225+c3E225+c3F225;
assign A3225=(C3225>=0)?1:0;

assign P4225=A3225;

ninexnine_unit ninexnine_unit_4064(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30006)
);

ninexnine_unit ninexnine_unit_4065(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31006)
);

ninexnine_unit ninexnine_unit_4066(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32006)
);

ninexnine_unit ninexnine_unit_4067(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33006)
);

ninexnine_unit ninexnine_unit_4068(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34006)
);

ninexnine_unit ninexnine_unit_4069(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35006)
);

ninexnine_unit ninexnine_unit_4070(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36006)
);

ninexnine_unit ninexnine_unit_4071(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37006)
);

ninexnine_unit ninexnine_unit_4072(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38006)
);

ninexnine_unit ninexnine_unit_4073(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39006)
);

ninexnine_unit ninexnine_unit_4074(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A006)
);

ninexnine_unit ninexnine_unit_4075(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B006)
);

ninexnine_unit ninexnine_unit_4076(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C006)
);

ninexnine_unit ninexnine_unit_4077(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D006)
);

ninexnine_unit ninexnine_unit_4078(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E006)
);

ninexnine_unit ninexnine_unit_4079(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F006)
);

assign C3006=c30006+c31006+c32006+c33006+c34006+c35006+c36006+c37006+c38006+c39006+c3A006+c3B006+c3C006+c3D006+c3E006+c3F006;
assign A3006=(C3006>=0)?1:0;

assign P4006=A3006;

ninexnine_unit ninexnine_unit_4080(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30016)
);

ninexnine_unit ninexnine_unit_4081(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31016)
);

ninexnine_unit ninexnine_unit_4082(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32016)
);

ninexnine_unit ninexnine_unit_4083(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33016)
);

ninexnine_unit ninexnine_unit_4084(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34016)
);

ninexnine_unit ninexnine_unit_4085(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35016)
);

ninexnine_unit ninexnine_unit_4086(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36016)
);

ninexnine_unit ninexnine_unit_4087(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37016)
);

ninexnine_unit ninexnine_unit_4088(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38016)
);

ninexnine_unit ninexnine_unit_4089(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39016)
);

ninexnine_unit ninexnine_unit_4090(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A016)
);

ninexnine_unit ninexnine_unit_4091(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B016)
);

ninexnine_unit ninexnine_unit_4092(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C016)
);

ninexnine_unit ninexnine_unit_4093(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D016)
);

ninexnine_unit ninexnine_unit_4094(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E016)
);

ninexnine_unit ninexnine_unit_4095(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F016)
);

assign C3016=c30016+c31016+c32016+c33016+c34016+c35016+c36016+c37016+c38016+c39016+c3A016+c3B016+c3C016+c3D016+c3E016+c3F016;
assign A3016=(C3016>=0)?1:0;

assign P4016=A3016;

ninexnine_unit ninexnine_unit_4096(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30026)
);

ninexnine_unit ninexnine_unit_4097(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31026)
);

ninexnine_unit ninexnine_unit_4098(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32026)
);

ninexnine_unit ninexnine_unit_4099(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33026)
);

ninexnine_unit ninexnine_unit_4100(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34026)
);

ninexnine_unit ninexnine_unit_4101(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35026)
);

ninexnine_unit ninexnine_unit_4102(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36026)
);

ninexnine_unit ninexnine_unit_4103(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37026)
);

ninexnine_unit ninexnine_unit_4104(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38026)
);

ninexnine_unit ninexnine_unit_4105(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39026)
);

ninexnine_unit ninexnine_unit_4106(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A026)
);

ninexnine_unit ninexnine_unit_4107(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B026)
);

ninexnine_unit ninexnine_unit_4108(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C026)
);

ninexnine_unit ninexnine_unit_4109(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D026)
);

ninexnine_unit ninexnine_unit_4110(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E026)
);

ninexnine_unit ninexnine_unit_4111(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F026)
);

assign C3026=c30026+c31026+c32026+c33026+c34026+c35026+c36026+c37026+c38026+c39026+c3A026+c3B026+c3C026+c3D026+c3E026+c3F026;
assign A3026=(C3026>=0)?1:0;

assign P4026=A3026;

ninexnine_unit ninexnine_unit_4112(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30106)
);

ninexnine_unit ninexnine_unit_4113(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31106)
);

ninexnine_unit ninexnine_unit_4114(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32106)
);

ninexnine_unit ninexnine_unit_4115(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33106)
);

ninexnine_unit ninexnine_unit_4116(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34106)
);

ninexnine_unit ninexnine_unit_4117(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35106)
);

ninexnine_unit ninexnine_unit_4118(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36106)
);

ninexnine_unit ninexnine_unit_4119(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37106)
);

ninexnine_unit ninexnine_unit_4120(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38106)
);

ninexnine_unit ninexnine_unit_4121(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39106)
);

ninexnine_unit ninexnine_unit_4122(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A106)
);

ninexnine_unit ninexnine_unit_4123(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B106)
);

ninexnine_unit ninexnine_unit_4124(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C106)
);

ninexnine_unit ninexnine_unit_4125(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D106)
);

ninexnine_unit ninexnine_unit_4126(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E106)
);

ninexnine_unit ninexnine_unit_4127(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F106)
);

assign C3106=c30106+c31106+c32106+c33106+c34106+c35106+c36106+c37106+c38106+c39106+c3A106+c3B106+c3C106+c3D106+c3E106+c3F106;
assign A3106=(C3106>=0)?1:0;

assign P4106=A3106;

ninexnine_unit ninexnine_unit_4128(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30116)
);

ninexnine_unit ninexnine_unit_4129(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31116)
);

ninexnine_unit ninexnine_unit_4130(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32116)
);

ninexnine_unit ninexnine_unit_4131(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33116)
);

ninexnine_unit ninexnine_unit_4132(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34116)
);

ninexnine_unit ninexnine_unit_4133(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35116)
);

ninexnine_unit ninexnine_unit_4134(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36116)
);

ninexnine_unit ninexnine_unit_4135(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37116)
);

ninexnine_unit ninexnine_unit_4136(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38116)
);

ninexnine_unit ninexnine_unit_4137(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39116)
);

ninexnine_unit ninexnine_unit_4138(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A116)
);

ninexnine_unit ninexnine_unit_4139(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B116)
);

ninexnine_unit ninexnine_unit_4140(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C116)
);

ninexnine_unit ninexnine_unit_4141(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D116)
);

ninexnine_unit ninexnine_unit_4142(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E116)
);

ninexnine_unit ninexnine_unit_4143(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F116)
);

assign C3116=c30116+c31116+c32116+c33116+c34116+c35116+c36116+c37116+c38116+c39116+c3A116+c3B116+c3C116+c3D116+c3E116+c3F116;
assign A3116=(C3116>=0)?1:0;

assign P4116=A3116;

ninexnine_unit ninexnine_unit_4144(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30126)
);

ninexnine_unit ninexnine_unit_4145(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31126)
);

ninexnine_unit ninexnine_unit_4146(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32126)
);

ninexnine_unit ninexnine_unit_4147(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33126)
);

ninexnine_unit ninexnine_unit_4148(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34126)
);

ninexnine_unit ninexnine_unit_4149(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35126)
);

ninexnine_unit ninexnine_unit_4150(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36126)
);

ninexnine_unit ninexnine_unit_4151(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37126)
);

ninexnine_unit ninexnine_unit_4152(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38126)
);

ninexnine_unit ninexnine_unit_4153(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39126)
);

ninexnine_unit ninexnine_unit_4154(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A126)
);

ninexnine_unit ninexnine_unit_4155(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B126)
);

ninexnine_unit ninexnine_unit_4156(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C126)
);

ninexnine_unit ninexnine_unit_4157(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D126)
);

ninexnine_unit ninexnine_unit_4158(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E126)
);

ninexnine_unit ninexnine_unit_4159(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F126)
);

assign C3126=c30126+c31126+c32126+c33126+c34126+c35126+c36126+c37126+c38126+c39126+c3A126+c3B126+c3C126+c3D126+c3E126+c3F126;
assign A3126=(C3126>=0)?1:0;

assign P4126=A3126;

ninexnine_unit ninexnine_unit_4160(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30206)
);

ninexnine_unit ninexnine_unit_4161(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31206)
);

ninexnine_unit ninexnine_unit_4162(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32206)
);

ninexnine_unit ninexnine_unit_4163(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33206)
);

ninexnine_unit ninexnine_unit_4164(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34206)
);

ninexnine_unit ninexnine_unit_4165(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35206)
);

ninexnine_unit ninexnine_unit_4166(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36206)
);

ninexnine_unit ninexnine_unit_4167(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37206)
);

ninexnine_unit ninexnine_unit_4168(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38206)
);

ninexnine_unit ninexnine_unit_4169(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39206)
);

ninexnine_unit ninexnine_unit_4170(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A206)
);

ninexnine_unit ninexnine_unit_4171(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B206)
);

ninexnine_unit ninexnine_unit_4172(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C206)
);

ninexnine_unit ninexnine_unit_4173(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D206)
);

ninexnine_unit ninexnine_unit_4174(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E206)
);

ninexnine_unit ninexnine_unit_4175(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F206)
);

assign C3206=c30206+c31206+c32206+c33206+c34206+c35206+c36206+c37206+c38206+c39206+c3A206+c3B206+c3C206+c3D206+c3E206+c3F206;
assign A3206=(C3206>=0)?1:0;

assign P4206=A3206;

ninexnine_unit ninexnine_unit_4176(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30216)
);

ninexnine_unit ninexnine_unit_4177(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31216)
);

ninexnine_unit ninexnine_unit_4178(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32216)
);

ninexnine_unit ninexnine_unit_4179(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33216)
);

ninexnine_unit ninexnine_unit_4180(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34216)
);

ninexnine_unit ninexnine_unit_4181(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35216)
);

ninexnine_unit ninexnine_unit_4182(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36216)
);

ninexnine_unit ninexnine_unit_4183(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37216)
);

ninexnine_unit ninexnine_unit_4184(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38216)
);

ninexnine_unit ninexnine_unit_4185(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39216)
);

ninexnine_unit ninexnine_unit_4186(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A216)
);

ninexnine_unit ninexnine_unit_4187(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B216)
);

ninexnine_unit ninexnine_unit_4188(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C216)
);

ninexnine_unit ninexnine_unit_4189(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D216)
);

ninexnine_unit ninexnine_unit_4190(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E216)
);

ninexnine_unit ninexnine_unit_4191(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F216)
);

assign C3216=c30216+c31216+c32216+c33216+c34216+c35216+c36216+c37216+c38216+c39216+c3A216+c3B216+c3C216+c3D216+c3E216+c3F216;
assign A3216=(C3216>=0)?1:0;

assign P4216=A3216;

ninexnine_unit ninexnine_unit_4192(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W36000),
				.b1(W36010),
				.b2(W36020),
				.b3(W36100),
				.b4(W36110),
				.b5(W36120),
				.b6(W36200),
				.b7(W36210),
				.b8(W36220),
				.c(c30226)
);

ninexnine_unit ninexnine_unit_4193(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W36001),
				.b1(W36011),
				.b2(W36021),
				.b3(W36101),
				.b4(W36111),
				.b5(W36121),
				.b6(W36201),
				.b7(W36211),
				.b8(W36221),
				.c(c31226)
);

ninexnine_unit ninexnine_unit_4194(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W36002),
				.b1(W36012),
				.b2(W36022),
				.b3(W36102),
				.b4(W36112),
				.b5(W36122),
				.b6(W36202),
				.b7(W36212),
				.b8(W36222),
				.c(c32226)
);

ninexnine_unit ninexnine_unit_4195(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W36003),
				.b1(W36013),
				.b2(W36023),
				.b3(W36103),
				.b4(W36113),
				.b5(W36123),
				.b6(W36203),
				.b7(W36213),
				.b8(W36223),
				.c(c33226)
);

ninexnine_unit ninexnine_unit_4196(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W36004),
				.b1(W36014),
				.b2(W36024),
				.b3(W36104),
				.b4(W36114),
				.b5(W36124),
				.b6(W36204),
				.b7(W36214),
				.b8(W36224),
				.c(c34226)
);

ninexnine_unit ninexnine_unit_4197(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W36005),
				.b1(W36015),
				.b2(W36025),
				.b3(W36105),
				.b4(W36115),
				.b5(W36125),
				.b6(W36205),
				.b7(W36215),
				.b8(W36225),
				.c(c35226)
);

ninexnine_unit ninexnine_unit_4198(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W36006),
				.b1(W36016),
				.b2(W36026),
				.b3(W36106),
				.b4(W36116),
				.b5(W36126),
				.b6(W36206),
				.b7(W36216),
				.b8(W36226),
				.c(c36226)
);

ninexnine_unit ninexnine_unit_4199(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W36007),
				.b1(W36017),
				.b2(W36027),
				.b3(W36107),
				.b4(W36117),
				.b5(W36127),
				.b6(W36207),
				.b7(W36217),
				.b8(W36227),
				.c(c37226)
);

ninexnine_unit ninexnine_unit_4200(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W36008),
				.b1(W36018),
				.b2(W36028),
				.b3(W36108),
				.b4(W36118),
				.b5(W36128),
				.b6(W36208),
				.b7(W36218),
				.b8(W36228),
				.c(c38226)
);

ninexnine_unit ninexnine_unit_4201(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W36009),
				.b1(W36019),
				.b2(W36029),
				.b3(W36109),
				.b4(W36119),
				.b5(W36129),
				.b6(W36209),
				.b7(W36219),
				.b8(W36229),
				.c(c39226)
);

ninexnine_unit ninexnine_unit_4202(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3600A),
				.b1(W3601A),
				.b2(W3602A),
				.b3(W3610A),
				.b4(W3611A),
				.b5(W3612A),
				.b6(W3620A),
				.b7(W3621A),
				.b8(W3622A),
				.c(c3A226)
);

ninexnine_unit ninexnine_unit_4203(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3600B),
				.b1(W3601B),
				.b2(W3602B),
				.b3(W3610B),
				.b4(W3611B),
				.b5(W3612B),
				.b6(W3620B),
				.b7(W3621B),
				.b8(W3622B),
				.c(c3B226)
);

ninexnine_unit ninexnine_unit_4204(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3600C),
				.b1(W3601C),
				.b2(W3602C),
				.b3(W3610C),
				.b4(W3611C),
				.b5(W3612C),
				.b6(W3620C),
				.b7(W3621C),
				.b8(W3622C),
				.c(c3C226)
);

ninexnine_unit ninexnine_unit_4205(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3600D),
				.b1(W3601D),
				.b2(W3602D),
				.b3(W3610D),
				.b4(W3611D),
				.b5(W3612D),
				.b6(W3620D),
				.b7(W3621D),
				.b8(W3622D),
				.c(c3D226)
);

ninexnine_unit ninexnine_unit_4206(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3600E),
				.b1(W3601E),
				.b2(W3602E),
				.b3(W3610E),
				.b4(W3611E),
				.b5(W3612E),
				.b6(W3620E),
				.b7(W3621E),
				.b8(W3622E),
				.c(c3E226)
);

ninexnine_unit ninexnine_unit_4207(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3600F),
				.b1(W3601F),
				.b2(W3602F),
				.b3(W3610F),
				.b4(W3611F),
				.b5(W3612F),
				.b6(W3620F),
				.b7(W3621F),
				.b8(W3622F),
				.c(c3F226)
);

assign C3226=c30226+c31226+c32226+c33226+c34226+c35226+c36226+c37226+c38226+c39226+c3A226+c3B226+c3C226+c3D226+c3E226+c3F226;
assign A3226=(C3226>=0)?1:0;

assign P4226=A3226;

ninexnine_unit ninexnine_unit_4208(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30007)
);

ninexnine_unit ninexnine_unit_4209(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31007)
);

ninexnine_unit ninexnine_unit_4210(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32007)
);

ninexnine_unit ninexnine_unit_4211(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33007)
);

ninexnine_unit ninexnine_unit_4212(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34007)
);

ninexnine_unit ninexnine_unit_4213(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35007)
);

ninexnine_unit ninexnine_unit_4214(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36007)
);

ninexnine_unit ninexnine_unit_4215(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37007)
);

ninexnine_unit ninexnine_unit_4216(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38007)
);

ninexnine_unit ninexnine_unit_4217(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39007)
);

ninexnine_unit ninexnine_unit_4218(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A007)
);

ninexnine_unit ninexnine_unit_4219(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B007)
);

ninexnine_unit ninexnine_unit_4220(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C007)
);

ninexnine_unit ninexnine_unit_4221(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D007)
);

ninexnine_unit ninexnine_unit_4222(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E007)
);

ninexnine_unit ninexnine_unit_4223(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F007)
);

assign C3007=c30007+c31007+c32007+c33007+c34007+c35007+c36007+c37007+c38007+c39007+c3A007+c3B007+c3C007+c3D007+c3E007+c3F007;
assign A3007=(C3007>=0)?1:0;

assign P4007=A3007;

ninexnine_unit ninexnine_unit_4224(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30017)
);

ninexnine_unit ninexnine_unit_4225(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31017)
);

ninexnine_unit ninexnine_unit_4226(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32017)
);

ninexnine_unit ninexnine_unit_4227(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33017)
);

ninexnine_unit ninexnine_unit_4228(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34017)
);

ninexnine_unit ninexnine_unit_4229(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35017)
);

ninexnine_unit ninexnine_unit_4230(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36017)
);

ninexnine_unit ninexnine_unit_4231(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37017)
);

ninexnine_unit ninexnine_unit_4232(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38017)
);

ninexnine_unit ninexnine_unit_4233(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39017)
);

ninexnine_unit ninexnine_unit_4234(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A017)
);

ninexnine_unit ninexnine_unit_4235(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B017)
);

ninexnine_unit ninexnine_unit_4236(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C017)
);

ninexnine_unit ninexnine_unit_4237(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D017)
);

ninexnine_unit ninexnine_unit_4238(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E017)
);

ninexnine_unit ninexnine_unit_4239(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F017)
);

assign C3017=c30017+c31017+c32017+c33017+c34017+c35017+c36017+c37017+c38017+c39017+c3A017+c3B017+c3C017+c3D017+c3E017+c3F017;
assign A3017=(C3017>=0)?1:0;

assign P4017=A3017;

ninexnine_unit ninexnine_unit_4240(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30027)
);

ninexnine_unit ninexnine_unit_4241(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31027)
);

ninexnine_unit ninexnine_unit_4242(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32027)
);

ninexnine_unit ninexnine_unit_4243(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33027)
);

ninexnine_unit ninexnine_unit_4244(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34027)
);

ninexnine_unit ninexnine_unit_4245(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35027)
);

ninexnine_unit ninexnine_unit_4246(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36027)
);

ninexnine_unit ninexnine_unit_4247(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37027)
);

ninexnine_unit ninexnine_unit_4248(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38027)
);

ninexnine_unit ninexnine_unit_4249(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39027)
);

ninexnine_unit ninexnine_unit_4250(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A027)
);

ninexnine_unit ninexnine_unit_4251(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B027)
);

ninexnine_unit ninexnine_unit_4252(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C027)
);

ninexnine_unit ninexnine_unit_4253(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D027)
);

ninexnine_unit ninexnine_unit_4254(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E027)
);

ninexnine_unit ninexnine_unit_4255(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F027)
);

assign C3027=c30027+c31027+c32027+c33027+c34027+c35027+c36027+c37027+c38027+c39027+c3A027+c3B027+c3C027+c3D027+c3E027+c3F027;
assign A3027=(C3027>=0)?1:0;

assign P4027=A3027;

ninexnine_unit ninexnine_unit_4256(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30107)
);

ninexnine_unit ninexnine_unit_4257(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31107)
);

ninexnine_unit ninexnine_unit_4258(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32107)
);

ninexnine_unit ninexnine_unit_4259(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33107)
);

ninexnine_unit ninexnine_unit_4260(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34107)
);

ninexnine_unit ninexnine_unit_4261(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35107)
);

ninexnine_unit ninexnine_unit_4262(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36107)
);

ninexnine_unit ninexnine_unit_4263(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37107)
);

ninexnine_unit ninexnine_unit_4264(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38107)
);

ninexnine_unit ninexnine_unit_4265(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39107)
);

ninexnine_unit ninexnine_unit_4266(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A107)
);

ninexnine_unit ninexnine_unit_4267(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B107)
);

ninexnine_unit ninexnine_unit_4268(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C107)
);

ninexnine_unit ninexnine_unit_4269(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D107)
);

ninexnine_unit ninexnine_unit_4270(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E107)
);

ninexnine_unit ninexnine_unit_4271(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F107)
);

assign C3107=c30107+c31107+c32107+c33107+c34107+c35107+c36107+c37107+c38107+c39107+c3A107+c3B107+c3C107+c3D107+c3E107+c3F107;
assign A3107=(C3107>=0)?1:0;

assign P4107=A3107;

ninexnine_unit ninexnine_unit_4272(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30117)
);

ninexnine_unit ninexnine_unit_4273(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31117)
);

ninexnine_unit ninexnine_unit_4274(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32117)
);

ninexnine_unit ninexnine_unit_4275(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33117)
);

ninexnine_unit ninexnine_unit_4276(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34117)
);

ninexnine_unit ninexnine_unit_4277(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35117)
);

ninexnine_unit ninexnine_unit_4278(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36117)
);

ninexnine_unit ninexnine_unit_4279(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37117)
);

ninexnine_unit ninexnine_unit_4280(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38117)
);

ninexnine_unit ninexnine_unit_4281(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39117)
);

ninexnine_unit ninexnine_unit_4282(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A117)
);

ninexnine_unit ninexnine_unit_4283(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B117)
);

ninexnine_unit ninexnine_unit_4284(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C117)
);

ninexnine_unit ninexnine_unit_4285(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D117)
);

ninexnine_unit ninexnine_unit_4286(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E117)
);

ninexnine_unit ninexnine_unit_4287(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F117)
);

assign C3117=c30117+c31117+c32117+c33117+c34117+c35117+c36117+c37117+c38117+c39117+c3A117+c3B117+c3C117+c3D117+c3E117+c3F117;
assign A3117=(C3117>=0)?1:0;

assign P4117=A3117;

ninexnine_unit ninexnine_unit_4288(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30127)
);

ninexnine_unit ninexnine_unit_4289(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31127)
);

ninexnine_unit ninexnine_unit_4290(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32127)
);

ninexnine_unit ninexnine_unit_4291(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33127)
);

ninexnine_unit ninexnine_unit_4292(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34127)
);

ninexnine_unit ninexnine_unit_4293(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35127)
);

ninexnine_unit ninexnine_unit_4294(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36127)
);

ninexnine_unit ninexnine_unit_4295(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37127)
);

ninexnine_unit ninexnine_unit_4296(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38127)
);

ninexnine_unit ninexnine_unit_4297(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39127)
);

ninexnine_unit ninexnine_unit_4298(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A127)
);

ninexnine_unit ninexnine_unit_4299(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B127)
);

ninexnine_unit ninexnine_unit_4300(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C127)
);

ninexnine_unit ninexnine_unit_4301(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D127)
);

ninexnine_unit ninexnine_unit_4302(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E127)
);

ninexnine_unit ninexnine_unit_4303(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F127)
);

assign C3127=c30127+c31127+c32127+c33127+c34127+c35127+c36127+c37127+c38127+c39127+c3A127+c3B127+c3C127+c3D127+c3E127+c3F127;
assign A3127=(C3127>=0)?1:0;

assign P4127=A3127;

ninexnine_unit ninexnine_unit_4304(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30207)
);

ninexnine_unit ninexnine_unit_4305(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31207)
);

ninexnine_unit ninexnine_unit_4306(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32207)
);

ninexnine_unit ninexnine_unit_4307(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33207)
);

ninexnine_unit ninexnine_unit_4308(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34207)
);

ninexnine_unit ninexnine_unit_4309(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35207)
);

ninexnine_unit ninexnine_unit_4310(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36207)
);

ninexnine_unit ninexnine_unit_4311(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37207)
);

ninexnine_unit ninexnine_unit_4312(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38207)
);

ninexnine_unit ninexnine_unit_4313(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39207)
);

ninexnine_unit ninexnine_unit_4314(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A207)
);

ninexnine_unit ninexnine_unit_4315(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B207)
);

ninexnine_unit ninexnine_unit_4316(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C207)
);

ninexnine_unit ninexnine_unit_4317(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D207)
);

ninexnine_unit ninexnine_unit_4318(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E207)
);

ninexnine_unit ninexnine_unit_4319(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F207)
);

assign C3207=c30207+c31207+c32207+c33207+c34207+c35207+c36207+c37207+c38207+c39207+c3A207+c3B207+c3C207+c3D207+c3E207+c3F207;
assign A3207=(C3207>=0)?1:0;

assign P4207=A3207;

ninexnine_unit ninexnine_unit_4320(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30217)
);

ninexnine_unit ninexnine_unit_4321(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31217)
);

ninexnine_unit ninexnine_unit_4322(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32217)
);

ninexnine_unit ninexnine_unit_4323(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33217)
);

ninexnine_unit ninexnine_unit_4324(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34217)
);

ninexnine_unit ninexnine_unit_4325(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35217)
);

ninexnine_unit ninexnine_unit_4326(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36217)
);

ninexnine_unit ninexnine_unit_4327(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37217)
);

ninexnine_unit ninexnine_unit_4328(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38217)
);

ninexnine_unit ninexnine_unit_4329(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39217)
);

ninexnine_unit ninexnine_unit_4330(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A217)
);

ninexnine_unit ninexnine_unit_4331(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B217)
);

ninexnine_unit ninexnine_unit_4332(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C217)
);

ninexnine_unit ninexnine_unit_4333(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D217)
);

ninexnine_unit ninexnine_unit_4334(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E217)
);

ninexnine_unit ninexnine_unit_4335(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F217)
);

assign C3217=c30217+c31217+c32217+c33217+c34217+c35217+c36217+c37217+c38217+c39217+c3A217+c3B217+c3C217+c3D217+c3E217+c3F217;
assign A3217=(C3217>=0)?1:0;

assign P4217=A3217;

ninexnine_unit ninexnine_unit_4336(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W37000),
				.b1(W37010),
				.b2(W37020),
				.b3(W37100),
				.b4(W37110),
				.b5(W37120),
				.b6(W37200),
				.b7(W37210),
				.b8(W37220),
				.c(c30227)
);

ninexnine_unit ninexnine_unit_4337(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W37001),
				.b1(W37011),
				.b2(W37021),
				.b3(W37101),
				.b4(W37111),
				.b5(W37121),
				.b6(W37201),
				.b7(W37211),
				.b8(W37221),
				.c(c31227)
);

ninexnine_unit ninexnine_unit_4338(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W37002),
				.b1(W37012),
				.b2(W37022),
				.b3(W37102),
				.b4(W37112),
				.b5(W37122),
				.b6(W37202),
				.b7(W37212),
				.b8(W37222),
				.c(c32227)
);

ninexnine_unit ninexnine_unit_4339(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W37003),
				.b1(W37013),
				.b2(W37023),
				.b3(W37103),
				.b4(W37113),
				.b5(W37123),
				.b6(W37203),
				.b7(W37213),
				.b8(W37223),
				.c(c33227)
);

ninexnine_unit ninexnine_unit_4340(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W37004),
				.b1(W37014),
				.b2(W37024),
				.b3(W37104),
				.b4(W37114),
				.b5(W37124),
				.b6(W37204),
				.b7(W37214),
				.b8(W37224),
				.c(c34227)
);

ninexnine_unit ninexnine_unit_4341(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W37005),
				.b1(W37015),
				.b2(W37025),
				.b3(W37105),
				.b4(W37115),
				.b5(W37125),
				.b6(W37205),
				.b7(W37215),
				.b8(W37225),
				.c(c35227)
);

ninexnine_unit ninexnine_unit_4342(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W37006),
				.b1(W37016),
				.b2(W37026),
				.b3(W37106),
				.b4(W37116),
				.b5(W37126),
				.b6(W37206),
				.b7(W37216),
				.b8(W37226),
				.c(c36227)
);

ninexnine_unit ninexnine_unit_4343(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W37007),
				.b1(W37017),
				.b2(W37027),
				.b3(W37107),
				.b4(W37117),
				.b5(W37127),
				.b6(W37207),
				.b7(W37217),
				.b8(W37227),
				.c(c37227)
);

ninexnine_unit ninexnine_unit_4344(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W37008),
				.b1(W37018),
				.b2(W37028),
				.b3(W37108),
				.b4(W37118),
				.b5(W37128),
				.b6(W37208),
				.b7(W37218),
				.b8(W37228),
				.c(c38227)
);

ninexnine_unit ninexnine_unit_4345(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W37009),
				.b1(W37019),
				.b2(W37029),
				.b3(W37109),
				.b4(W37119),
				.b5(W37129),
				.b6(W37209),
				.b7(W37219),
				.b8(W37229),
				.c(c39227)
);

ninexnine_unit ninexnine_unit_4346(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3700A),
				.b1(W3701A),
				.b2(W3702A),
				.b3(W3710A),
				.b4(W3711A),
				.b5(W3712A),
				.b6(W3720A),
				.b7(W3721A),
				.b8(W3722A),
				.c(c3A227)
);

ninexnine_unit ninexnine_unit_4347(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3700B),
				.b1(W3701B),
				.b2(W3702B),
				.b3(W3710B),
				.b4(W3711B),
				.b5(W3712B),
				.b6(W3720B),
				.b7(W3721B),
				.b8(W3722B),
				.c(c3B227)
);

ninexnine_unit ninexnine_unit_4348(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3700C),
				.b1(W3701C),
				.b2(W3702C),
				.b3(W3710C),
				.b4(W3711C),
				.b5(W3712C),
				.b6(W3720C),
				.b7(W3721C),
				.b8(W3722C),
				.c(c3C227)
);

ninexnine_unit ninexnine_unit_4349(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3700D),
				.b1(W3701D),
				.b2(W3702D),
				.b3(W3710D),
				.b4(W3711D),
				.b5(W3712D),
				.b6(W3720D),
				.b7(W3721D),
				.b8(W3722D),
				.c(c3D227)
);

ninexnine_unit ninexnine_unit_4350(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3700E),
				.b1(W3701E),
				.b2(W3702E),
				.b3(W3710E),
				.b4(W3711E),
				.b5(W3712E),
				.b6(W3720E),
				.b7(W3721E),
				.b8(W3722E),
				.c(c3E227)
);

ninexnine_unit ninexnine_unit_4351(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3700F),
				.b1(W3701F),
				.b2(W3702F),
				.b3(W3710F),
				.b4(W3711F),
				.b5(W3712F),
				.b6(W3720F),
				.b7(W3721F),
				.b8(W3722F),
				.c(c3F227)
);

assign C3227=c30227+c31227+c32227+c33227+c34227+c35227+c36227+c37227+c38227+c39227+c3A227+c3B227+c3C227+c3D227+c3E227+c3F227;
assign A3227=(C3227>=0)?1:0;

assign P4227=A3227;

ninexnine_unit ninexnine_unit_4352(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30008)
);

ninexnine_unit ninexnine_unit_4353(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31008)
);

ninexnine_unit ninexnine_unit_4354(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32008)
);

ninexnine_unit ninexnine_unit_4355(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33008)
);

ninexnine_unit ninexnine_unit_4356(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34008)
);

ninexnine_unit ninexnine_unit_4357(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35008)
);

ninexnine_unit ninexnine_unit_4358(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36008)
);

ninexnine_unit ninexnine_unit_4359(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37008)
);

ninexnine_unit ninexnine_unit_4360(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38008)
);

ninexnine_unit ninexnine_unit_4361(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39008)
);

ninexnine_unit ninexnine_unit_4362(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A008)
);

ninexnine_unit ninexnine_unit_4363(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B008)
);

ninexnine_unit ninexnine_unit_4364(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C008)
);

ninexnine_unit ninexnine_unit_4365(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D008)
);

ninexnine_unit ninexnine_unit_4366(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E008)
);

ninexnine_unit ninexnine_unit_4367(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F008)
);

assign C3008=c30008+c31008+c32008+c33008+c34008+c35008+c36008+c37008+c38008+c39008+c3A008+c3B008+c3C008+c3D008+c3E008+c3F008;
assign A3008=(C3008>=0)?1:0;

assign P4008=A3008;

ninexnine_unit ninexnine_unit_4368(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30018)
);

ninexnine_unit ninexnine_unit_4369(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31018)
);

ninexnine_unit ninexnine_unit_4370(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32018)
);

ninexnine_unit ninexnine_unit_4371(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33018)
);

ninexnine_unit ninexnine_unit_4372(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34018)
);

ninexnine_unit ninexnine_unit_4373(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35018)
);

ninexnine_unit ninexnine_unit_4374(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36018)
);

ninexnine_unit ninexnine_unit_4375(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37018)
);

ninexnine_unit ninexnine_unit_4376(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38018)
);

ninexnine_unit ninexnine_unit_4377(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39018)
);

ninexnine_unit ninexnine_unit_4378(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A018)
);

ninexnine_unit ninexnine_unit_4379(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B018)
);

ninexnine_unit ninexnine_unit_4380(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C018)
);

ninexnine_unit ninexnine_unit_4381(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D018)
);

ninexnine_unit ninexnine_unit_4382(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E018)
);

ninexnine_unit ninexnine_unit_4383(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F018)
);

assign C3018=c30018+c31018+c32018+c33018+c34018+c35018+c36018+c37018+c38018+c39018+c3A018+c3B018+c3C018+c3D018+c3E018+c3F018;
assign A3018=(C3018>=0)?1:0;

assign P4018=A3018;

ninexnine_unit ninexnine_unit_4384(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30028)
);

ninexnine_unit ninexnine_unit_4385(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31028)
);

ninexnine_unit ninexnine_unit_4386(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32028)
);

ninexnine_unit ninexnine_unit_4387(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33028)
);

ninexnine_unit ninexnine_unit_4388(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34028)
);

ninexnine_unit ninexnine_unit_4389(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35028)
);

ninexnine_unit ninexnine_unit_4390(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36028)
);

ninexnine_unit ninexnine_unit_4391(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37028)
);

ninexnine_unit ninexnine_unit_4392(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38028)
);

ninexnine_unit ninexnine_unit_4393(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39028)
);

ninexnine_unit ninexnine_unit_4394(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A028)
);

ninexnine_unit ninexnine_unit_4395(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B028)
);

ninexnine_unit ninexnine_unit_4396(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C028)
);

ninexnine_unit ninexnine_unit_4397(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D028)
);

ninexnine_unit ninexnine_unit_4398(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E028)
);

ninexnine_unit ninexnine_unit_4399(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F028)
);

assign C3028=c30028+c31028+c32028+c33028+c34028+c35028+c36028+c37028+c38028+c39028+c3A028+c3B028+c3C028+c3D028+c3E028+c3F028;
assign A3028=(C3028>=0)?1:0;

assign P4028=A3028;

ninexnine_unit ninexnine_unit_4400(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30108)
);

ninexnine_unit ninexnine_unit_4401(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31108)
);

ninexnine_unit ninexnine_unit_4402(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32108)
);

ninexnine_unit ninexnine_unit_4403(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33108)
);

ninexnine_unit ninexnine_unit_4404(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34108)
);

ninexnine_unit ninexnine_unit_4405(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35108)
);

ninexnine_unit ninexnine_unit_4406(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36108)
);

ninexnine_unit ninexnine_unit_4407(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37108)
);

ninexnine_unit ninexnine_unit_4408(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38108)
);

ninexnine_unit ninexnine_unit_4409(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39108)
);

ninexnine_unit ninexnine_unit_4410(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A108)
);

ninexnine_unit ninexnine_unit_4411(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B108)
);

ninexnine_unit ninexnine_unit_4412(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C108)
);

ninexnine_unit ninexnine_unit_4413(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D108)
);

ninexnine_unit ninexnine_unit_4414(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E108)
);

ninexnine_unit ninexnine_unit_4415(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F108)
);

assign C3108=c30108+c31108+c32108+c33108+c34108+c35108+c36108+c37108+c38108+c39108+c3A108+c3B108+c3C108+c3D108+c3E108+c3F108;
assign A3108=(C3108>=0)?1:0;

assign P4108=A3108;

ninexnine_unit ninexnine_unit_4416(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30118)
);

ninexnine_unit ninexnine_unit_4417(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31118)
);

ninexnine_unit ninexnine_unit_4418(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32118)
);

ninexnine_unit ninexnine_unit_4419(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33118)
);

ninexnine_unit ninexnine_unit_4420(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34118)
);

ninexnine_unit ninexnine_unit_4421(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35118)
);

ninexnine_unit ninexnine_unit_4422(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36118)
);

ninexnine_unit ninexnine_unit_4423(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37118)
);

ninexnine_unit ninexnine_unit_4424(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38118)
);

ninexnine_unit ninexnine_unit_4425(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39118)
);

ninexnine_unit ninexnine_unit_4426(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A118)
);

ninexnine_unit ninexnine_unit_4427(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B118)
);

ninexnine_unit ninexnine_unit_4428(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C118)
);

ninexnine_unit ninexnine_unit_4429(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D118)
);

ninexnine_unit ninexnine_unit_4430(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E118)
);

ninexnine_unit ninexnine_unit_4431(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F118)
);

assign C3118=c30118+c31118+c32118+c33118+c34118+c35118+c36118+c37118+c38118+c39118+c3A118+c3B118+c3C118+c3D118+c3E118+c3F118;
assign A3118=(C3118>=0)?1:0;

assign P4118=A3118;

ninexnine_unit ninexnine_unit_4432(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30128)
);

ninexnine_unit ninexnine_unit_4433(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31128)
);

ninexnine_unit ninexnine_unit_4434(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32128)
);

ninexnine_unit ninexnine_unit_4435(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33128)
);

ninexnine_unit ninexnine_unit_4436(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34128)
);

ninexnine_unit ninexnine_unit_4437(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35128)
);

ninexnine_unit ninexnine_unit_4438(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36128)
);

ninexnine_unit ninexnine_unit_4439(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37128)
);

ninexnine_unit ninexnine_unit_4440(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38128)
);

ninexnine_unit ninexnine_unit_4441(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39128)
);

ninexnine_unit ninexnine_unit_4442(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A128)
);

ninexnine_unit ninexnine_unit_4443(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B128)
);

ninexnine_unit ninexnine_unit_4444(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C128)
);

ninexnine_unit ninexnine_unit_4445(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D128)
);

ninexnine_unit ninexnine_unit_4446(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E128)
);

ninexnine_unit ninexnine_unit_4447(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F128)
);

assign C3128=c30128+c31128+c32128+c33128+c34128+c35128+c36128+c37128+c38128+c39128+c3A128+c3B128+c3C128+c3D128+c3E128+c3F128;
assign A3128=(C3128>=0)?1:0;

assign P4128=A3128;

ninexnine_unit ninexnine_unit_4448(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30208)
);

ninexnine_unit ninexnine_unit_4449(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31208)
);

ninexnine_unit ninexnine_unit_4450(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32208)
);

ninexnine_unit ninexnine_unit_4451(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33208)
);

ninexnine_unit ninexnine_unit_4452(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34208)
);

ninexnine_unit ninexnine_unit_4453(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35208)
);

ninexnine_unit ninexnine_unit_4454(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36208)
);

ninexnine_unit ninexnine_unit_4455(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37208)
);

ninexnine_unit ninexnine_unit_4456(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38208)
);

ninexnine_unit ninexnine_unit_4457(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39208)
);

ninexnine_unit ninexnine_unit_4458(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A208)
);

ninexnine_unit ninexnine_unit_4459(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B208)
);

ninexnine_unit ninexnine_unit_4460(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C208)
);

ninexnine_unit ninexnine_unit_4461(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D208)
);

ninexnine_unit ninexnine_unit_4462(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E208)
);

ninexnine_unit ninexnine_unit_4463(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F208)
);

assign C3208=c30208+c31208+c32208+c33208+c34208+c35208+c36208+c37208+c38208+c39208+c3A208+c3B208+c3C208+c3D208+c3E208+c3F208;
assign A3208=(C3208>=0)?1:0;

assign P4208=A3208;

ninexnine_unit ninexnine_unit_4464(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30218)
);

ninexnine_unit ninexnine_unit_4465(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31218)
);

ninexnine_unit ninexnine_unit_4466(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32218)
);

ninexnine_unit ninexnine_unit_4467(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33218)
);

ninexnine_unit ninexnine_unit_4468(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34218)
);

ninexnine_unit ninexnine_unit_4469(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35218)
);

ninexnine_unit ninexnine_unit_4470(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36218)
);

ninexnine_unit ninexnine_unit_4471(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37218)
);

ninexnine_unit ninexnine_unit_4472(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38218)
);

ninexnine_unit ninexnine_unit_4473(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39218)
);

ninexnine_unit ninexnine_unit_4474(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A218)
);

ninexnine_unit ninexnine_unit_4475(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B218)
);

ninexnine_unit ninexnine_unit_4476(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C218)
);

ninexnine_unit ninexnine_unit_4477(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D218)
);

ninexnine_unit ninexnine_unit_4478(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E218)
);

ninexnine_unit ninexnine_unit_4479(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F218)
);

assign C3218=c30218+c31218+c32218+c33218+c34218+c35218+c36218+c37218+c38218+c39218+c3A218+c3B218+c3C218+c3D218+c3E218+c3F218;
assign A3218=(C3218>=0)?1:0;

assign P4218=A3218;

ninexnine_unit ninexnine_unit_4480(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W38000),
				.b1(W38010),
				.b2(W38020),
				.b3(W38100),
				.b4(W38110),
				.b5(W38120),
				.b6(W38200),
				.b7(W38210),
				.b8(W38220),
				.c(c30228)
);

ninexnine_unit ninexnine_unit_4481(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W38001),
				.b1(W38011),
				.b2(W38021),
				.b3(W38101),
				.b4(W38111),
				.b5(W38121),
				.b6(W38201),
				.b7(W38211),
				.b8(W38221),
				.c(c31228)
);

ninexnine_unit ninexnine_unit_4482(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W38002),
				.b1(W38012),
				.b2(W38022),
				.b3(W38102),
				.b4(W38112),
				.b5(W38122),
				.b6(W38202),
				.b7(W38212),
				.b8(W38222),
				.c(c32228)
);

ninexnine_unit ninexnine_unit_4483(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W38003),
				.b1(W38013),
				.b2(W38023),
				.b3(W38103),
				.b4(W38113),
				.b5(W38123),
				.b6(W38203),
				.b7(W38213),
				.b8(W38223),
				.c(c33228)
);

ninexnine_unit ninexnine_unit_4484(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W38004),
				.b1(W38014),
				.b2(W38024),
				.b3(W38104),
				.b4(W38114),
				.b5(W38124),
				.b6(W38204),
				.b7(W38214),
				.b8(W38224),
				.c(c34228)
);

ninexnine_unit ninexnine_unit_4485(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W38005),
				.b1(W38015),
				.b2(W38025),
				.b3(W38105),
				.b4(W38115),
				.b5(W38125),
				.b6(W38205),
				.b7(W38215),
				.b8(W38225),
				.c(c35228)
);

ninexnine_unit ninexnine_unit_4486(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W38006),
				.b1(W38016),
				.b2(W38026),
				.b3(W38106),
				.b4(W38116),
				.b5(W38126),
				.b6(W38206),
				.b7(W38216),
				.b8(W38226),
				.c(c36228)
);

ninexnine_unit ninexnine_unit_4487(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W38007),
				.b1(W38017),
				.b2(W38027),
				.b3(W38107),
				.b4(W38117),
				.b5(W38127),
				.b6(W38207),
				.b7(W38217),
				.b8(W38227),
				.c(c37228)
);

ninexnine_unit ninexnine_unit_4488(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W38008),
				.b1(W38018),
				.b2(W38028),
				.b3(W38108),
				.b4(W38118),
				.b5(W38128),
				.b6(W38208),
				.b7(W38218),
				.b8(W38228),
				.c(c38228)
);

ninexnine_unit ninexnine_unit_4489(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W38009),
				.b1(W38019),
				.b2(W38029),
				.b3(W38109),
				.b4(W38119),
				.b5(W38129),
				.b6(W38209),
				.b7(W38219),
				.b8(W38229),
				.c(c39228)
);

ninexnine_unit ninexnine_unit_4490(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3800A),
				.b1(W3801A),
				.b2(W3802A),
				.b3(W3810A),
				.b4(W3811A),
				.b5(W3812A),
				.b6(W3820A),
				.b7(W3821A),
				.b8(W3822A),
				.c(c3A228)
);

ninexnine_unit ninexnine_unit_4491(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3800B),
				.b1(W3801B),
				.b2(W3802B),
				.b3(W3810B),
				.b4(W3811B),
				.b5(W3812B),
				.b6(W3820B),
				.b7(W3821B),
				.b8(W3822B),
				.c(c3B228)
);

ninexnine_unit ninexnine_unit_4492(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3800C),
				.b1(W3801C),
				.b2(W3802C),
				.b3(W3810C),
				.b4(W3811C),
				.b5(W3812C),
				.b6(W3820C),
				.b7(W3821C),
				.b8(W3822C),
				.c(c3C228)
);

ninexnine_unit ninexnine_unit_4493(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3800D),
				.b1(W3801D),
				.b2(W3802D),
				.b3(W3810D),
				.b4(W3811D),
				.b5(W3812D),
				.b6(W3820D),
				.b7(W3821D),
				.b8(W3822D),
				.c(c3D228)
);

ninexnine_unit ninexnine_unit_4494(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3800E),
				.b1(W3801E),
				.b2(W3802E),
				.b3(W3810E),
				.b4(W3811E),
				.b5(W3812E),
				.b6(W3820E),
				.b7(W3821E),
				.b8(W3822E),
				.c(c3E228)
);

ninexnine_unit ninexnine_unit_4495(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3800F),
				.b1(W3801F),
				.b2(W3802F),
				.b3(W3810F),
				.b4(W3811F),
				.b5(W3812F),
				.b6(W3820F),
				.b7(W3821F),
				.b8(W3822F),
				.c(c3F228)
);

assign C3228=c30228+c31228+c32228+c33228+c34228+c35228+c36228+c37228+c38228+c39228+c3A228+c3B228+c3C228+c3D228+c3E228+c3F228;
assign A3228=(C3228>=0)?1:0;

assign P4228=A3228;

ninexnine_unit ninexnine_unit_4496(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30009)
);

ninexnine_unit ninexnine_unit_4497(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31009)
);

ninexnine_unit ninexnine_unit_4498(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32009)
);

ninexnine_unit ninexnine_unit_4499(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33009)
);

ninexnine_unit ninexnine_unit_4500(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34009)
);

ninexnine_unit ninexnine_unit_4501(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35009)
);

ninexnine_unit ninexnine_unit_4502(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36009)
);

ninexnine_unit ninexnine_unit_4503(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37009)
);

ninexnine_unit ninexnine_unit_4504(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38009)
);

ninexnine_unit ninexnine_unit_4505(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39009)
);

ninexnine_unit ninexnine_unit_4506(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A009)
);

ninexnine_unit ninexnine_unit_4507(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B009)
);

ninexnine_unit ninexnine_unit_4508(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C009)
);

ninexnine_unit ninexnine_unit_4509(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D009)
);

ninexnine_unit ninexnine_unit_4510(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E009)
);

ninexnine_unit ninexnine_unit_4511(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F009)
);

assign C3009=c30009+c31009+c32009+c33009+c34009+c35009+c36009+c37009+c38009+c39009+c3A009+c3B009+c3C009+c3D009+c3E009+c3F009;
assign A3009=(C3009>=0)?1:0;

assign P4009=A3009;

ninexnine_unit ninexnine_unit_4512(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30019)
);

ninexnine_unit ninexnine_unit_4513(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31019)
);

ninexnine_unit ninexnine_unit_4514(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32019)
);

ninexnine_unit ninexnine_unit_4515(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33019)
);

ninexnine_unit ninexnine_unit_4516(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34019)
);

ninexnine_unit ninexnine_unit_4517(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35019)
);

ninexnine_unit ninexnine_unit_4518(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36019)
);

ninexnine_unit ninexnine_unit_4519(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37019)
);

ninexnine_unit ninexnine_unit_4520(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38019)
);

ninexnine_unit ninexnine_unit_4521(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39019)
);

ninexnine_unit ninexnine_unit_4522(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A019)
);

ninexnine_unit ninexnine_unit_4523(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B019)
);

ninexnine_unit ninexnine_unit_4524(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C019)
);

ninexnine_unit ninexnine_unit_4525(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D019)
);

ninexnine_unit ninexnine_unit_4526(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E019)
);

ninexnine_unit ninexnine_unit_4527(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F019)
);

assign C3019=c30019+c31019+c32019+c33019+c34019+c35019+c36019+c37019+c38019+c39019+c3A019+c3B019+c3C019+c3D019+c3E019+c3F019;
assign A3019=(C3019>=0)?1:0;

assign P4019=A3019;

ninexnine_unit ninexnine_unit_4528(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30029)
);

ninexnine_unit ninexnine_unit_4529(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31029)
);

ninexnine_unit ninexnine_unit_4530(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32029)
);

ninexnine_unit ninexnine_unit_4531(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33029)
);

ninexnine_unit ninexnine_unit_4532(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34029)
);

ninexnine_unit ninexnine_unit_4533(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35029)
);

ninexnine_unit ninexnine_unit_4534(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36029)
);

ninexnine_unit ninexnine_unit_4535(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37029)
);

ninexnine_unit ninexnine_unit_4536(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38029)
);

ninexnine_unit ninexnine_unit_4537(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39029)
);

ninexnine_unit ninexnine_unit_4538(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A029)
);

ninexnine_unit ninexnine_unit_4539(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B029)
);

ninexnine_unit ninexnine_unit_4540(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C029)
);

ninexnine_unit ninexnine_unit_4541(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D029)
);

ninexnine_unit ninexnine_unit_4542(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E029)
);

ninexnine_unit ninexnine_unit_4543(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F029)
);

assign C3029=c30029+c31029+c32029+c33029+c34029+c35029+c36029+c37029+c38029+c39029+c3A029+c3B029+c3C029+c3D029+c3E029+c3F029;
assign A3029=(C3029>=0)?1:0;

assign P4029=A3029;

ninexnine_unit ninexnine_unit_4544(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30109)
);

ninexnine_unit ninexnine_unit_4545(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31109)
);

ninexnine_unit ninexnine_unit_4546(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32109)
);

ninexnine_unit ninexnine_unit_4547(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33109)
);

ninexnine_unit ninexnine_unit_4548(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34109)
);

ninexnine_unit ninexnine_unit_4549(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35109)
);

ninexnine_unit ninexnine_unit_4550(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36109)
);

ninexnine_unit ninexnine_unit_4551(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37109)
);

ninexnine_unit ninexnine_unit_4552(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38109)
);

ninexnine_unit ninexnine_unit_4553(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39109)
);

ninexnine_unit ninexnine_unit_4554(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A109)
);

ninexnine_unit ninexnine_unit_4555(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B109)
);

ninexnine_unit ninexnine_unit_4556(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C109)
);

ninexnine_unit ninexnine_unit_4557(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D109)
);

ninexnine_unit ninexnine_unit_4558(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E109)
);

ninexnine_unit ninexnine_unit_4559(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F109)
);

assign C3109=c30109+c31109+c32109+c33109+c34109+c35109+c36109+c37109+c38109+c39109+c3A109+c3B109+c3C109+c3D109+c3E109+c3F109;
assign A3109=(C3109>=0)?1:0;

assign P4109=A3109;

ninexnine_unit ninexnine_unit_4560(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30119)
);

ninexnine_unit ninexnine_unit_4561(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31119)
);

ninexnine_unit ninexnine_unit_4562(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32119)
);

ninexnine_unit ninexnine_unit_4563(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33119)
);

ninexnine_unit ninexnine_unit_4564(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34119)
);

ninexnine_unit ninexnine_unit_4565(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35119)
);

ninexnine_unit ninexnine_unit_4566(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36119)
);

ninexnine_unit ninexnine_unit_4567(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37119)
);

ninexnine_unit ninexnine_unit_4568(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38119)
);

ninexnine_unit ninexnine_unit_4569(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39119)
);

ninexnine_unit ninexnine_unit_4570(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A119)
);

ninexnine_unit ninexnine_unit_4571(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B119)
);

ninexnine_unit ninexnine_unit_4572(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C119)
);

ninexnine_unit ninexnine_unit_4573(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D119)
);

ninexnine_unit ninexnine_unit_4574(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E119)
);

ninexnine_unit ninexnine_unit_4575(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F119)
);

assign C3119=c30119+c31119+c32119+c33119+c34119+c35119+c36119+c37119+c38119+c39119+c3A119+c3B119+c3C119+c3D119+c3E119+c3F119;
assign A3119=(C3119>=0)?1:0;

assign P4119=A3119;

ninexnine_unit ninexnine_unit_4576(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30129)
);

ninexnine_unit ninexnine_unit_4577(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31129)
);

ninexnine_unit ninexnine_unit_4578(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32129)
);

ninexnine_unit ninexnine_unit_4579(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33129)
);

ninexnine_unit ninexnine_unit_4580(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34129)
);

ninexnine_unit ninexnine_unit_4581(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35129)
);

ninexnine_unit ninexnine_unit_4582(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36129)
);

ninexnine_unit ninexnine_unit_4583(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37129)
);

ninexnine_unit ninexnine_unit_4584(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38129)
);

ninexnine_unit ninexnine_unit_4585(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39129)
);

ninexnine_unit ninexnine_unit_4586(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A129)
);

ninexnine_unit ninexnine_unit_4587(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B129)
);

ninexnine_unit ninexnine_unit_4588(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C129)
);

ninexnine_unit ninexnine_unit_4589(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D129)
);

ninexnine_unit ninexnine_unit_4590(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E129)
);

ninexnine_unit ninexnine_unit_4591(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F129)
);

assign C3129=c30129+c31129+c32129+c33129+c34129+c35129+c36129+c37129+c38129+c39129+c3A129+c3B129+c3C129+c3D129+c3E129+c3F129;
assign A3129=(C3129>=0)?1:0;

assign P4129=A3129;

ninexnine_unit ninexnine_unit_4592(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30209)
);

ninexnine_unit ninexnine_unit_4593(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31209)
);

ninexnine_unit ninexnine_unit_4594(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32209)
);

ninexnine_unit ninexnine_unit_4595(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33209)
);

ninexnine_unit ninexnine_unit_4596(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34209)
);

ninexnine_unit ninexnine_unit_4597(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35209)
);

ninexnine_unit ninexnine_unit_4598(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36209)
);

ninexnine_unit ninexnine_unit_4599(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37209)
);

ninexnine_unit ninexnine_unit_4600(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38209)
);

ninexnine_unit ninexnine_unit_4601(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39209)
);

ninexnine_unit ninexnine_unit_4602(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A209)
);

ninexnine_unit ninexnine_unit_4603(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B209)
);

ninexnine_unit ninexnine_unit_4604(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C209)
);

ninexnine_unit ninexnine_unit_4605(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D209)
);

ninexnine_unit ninexnine_unit_4606(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E209)
);

ninexnine_unit ninexnine_unit_4607(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F209)
);

assign C3209=c30209+c31209+c32209+c33209+c34209+c35209+c36209+c37209+c38209+c39209+c3A209+c3B209+c3C209+c3D209+c3E209+c3F209;
assign A3209=(C3209>=0)?1:0;

assign P4209=A3209;

ninexnine_unit ninexnine_unit_4608(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30219)
);

ninexnine_unit ninexnine_unit_4609(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31219)
);

ninexnine_unit ninexnine_unit_4610(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32219)
);

ninexnine_unit ninexnine_unit_4611(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33219)
);

ninexnine_unit ninexnine_unit_4612(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34219)
);

ninexnine_unit ninexnine_unit_4613(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35219)
);

ninexnine_unit ninexnine_unit_4614(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36219)
);

ninexnine_unit ninexnine_unit_4615(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37219)
);

ninexnine_unit ninexnine_unit_4616(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38219)
);

ninexnine_unit ninexnine_unit_4617(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39219)
);

ninexnine_unit ninexnine_unit_4618(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A219)
);

ninexnine_unit ninexnine_unit_4619(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B219)
);

ninexnine_unit ninexnine_unit_4620(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C219)
);

ninexnine_unit ninexnine_unit_4621(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D219)
);

ninexnine_unit ninexnine_unit_4622(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E219)
);

ninexnine_unit ninexnine_unit_4623(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F219)
);

assign C3219=c30219+c31219+c32219+c33219+c34219+c35219+c36219+c37219+c38219+c39219+c3A219+c3B219+c3C219+c3D219+c3E219+c3F219;
assign A3219=(C3219>=0)?1:0;

assign P4219=A3219;

ninexnine_unit ninexnine_unit_4624(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W39000),
				.b1(W39010),
				.b2(W39020),
				.b3(W39100),
				.b4(W39110),
				.b5(W39120),
				.b6(W39200),
				.b7(W39210),
				.b8(W39220),
				.c(c30229)
);

ninexnine_unit ninexnine_unit_4625(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W39001),
				.b1(W39011),
				.b2(W39021),
				.b3(W39101),
				.b4(W39111),
				.b5(W39121),
				.b6(W39201),
				.b7(W39211),
				.b8(W39221),
				.c(c31229)
);

ninexnine_unit ninexnine_unit_4626(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W39002),
				.b1(W39012),
				.b2(W39022),
				.b3(W39102),
				.b4(W39112),
				.b5(W39122),
				.b6(W39202),
				.b7(W39212),
				.b8(W39222),
				.c(c32229)
);

ninexnine_unit ninexnine_unit_4627(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W39003),
				.b1(W39013),
				.b2(W39023),
				.b3(W39103),
				.b4(W39113),
				.b5(W39123),
				.b6(W39203),
				.b7(W39213),
				.b8(W39223),
				.c(c33229)
);

ninexnine_unit ninexnine_unit_4628(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W39004),
				.b1(W39014),
				.b2(W39024),
				.b3(W39104),
				.b4(W39114),
				.b5(W39124),
				.b6(W39204),
				.b7(W39214),
				.b8(W39224),
				.c(c34229)
);

ninexnine_unit ninexnine_unit_4629(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W39005),
				.b1(W39015),
				.b2(W39025),
				.b3(W39105),
				.b4(W39115),
				.b5(W39125),
				.b6(W39205),
				.b7(W39215),
				.b8(W39225),
				.c(c35229)
);

ninexnine_unit ninexnine_unit_4630(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W39006),
				.b1(W39016),
				.b2(W39026),
				.b3(W39106),
				.b4(W39116),
				.b5(W39126),
				.b6(W39206),
				.b7(W39216),
				.b8(W39226),
				.c(c36229)
);

ninexnine_unit ninexnine_unit_4631(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W39007),
				.b1(W39017),
				.b2(W39027),
				.b3(W39107),
				.b4(W39117),
				.b5(W39127),
				.b6(W39207),
				.b7(W39217),
				.b8(W39227),
				.c(c37229)
);

ninexnine_unit ninexnine_unit_4632(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W39008),
				.b1(W39018),
				.b2(W39028),
				.b3(W39108),
				.b4(W39118),
				.b5(W39128),
				.b6(W39208),
				.b7(W39218),
				.b8(W39228),
				.c(c38229)
);

ninexnine_unit ninexnine_unit_4633(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W39009),
				.b1(W39019),
				.b2(W39029),
				.b3(W39109),
				.b4(W39119),
				.b5(W39129),
				.b6(W39209),
				.b7(W39219),
				.b8(W39229),
				.c(c39229)
);

ninexnine_unit ninexnine_unit_4634(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3900A),
				.b1(W3901A),
				.b2(W3902A),
				.b3(W3910A),
				.b4(W3911A),
				.b5(W3912A),
				.b6(W3920A),
				.b7(W3921A),
				.b8(W3922A),
				.c(c3A229)
);

ninexnine_unit ninexnine_unit_4635(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3900B),
				.b1(W3901B),
				.b2(W3902B),
				.b3(W3910B),
				.b4(W3911B),
				.b5(W3912B),
				.b6(W3920B),
				.b7(W3921B),
				.b8(W3922B),
				.c(c3B229)
);

ninexnine_unit ninexnine_unit_4636(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3900C),
				.b1(W3901C),
				.b2(W3902C),
				.b3(W3910C),
				.b4(W3911C),
				.b5(W3912C),
				.b6(W3920C),
				.b7(W3921C),
				.b8(W3922C),
				.c(c3C229)
);

ninexnine_unit ninexnine_unit_4637(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3900D),
				.b1(W3901D),
				.b2(W3902D),
				.b3(W3910D),
				.b4(W3911D),
				.b5(W3912D),
				.b6(W3920D),
				.b7(W3921D),
				.b8(W3922D),
				.c(c3D229)
);

ninexnine_unit ninexnine_unit_4638(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3900E),
				.b1(W3901E),
				.b2(W3902E),
				.b3(W3910E),
				.b4(W3911E),
				.b5(W3912E),
				.b6(W3920E),
				.b7(W3921E),
				.b8(W3922E),
				.c(c3E229)
);

ninexnine_unit ninexnine_unit_4639(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3900F),
				.b1(W3901F),
				.b2(W3902F),
				.b3(W3910F),
				.b4(W3911F),
				.b5(W3912F),
				.b6(W3920F),
				.b7(W3921F),
				.b8(W3922F),
				.c(c3F229)
);

assign C3229=c30229+c31229+c32229+c33229+c34229+c35229+c36229+c37229+c38229+c39229+c3A229+c3B229+c3C229+c3D229+c3E229+c3F229;
assign A3229=(C3229>=0)?1:0;

assign P4229=A3229;

ninexnine_unit ninexnine_unit_4640(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3000A)
);

ninexnine_unit ninexnine_unit_4641(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3100A)
);

ninexnine_unit ninexnine_unit_4642(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3200A)
);

ninexnine_unit ninexnine_unit_4643(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3300A)
);

ninexnine_unit ninexnine_unit_4644(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3400A)
);

ninexnine_unit ninexnine_unit_4645(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3500A)
);

ninexnine_unit ninexnine_unit_4646(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3600A)
);

ninexnine_unit ninexnine_unit_4647(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3700A)
);

ninexnine_unit ninexnine_unit_4648(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3800A)
);

ninexnine_unit ninexnine_unit_4649(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3900A)
);

ninexnine_unit ninexnine_unit_4650(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A00A)
);

ninexnine_unit ninexnine_unit_4651(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B00A)
);

ninexnine_unit ninexnine_unit_4652(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C00A)
);

ninexnine_unit ninexnine_unit_4653(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D00A)
);

ninexnine_unit ninexnine_unit_4654(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E00A)
);

ninexnine_unit ninexnine_unit_4655(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F00A)
);

assign C300A=c3000A+c3100A+c3200A+c3300A+c3400A+c3500A+c3600A+c3700A+c3800A+c3900A+c3A00A+c3B00A+c3C00A+c3D00A+c3E00A+c3F00A;
assign A300A=(C300A>=0)?1:0;

assign P400A=A300A;

ninexnine_unit ninexnine_unit_4656(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3001A)
);

ninexnine_unit ninexnine_unit_4657(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3101A)
);

ninexnine_unit ninexnine_unit_4658(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3201A)
);

ninexnine_unit ninexnine_unit_4659(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3301A)
);

ninexnine_unit ninexnine_unit_4660(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3401A)
);

ninexnine_unit ninexnine_unit_4661(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3501A)
);

ninexnine_unit ninexnine_unit_4662(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3601A)
);

ninexnine_unit ninexnine_unit_4663(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3701A)
);

ninexnine_unit ninexnine_unit_4664(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3801A)
);

ninexnine_unit ninexnine_unit_4665(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3901A)
);

ninexnine_unit ninexnine_unit_4666(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A01A)
);

ninexnine_unit ninexnine_unit_4667(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B01A)
);

ninexnine_unit ninexnine_unit_4668(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C01A)
);

ninexnine_unit ninexnine_unit_4669(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D01A)
);

ninexnine_unit ninexnine_unit_4670(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E01A)
);

ninexnine_unit ninexnine_unit_4671(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F01A)
);

assign C301A=c3001A+c3101A+c3201A+c3301A+c3401A+c3501A+c3601A+c3701A+c3801A+c3901A+c3A01A+c3B01A+c3C01A+c3D01A+c3E01A+c3F01A;
assign A301A=(C301A>=0)?1:0;

assign P401A=A301A;

ninexnine_unit ninexnine_unit_4672(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3002A)
);

ninexnine_unit ninexnine_unit_4673(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3102A)
);

ninexnine_unit ninexnine_unit_4674(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3202A)
);

ninexnine_unit ninexnine_unit_4675(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3302A)
);

ninexnine_unit ninexnine_unit_4676(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3402A)
);

ninexnine_unit ninexnine_unit_4677(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3502A)
);

ninexnine_unit ninexnine_unit_4678(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3602A)
);

ninexnine_unit ninexnine_unit_4679(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3702A)
);

ninexnine_unit ninexnine_unit_4680(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3802A)
);

ninexnine_unit ninexnine_unit_4681(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3902A)
);

ninexnine_unit ninexnine_unit_4682(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A02A)
);

ninexnine_unit ninexnine_unit_4683(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B02A)
);

ninexnine_unit ninexnine_unit_4684(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C02A)
);

ninexnine_unit ninexnine_unit_4685(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D02A)
);

ninexnine_unit ninexnine_unit_4686(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E02A)
);

ninexnine_unit ninexnine_unit_4687(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F02A)
);

assign C302A=c3002A+c3102A+c3202A+c3302A+c3402A+c3502A+c3602A+c3702A+c3802A+c3902A+c3A02A+c3B02A+c3C02A+c3D02A+c3E02A+c3F02A;
assign A302A=(C302A>=0)?1:0;

assign P402A=A302A;

ninexnine_unit ninexnine_unit_4688(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3010A)
);

ninexnine_unit ninexnine_unit_4689(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3110A)
);

ninexnine_unit ninexnine_unit_4690(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3210A)
);

ninexnine_unit ninexnine_unit_4691(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3310A)
);

ninexnine_unit ninexnine_unit_4692(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3410A)
);

ninexnine_unit ninexnine_unit_4693(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3510A)
);

ninexnine_unit ninexnine_unit_4694(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3610A)
);

ninexnine_unit ninexnine_unit_4695(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3710A)
);

ninexnine_unit ninexnine_unit_4696(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3810A)
);

ninexnine_unit ninexnine_unit_4697(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3910A)
);

ninexnine_unit ninexnine_unit_4698(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A10A)
);

ninexnine_unit ninexnine_unit_4699(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B10A)
);

ninexnine_unit ninexnine_unit_4700(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C10A)
);

ninexnine_unit ninexnine_unit_4701(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D10A)
);

ninexnine_unit ninexnine_unit_4702(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E10A)
);

ninexnine_unit ninexnine_unit_4703(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F10A)
);

assign C310A=c3010A+c3110A+c3210A+c3310A+c3410A+c3510A+c3610A+c3710A+c3810A+c3910A+c3A10A+c3B10A+c3C10A+c3D10A+c3E10A+c3F10A;
assign A310A=(C310A>=0)?1:0;

assign P410A=A310A;

ninexnine_unit ninexnine_unit_4704(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3011A)
);

ninexnine_unit ninexnine_unit_4705(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3111A)
);

ninexnine_unit ninexnine_unit_4706(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3211A)
);

ninexnine_unit ninexnine_unit_4707(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3311A)
);

ninexnine_unit ninexnine_unit_4708(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3411A)
);

ninexnine_unit ninexnine_unit_4709(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3511A)
);

ninexnine_unit ninexnine_unit_4710(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3611A)
);

ninexnine_unit ninexnine_unit_4711(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3711A)
);

ninexnine_unit ninexnine_unit_4712(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3811A)
);

ninexnine_unit ninexnine_unit_4713(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3911A)
);

ninexnine_unit ninexnine_unit_4714(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A11A)
);

ninexnine_unit ninexnine_unit_4715(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B11A)
);

ninexnine_unit ninexnine_unit_4716(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C11A)
);

ninexnine_unit ninexnine_unit_4717(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D11A)
);

ninexnine_unit ninexnine_unit_4718(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E11A)
);

ninexnine_unit ninexnine_unit_4719(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F11A)
);

assign C311A=c3011A+c3111A+c3211A+c3311A+c3411A+c3511A+c3611A+c3711A+c3811A+c3911A+c3A11A+c3B11A+c3C11A+c3D11A+c3E11A+c3F11A;
assign A311A=(C311A>=0)?1:0;

assign P411A=A311A;

ninexnine_unit ninexnine_unit_4720(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3012A)
);

ninexnine_unit ninexnine_unit_4721(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3112A)
);

ninexnine_unit ninexnine_unit_4722(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3212A)
);

ninexnine_unit ninexnine_unit_4723(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3312A)
);

ninexnine_unit ninexnine_unit_4724(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3412A)
);

ninexnine_unit ninexnine_unit_4725(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3512A)
);

ninexnine_unit ninexnine_unit_4726(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3612A)
);

ninexnine_unit ninexnine_unit_4727(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3712A)
);

ninexnine_unit ninexnine_unit_4728(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3812A)
);

ninexnine_unit ninexnine_unit_4729(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3912A)
);

ninexnine_unit ninexnine_unit_4730(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A12A)
);

ninexnine_unit ninexnine_unit_4731(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B12A)
);

ninexnine_unit ninexnine_unit_4732(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C12A)
);

ninexnine_unit ninexnine_unit_4733(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D12A)
);

ninexnine_unit ninexnine_unit_4734(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E12A)
);

ninexnine_unit ninexnine_unit_4735(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F12A)
);

assign C312A=c3012A+c3112A+c3212A+c3312A+c3412A+c3512A+c3612A+c3712A+c3812A+c3912A+c3A12A+c3B12A+c3C12A+c3D12A+c3E12A+c3F12A;
assign A312A=(C312A>=0)?1:0;

assign P412A=A312A;

ninexnine_unit ninexnine_unit_4736(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3020A)
);

ninexnine_unit ninexnine_unit_4737(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3120A)
);

ninexnine_unit ninexnine_unit_4738(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3220A)
);

ninexnine_unit ninexnine_unit_4739(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3320A)
);

ninexnine_unit ninexnine_unit_4740(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3420A)
);

ninexnine_unit ninexnine_unit_4741(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3520A)
);

ninexnine_unit ninexnine_unit_4742(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3620A)
);

ninexnine_unit ninexnine_unit_4743(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3720A)
);

ninexnine_unit ninexnine_unit_4744(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3820A)
);

ninexnine_unit ninexnine_unit_4745(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3920A)
);

ninexnine_unit ninexnine_unit_4746(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A20A)
);

ninexnine_unit ninexnine_unit_4747(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B20A)
);

ninexnine_unit ninexnine_unit_4748(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C20A)
);

ninexnine_unit ninexnine_unit_4749(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D20A)
);

ninexnine_unit ninexnine_unit_4750(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E20A)
);

ninexnine_unit ninexnine_unit_4751(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F20A)
);

assign C320A=c3020A+c3120A+c3220A+c3320A+c3420A+c3520A+c3620A+c3720A+c3820A+c3920A+c3A20A+c3B20A+c3C20A+c3D20A+c3E20A+c3F20A;
assign A320A=(C320A>=0)?1:0;

assign P420A=A320A;

ninexnine_unit ninexnine_unit_4752(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3021A)
);

ninexnine_unit ninexnine_unit_4753(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3121A)
);

ninexnine_unit ninexnine_unit_4754(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3221A)
);

ninexnine_unit ninexnine_unit_4755(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3321A)
);

ninexnine_unit ninexnine_unit_4756(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3421A)
);

ninexnine_unit ninexnine_unit_4757(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3521A)
);

ninexnine_unit ninexnine_unit_4758(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3621A)
);

ninexnine_unit ninexnine_unit_4759(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3721A)
);

ninexnine_unit ninexnine_unit_4760(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3821A)
);

ninexnine_unit ninexnine_unit_4761(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3921A)
);

ninexnine_unit ninexnine_unit_4762(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A21A)
);

ninexnine_unit ninexnine_unit_4763(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B21A)
);

ninexnine_unit ninexnine_unit_4764(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C21A)
);

ninexnine_unit ninexnine_unit_4765(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D21A)
);

ninexnine_unit ninexnine_unit_4766(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E21A)
);

ninexnine_unit ninexnine_unit_4767(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F21A)
);

assign C321A=c3021A+c3121A+c3221A+c3321A+c3421A+c3521A+c3621A+c3721A+c3821A+c3921A+c3A21A+c3B21A+c3C21A+c3D21A+c3E21A+c3F21A;
assign A321A=(C321A>=0)?1:0;

assign P421A=A321A;

ninexnine_unit ninexnine_unit_4768(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3A000),
				.b1(W3A010),
				.b2(W3A020),
				.b3(W3A100),
				.b4(W3A110),
				.b5(W3A120),
				.b6(W3A200),
				.b7(W3A210),
				.b8(W3A220),
				.c(c3022A)
);

ninexnine_unit ninexnine_unit_4769(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3A001),
				.b1(W3A011),
				.b2(W3A021),
				.b3(W3A101),
				.b4(W3A111),
				.b5(W3A121),
				.b6(W3A201),
				.b7(W3A211),
				.b8(W3A221),
				.c(c3122A)
);

ninexnine_unit ninexnine_unit_4770(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3A002),
				.b1(W3A012),
				.b2(W3A022),
				.b3(W3A102),
				.b4(W3A112),
				.b5(W3A122),
				.b6(W3A202),
				.b7(W3A212),
				.b8(W3A222),
				.c(c3222A)
);

ninexnine_unit ninexnine_unit_4771(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3A003),
				.b1(W3A013),
				.b2(W3A023),
				.b3(W3A103),
				.b4(W3A113),
				.b5(W3A123),
				.b6(W3A203),
				.b7(W3A213),
				.b8(W3A223),
				.c(c3322A)
);

ninexnine_unit ninexnine_unit_4772(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3A004),
				.b1(W3A014),
				.b2(W3A024),
				.b3(W3A104),
				.b4(W3A114),
				.b5(W3A124),
				.b6(W3A204),
				.b7(W3A214),
				.b8(W3A224),
				.c(c3422A)
);

ninexnine_unit ninexnine_unit_4773(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3A005),
				.b1(W3A015),
				.b2(W3A025),
				.b3(W3A105),
				.b4(W3A115),
				.b5(W3A125),
				.b6(W3A205),
				.b7(W3A215),
				.b8(W3A225),
				.c(c3522A)
);

ninexnine_unit ninexnine_unit_4774(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3A006),
				.b1(W3A016),
				.b2(W3A026),
				.b3(W3A106),
				.b4(W3A116),
				.b5(W3A126),
				.b6(W3A206),
				.b7(W3A216),
				.b8(W3A226),
				.c(c3622A)
);

ninexnine_unit ninexnine_unit_4775(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3A007),
				.b1(W3A017),
				.b2(W3A027),
				.b3(W3A107),
				.b4(W3A117),
				.b5(W3A127),
				.b6(W3A207),
				.b7(W3A217),
				.b8(W3A227),
				.c(c3722A)
);

ninexnine_unit ninexnine_unit_4776(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3A008),
				.b1(W3A018),
				.b2(W3A028),
				.b3(W3A108),
				.b4(W3A118),
				.b5(W3A128),
				.b6(W3A208),
				.b7(W3A218),
				.b8(W3A228),
				.c(c3822A)
);

ninexnine_unit ninexnine_unit_4777(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3A009),
				.b1(W3A019),
				.b2(W3A029),
				.b3(W3A109),
				.b4(W3A119),
				.b5(W3A129),
				.b6(W3A209),
				.b7(W3A219),
				.b8(W3A229),
				.c(c3922A)
);

ninexnine_unit ninexnine_unit_4778(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3A00A),
				.b1(W3A01A),
				.b2(W3A02A),
				.b3(W3A10A),
				.b4(W3A11A),
				.b5(W3A12A),
				.b6(W3A20A),
				.b7(W3A21A),
				.b8(W3A22A),
				.c(c3A22A)
);

ninexnine_unit ninexnine_unit_4779(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3A00B),
				.b1(W3A01B),
				.b2(W3A02B),
				.b3(W3A10B),
				.b4(W3A11B),
				.b5(W3A12B),
				.b6(W3A20B),
				.b7(W3A21B),
				.b8(W3A22B),
				.c(c3B22A)
);

ninexnine_unit ninexnine_unit_4780(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3A00C),
				.b1(W3A01C),
				.b2(W3A02C),
				.b3(W3A10C),
				.b4(W3A11C),
				.b5(W3A12C),
				.b6(W3A20C),
				.b7(W3A21C),
				.b8(W3A22C),
				.c(c3C22A)
);

ninexnine_unit ninexnine_unit_4781(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3A00D),
				.b1(W3A01D),
				.b2(W3A02D),
				.b3(W3A10D),
				.b4(W3A11D),
				.b5(W3A12D),
				.b6(W3A20D),
				.b7(W3A21D),
				.b8(W3A22D),
				.c(c3D22A)
);

ninexnine_unit ninexnine_unit_4782(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3A00E),
				.b1(W3A01E),
				.b2(W3A02E),
				.b3(W3A10E),
				.b4(W3A11E),
				.b5(W3A12E),
				.b6(W3A20E),
				.b7(W3A21E),
				.b8(W3A22E),
				.c(c3E22A)
);

ninexnine_unit ninexnine_unit_4783(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3A00F),
				.b1(W3A01F),
				.b2(W3A02F),
				.b3(W3A10F),
				.b4(W3A11F),
				.b5(W3A12F),
				.b6(W3A20F),
				.b7(W3A21F),
				.b8(W3A22F),
				.c(c3F22A)
);

assign C322A=c3022A+c3122A+c3222A+c3322A+c3422A+c3522A+c3622A+c3722A+c3822A+c3922A+c3A22A+c3B22A+c3C22A+c3D22A+c3E22A+c3F22A;
assign A322A=(C322A>=0)?1:0;

assign P422A=A322A;

ninexnine_unit ninexnine_unit_4784(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3000B)
);

ninexnine_unit ninexnine_unit_4785(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3100B)
);

ninexnine_unit ninexnine_unit_4786(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3200B)
);

ninexnine_unit ninexnine_unit_4787(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3300B)
);

ninexnine_unit ninexnine_unit_4788(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3400B)
);

ninexnine_unit ninexnine_unit_4789(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3500B)
);

ninexnine_unit ninexnine_unit_4790(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3600B)
);

ninexnine_unit ninexnine_unit_4791(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3700B)
);

ninexnine_unit ninexnine_unit_4792(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3800B)
);

ninexnine_unit ninexnine_unit_4793(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3900B)
);

ninexnine_unit ninexnine_unit_4794(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A00B)
);

ninexnine_unit ninexnine_unit_4795(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B00B)
);

ninexnine_unit ninexnine_unit_4796(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C00B)
);

ninexnine_unit ninexnine_unit_4797(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D00B)
);

ninexnine_unit ninexnine_unit_4798(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E00B)
);

ninexnine_unit ninexnine_unit_4799(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F00B)
);

assign C300B=c3000B+c3100B+c3200B+c3300B+c3400B+c3500B+c3600B+c3700B+c3800B+c3900B+c3A00B+c3B00B+c3C00B+c3D00B+c3E00B+c3F00B;
assign A300B=(C300B>=0)?1:0;

assign P400B=A300B;

ninexnine_unit ninexnine_unit_4800(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3001B)
);

ninexnine_unit ninexnine_unit_4801(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3101B)
);

ninexnine_unit ninexnine_unit_4802(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3201B)
);

ninexnine_unit ninexnine_unit_4803(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3301B)
);

ninexnine_unit ninexnine_unit_4804(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3401B)
);

ninexnine_unit ninexnine_unit_4805(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3501B)
);

ninexnine_unit ninexnine_unit_4806(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3601B)
);

ninexnine_unit ninexnine_unit_4807(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3701B)
);

ninexnine_unit ninexnine_unit_4808(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3801B)
);

ninexnine_unit ninexnine_unit_4809(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3901B)
);

ninexnine_unit ninexnine_unit_4810(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A01B)
);

ninexnine_unit ninexnine_unit_4811(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B01B)
);

ninexnine_unit ninexnine_unit_4812(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C01B)
);

ninexnine_unit ninexnine_unit_4813(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D01B)
);

ninexnine_unit ninexnine_unit_4814(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E01B)
);

ninexnine_unit ninexnine_unit_4815(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F01B)
);

assign C301B=c3001B+c3101B+c3201B+c3301B+c3401B+c3501B+c3601B+c3701B+c3801B+c3901B+c3A01B+c3B01B+c3C01B+c3D01B+c3E01B+c3F01B;
assign A301B=(C301B>=0)?1:0;

assign P401B=A301B;

ninexnine_unit ninexnine_unit_4816(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3002B)
);

ninexnine_unit ninexnine_unit_4817(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3102B)
);

ninexnine_unit ninexnine_unit_4818(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3202B)
);

ninexnine_unit ninexnine_unit_4819(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3302B)
);

ninexnine_unit ninexnine_unit_4820(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3402B)
);

ninexnine_unit ninexnine_unit_4821(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3502B)
);

ninexnine_unit ninexnine_unit_4822(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3602B)
);

ninexnine_unit ninexnine_unit_4823(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3702B)
);

ninexnine_unit ninexnine_unit_4824(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3802B)
);

ninexnine_unit ninexnine_unit_4825(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3902B)
);

ninexnine_unit ninexnine_unit_4826(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A02B)
);

ninexnine_unit ninexnine_unit_4827(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B02B)
);

ninexnine_unit ninexnine_unit_4828(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C02B)
);

ninexnine_unit ninexnine_unit_4829(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D02B)
);

ninexnine_unit ninexnine_unit_4830(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E02B)
);

ninexnine_unit ninexnine_unit_4831(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F02B)
);

assign C302B=c3002B+c3102B+c3202B+c3302B+c3402B+c3502B+c3602B+c3702B+c3802B+c3902B+c3A02B+c3B02B+c3C02B+c3D02B+c3E02B+c3F02B;
assign A302B=(C302B>=0)?1:0;

assign P402B=A302B;

ninexnine_unit ninexnine_unit_4832(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3010B)
);

ninexnine_unit ninexnine_unit_4833(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3110B)
);

ninexnine_unit ninexnine_unit_4834(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3210B)
);

ninexnine_unit ninexnine_unit_4835(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3310B)
);

ninexnine_unit ninexnine_unit_4836(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3410B)
);

ninexnine_unit ninexnine_unit_4837(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3510B)
);

ninexnine_unit ninexnine_unit_4838(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3610B)
);

ninexnine_unit ninexnine_unit_4839(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3710B)
);

ninexnine_unit ninexnine_unit_4840(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3810B)
);

ninexnine_unit ninexnine_unit_4841(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3910B)
);

ninexnine_unit ninexnine_unit_4842(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A10B)
);

ninexnine_unit ninexnine_unit_4843(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B10B)
);

ninexnine_unit ninexnine_unit_4844(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C10B)
);

ninexnine_unit ninexnine_unit_4845(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D10B)
);

ninexnine_unit ninexnine_unit_4846(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E10B)
);

ninexnine_unit ninexnine_unit_4847(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F10B)
);

assign C310B=c3010B+c3110B+c3210B+c3310B+c3410B+c3510B+c3610B+c3710B+c3810B+c3910B+c3A10B+c3B10B+c3C10B+c3D10B+c3E10B+c3F10B;
assign A310B=(C310B>=0)?1:0;

assign P410B=A310B;

ninexnine_unit ninexnine_unit_4848(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3011B)
);

ninexnine_unit ninexnine_unit_4849(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3111B)
);

ninexnine_unit ninexnine_unit_4850(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3211B)
);

ninexnine_unit ninexnine_unit_4851(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3311B)
);

ninexnine_unit ninexnine_unit_4852(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3411B)
);

ninexnine_unit ninexnine_unit_4853(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3511B)
);

ninexnine_unit ninexnine_unit_4854(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3611B)
);

ninexnine_unit ninexnine_unit_4855(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3711B)
);

ninexnine_unit ninexnine_unit_4856(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3811B)
);

ninexnine_unit ninexnine_unit_4857(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3911B)
);

ninexnine_unit ninexnine_unit_4858(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A11B)
);

ninexnine_unit ninexnine_unit_4859(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B11B)
);

ninexnine_unit ninexnine_unit_4860(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C11B)
);

ninexnine_unit ninexnine_unit_4861(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D11B)
);

ninexnine_unit ninexnine_unit_4862(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E11B)
);

ninexnine_unit ninexnine_unit_4863(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F11B)
);

assign C311B=c3011B+c3111B+c3211B+c3311B+c3411B+c3511B+c3611B+c3711B+c3811B+c3911B+c3A11B+c3B11B+c3C11B+c3D11B+c3E11B+c3F11B;
assign A311B=(C311B>=0)?1:0;

assign P411B=A311B;

ninexnine_unit ninexnine_unit_4864(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3012B)
);

ninexnine_unit ninexnine_unit_4865(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3112B)
);

ninexnine_unit ninexnine_unit_4866(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3212B)
);

ninexnine_unit ninexnine_unit_4867(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3312B)
);

ninexnine_unit ninexnine_unit_4868(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3412B)
);

ninexnine_unit ninexnine_unit_4869(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3512B)
);

ninexnine_unit ninexnine_unit_4870(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3612B)
);

ninexnine_unit ninexnine_unit_4871(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3712B)
);

ninexnine_unit ninexnine_unit_4872(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3812B)
);

ninexnine_unit ninexnine_unit_4873(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3912B)
);

ninexnine_unit ninexnine_unit_4874(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A12B)
);

ninexnine_unit ninexnine_unit_4875(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B12B)
);

ninexnine_unit ninexnine_unit_4876(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C12B)
);

ninexnine_unit ninexnine_unit_4877(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D12B)
);

ninexnine_unit ninexnine_unit_4878(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E12B)
);

ninexnine_unit ninexnine_unit_4879(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F12B)
);

assign C312B=c3012B+c3112B+c3212B+c3312B+c3412B+c3512B+c3612B+c3712B+c3812B+c3912B+c3A12B+c3B12B+c3C12B+c3D12B+c3E12B+c3F12B;
assign A312B=(C312B>=0)?1:0;

assign P412B=A312B;

ninexnine_unit ninexnine_unit_4880(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3020B)
);

ninexnine_unit ninexnine_unit_4881(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3120B)
);

ninexnine_unit ninexnine_unit_4882(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3220B)
);

ninexnine_unit ninexnine_unit_4883(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3320B)
);

ninexnine_unit ninexnine_unit_4884(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3420B)
);

ninexnine_unit ninexnine_unit_4885(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3520B)
);

ninexnine_unit ninexnine_unit_4886(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3620B)
);

ninexnine_unit ninexnine_unit_4887(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3720B)
);

ninexnine_unit ninexnine_unit_4888(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3820B)
);

ninexnine_unit ninexnine_unit_4889(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3920B)
);

ninexnine_unit ninexnine_unit_4890(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A20B)
);

ninexnine_unit ninexnine_unit_4891(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B20B)
);

ninexnine_unit ninexnine_unit_4892(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C20B)
);

ninexnine_unit ninexnine_unit_4893(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D20B)
);

ninexnine_unit ninexnine_unit_4894(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E20B)
);

ninexnine_unit ninexnine_unit_4895(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F20B)
);

assign C320B=c3020B+c3120B+c3220B+c3320B+c3420B+c3520B+c3620B+c3720B+c3820B+c3920B+c3A20B+c3B20B+c3C20B+c3D20B+c3E20B+c3F20B;
assign A320B=(C320B>=0)?1:0;

assign P420B=A320B;

ninexnine_unit ninexnine_unit_4896(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3021B)
);

ninexnine_unit ninexnine_unit_4897(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3121B)
);

ninexnine_unit ninexnine_unit_4898(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3221B)
);

ninexnine_unit ninexnine_unit_4899(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3321B)
);

ninexnine_unit ninexnine_unit_4900(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3421B)
);

ninexnine_unit ninexnine_unit_4901(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3521B)
);

ninexnine_unit ninexnine_unit_4902(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3621B)
);

ninexnine_unit ninexnine_unit_4903(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3721B)
);

ninexnine_unit ninexnine_unit_4904(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3821B)
);

ninexnine_unit ninexnine_unit_4905(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3921B)
);

ninexnine_unit ninexnine_unit_4906(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A21B)
);

ninexnine_unit ninexnine_unit_4907(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B21B)
);

ninexnine_unit ninexnine_unit_4908(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C21B)
);

ninexnine_unit ninexnine_unit_4909(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D21B)
);

ninexnine_unit ninexnine_unit_4910(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E21B)
);

ninexnine_unit ninexnine_unit_4911(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F21B)
);

assign C321B=c3021B+c3121B+c3221B+c3321B+c3421B+c3521B+c3621B+c3721B+c3821B+c3921B+c3A21B+c3B21B+c3C21B+c3D21B+c3E21B+c3F21B;
assign A321B=(C321B>=0)?1:0;

assign P421B=A321B;

ninexnine_unit ninexnine_unit_4912(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3B000),
				.b1(W3B010),
				.b2(W3B020),
				.b3(W3B100),
				.b4(W3B110),
				.b5(W3B120),
				.b6(W3B200),
				.b7(W3B210),
				.b8(W3B220),
				.c(c3022B)
);

ninexnine_unit ninexnine_unit_4913(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3B001),
				.b1(W3B011),
				.b2(W3B021),
				.b3(W3B101),
				.b4(W3B111),
				.b5(W3B121),
				.b6(W3B201),
				.b7(W3B211),
				.b8(W3B221),
				.c(c3122B)
);

ninexnine_unit ninexnine_unit_4914(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3B002),
				.b1(W3B012),
				.b2(W3B022),
				.b3(W3B102),
				.b4(W3B112),
				.b5(W3B122),
				.b6(W3B202),
				.b7(W3B212),
				.b8(W3B222),
				.c(c3222B)
);

ninexnine_unit ninexnine_unit_4915(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3B003),
				.b1(W3B013),
				.b2(W3B023),
				.b3(W3B103),
				.b4(W3B113),
				.b5(W3B123),
				.b6(W3B203),
				.b7(W3B213),
				.b8(W3B223),
				.c(c3322B)
);

ninexnine_unit ninexnine_unit_4916(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3B004),
				.b1(W3B014),
				.b2(W3B024),
				.b3(W3B104),
				.b4(W3B114),
				.b5(W3B124),
				.b6(W3B204),
				.b7(W3B214),
				.b8(W3B224),
				.c(c3422B)
);

ninexnine_unit ninexnine_unit_4917(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3B005),
				.b1(W3B015),
				.b2(W3B025),
				.b3(W3B105),
				.b4(W3B115),
				.b5(W3B125),
				.b6(W3B205),
				.b7(W3B215),
				.b8(W3B225),
				.c(c3522B)
);

ninexnine_unit ninexnine_unit_4918(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3B006),
				.b1(W3B016),
				.b2(W3B026),
				.b3(W3B106),
				.b4(W3B116),
				.b5(W3B126),
				.b6(W3B206),
				.b7(W3B216),
				.b8(W3B226),
				.c(c3622B)
);

ninexnine_unit ninexnine_unit_4919(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3B007),
				.b1(W3B017),
				.b2(W3B027),
				.b3(W3B107),
				.b4(W3B117),
				.b5(W3B127),
				.b6(W3B207),
				.b7(W3B217),
				.b8(W3B227),
				.c(c3722B)
);

ninexnine_unit ninexnine_unit_4920(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3B008),
				.b1(W3B018),
				.b2(W3B028),
				.b3(W3B108),
				.b4(W3B118),
				.b5(W3B128),
				.b6(W3B208),
				.b7(W3B218),
				.b8(W3B228),
				.c(c3822B)
);

ninexnine_unit ninexnine_unit_4921(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3B009),
				.b1(W3B019),
				.b2(W3B029),
				.b3(W3B109),
				.b4(W3B119),
				.b5(W3B129),
				.b6(W3B209),
				.b7(W3B219),
				.b8(W3B229),
				.c(c3922B)
);

ninexnine_unit ninexnine_unit_4922(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3B00A),
				.b1(W3B01A),
				.b2(W3B02A),
				.b3(W3B10A),
				.b4(W3B11A),
				.b5(W3B12A),
				.b6(W3B20A),
				.b7(W3B21A),
				.b8(W3B22A),
				.c(c3A22B)
);

ninexnine_unit ninexnine_unit_4923(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3B00B),
				.b1(W3B01B),
				.b2(W3B02B),
				.b3(W3B10B),
				.b4(W3B11B),
				.b5(W3B12B),
				.b6(W3B20B),
				.b7(W3B21B),
				.b8(W3B22B),
				.c(c3B22B)
);

ninexnine_unit ninexnine_unit_4924(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3B00C),
				.b1(W3B01C),
				.b2(W3B02C),
				.b3(W3B10C),
				.b4(W3B11C),
				.b5(W3B12C),
				.b6(W3B20C),
				.b7(W3B21C),
				.b8(W3B22C),
				.c(c3C22B)
);

ninexnine_unit ninexnine_unit_4925(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3B00D),
				.b1(W3B01D),
				.b2(W3B02D),
				.b3(W3B10D),
				.b4(W3B11D),
				.b5(W3B12D),
				.b6(W3B20D),
				.b7(W3B21D),
				.b8(W3B22D),
				.c(c3D22B)
);

ninexnine_unit ninexnine_unit_4926(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3B00E),
				.b1(W3B01E),
				.b2(W3B02E),
				.b3(W3B10E),
				.b4(W3B11E),
				.b5(W3B12E),
				.b6(W3B20E),
				.b7(W3B21E),
				.b8(W3B22E),
				.c(c3E22B)
);

ninexnine_unit ninexnine_unit_4927(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3B00F),
				.b1(W3B01F),
				.b2(W3B02F),
				.b3(W3B10F),
				.b4(W3B11F),
				.b5(W3B12F),
				.b6(W3B20F),
				.b7(W3B21F),
				.b8(W3B22F),
				.c(c3F22B)
);

assign C322B=c3022B+c3122B+c3222B+c3322B+c3422B+c3522B+c3622B+c3722B+c3822B+c3922B+c3A22B+c3B22B+c3C22B+c3D22B+c3E22B+c3F22B;
assign A322B=(C322B>=0)?1:0;

assign P422B=A322B;

ninexnine_unit ninexnine_unit_4928(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3000C)
);

ninexnine_unit ninexnine_unit_4929(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3100C)
);

ninexnine_unit ninexnine_unit_4930(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3200C)
);

ninexnine_unit ninexnine_unit_4931(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3300C)
);

ninexnine_unit ninexnine_unit_4932(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3400C)
);

ninexnine_unit ninexnine_unit_4933(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3500C)
);

ninexnine_unit ninexnine_unit_4934(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3600C)
);

ninexnine_unit ninexnine_unit_4935(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3700C)
);

ninexnine_unit ninexnine_unit_4936(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3800C)
);

ninexnine_unit ninexnine_unit_4937(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3900C)
);

ninexnine_unit ninexnine_unit_4938(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A00C)
);

ninexnine_unit ninexnine_unit_4939(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B00C)
);

ninexnine_unit ninexnine_unit_4940(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C00C)
);

ninexnine_unit ninexnine_unit_4941(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D00C)
);

ninexnine_unit ninexnine_unit_4942(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E00C)
);

ninexnine_unit ninexnine_unit_4943(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F00C)
);

assign C300C=c3000C+c3100C+c3200C+c3300C+c3400C+c3500C+c3600C+c3700C+c3800C+c3900C+c3A00C+c3B00C+c3C00C+c3D00C+c3E00C+c3F00C;
assign A300C=(C300C>=0)?1:0;

assign P400C=A300C;

ninexnine_unit ninexnine_unit_4944(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3001C)
);

ninexnine_unit ninexnine_unit_4945(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3101C)
);

ninexnine_unit ninexnine_unit_4946(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3201C)
);

ninexnine_unit ninexnine_unit_4947(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3301C)
);

ninexnine_unit ninexnine_unit_4948(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3401C)
);

ninexnine_unit ninexnine_unit_4949(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3501C)
);

ninexnine_unit ninexnine_unit_4950(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3601C)
);

ninexnine_unit ninexnine_unit_4951(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3701C)
);

ninexnine_unit ninexnine_unit_4952(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3801C)
);

ninexnine_unit ninexnine_unit_4953(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3901C)
);

ninexnine_unit ninexnine_unit_4954(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A01C)
);

ninexnine_unit ninexnine_unit_4955(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B01C)
);

ninexnine_unit ninexnine_unit_4956(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C01C)
);

ninexnine_unit ninexnine_unit_4957(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D01C)
);

ninexnine_unit ninexnine_unit_4958(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E01C)
);

ninexnine_unit ninexnine_unit_4959(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F01C)
);

assign C301C=c3001C+c3101C+c3201C+c3301C+c3401C+c3501C+c3601C+c3701C+c3801C+c3901C+c3A01C+c3B01C+c3C01C+c3D01C+c3E01C+c3F01C;
assign A301C=(C301C>=0)?1:0;

assign P401C=A301C;

ninexnine_unit ninexnine_unit_4960(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3002C)
);

ninexnine_unit ninexnine_unit_4961(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3102C)
);

ninexnine_unit ninexnine_unit_4962(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3202C)
);

ninexnine_unit ninexnine_unit_4963(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3302C)
);

ninexnine_unit ninexnine_unit_4964(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3402C)
);

ninexnine_unit ninexnine_unit_4965(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3502C)
);

ninexnine_unit ninexnine_unit_4966(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3602C)
);

ninexnine_unit ninexnine_unit_4967(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3702C)
);

ninexnine_unit ninexnine_unit_4968(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3802C)
);

ninexnine_unit ninexnine_unit_4969(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3902C)
);

ninexnine_unit ninexnine_unit_4970(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A02C)
);

ninexnine_unit ninexnine_unit_4971(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B02C)
);

ninexnine_unit ninexnine_unit_4972(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C02C)
);

ninexnine_unit ninexnine_unit_4973(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D02C)
);

ninexnine_unit ninexnine_unit_4974(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E02C)
);

ninexnine_unit ninexnine_unit_4975(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F02C)
);

assign C302C=c3002C+c3102C+c3202C+c3302C+c3402C+c3502C+c3602C+c3702C+c3802C+c3902C+c3A02C+c3B02C+c3C02C+c3D02C+c3E02C+c3F02C;
assign A302C=(C302C>=0)?1:0;

assign P402C=A302C;

ninexnine_unit ninexnine_unit_4976(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3010C)
);

ninexnine_unit ninexnine_unit_4977(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3110C)
);

ninexnine_unit ninexnine_unit_4978(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3210C)
);

ninexnine_unit ninexnine_unit_4979(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3310C)
);

ninexnine_unit ninexnine_unit_4980(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3410C)
);

ninexnine_unit ninexnine_unit_4981(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3510C)
);

ninexnine_unit ninexnine_unit_4982(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3610C)
);

ninexnine_unit ninexnine_unit_4983(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3710C)
);

ninexnine_unit ninexnine_unit_4984(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3810C)
);

ninexnine_unit ninexnine_unit_4985(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3910C)
);

ninexnine_unit ninexnine_unit_4986(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A10C)
);

ninexnine_unit ninexnine_unit_4987(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B10C)
);

ninexnine_unit ninexnine_unit_4988(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C10C)
);

ninexnine_unit ninexnine_unit_4989(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D10C)
);

ninexnine_unit ninexnine_unit_4990(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E10C)
);

ninexnine_unit ninexnine_unit_4991(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F10C)
);

assign C310C=c3010C+c3110C+c3210C+c3310C+c3410C+c3510C+c3610C+c3710C+c3810C+c3910C+c3A10C+c3B10C+c3C10C+c3D10C+c3E10C+c3F10C;
assign A310C=(C310C>=0)?1:0;

assign P410C=A310C;

ninexnine_unit ninexnine_unit_4992(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3011C)
);

ninexnine_unit ninexnine_unit_4993(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3111C)
);

ninexnine_unit ninexnine_unit_4994(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3211C)
);

ninexnine_unit ninexnine_unit_4995(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3311C)
);

ninexnine_unit ninexnine_unit_4996(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3411C)
);

ninexnine_unit ninexnine_unit_4997(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3511C)
);

ninexnine_unit ninexnine_unit_4998(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3611C)
);

ninexnine_unit ninexnine_unit_4999(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3711C)
);

ninexnine_unit ninexnine_unit_5000(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3811C)
);

ninexnine_unit ninexnine_unit_5001(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3911C)
);

ninexnine_unit ninexnine_unit_5002(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A11C)
);

ninexnine_unit ninexnine_unit_5003(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B11C)
);

ninexnine_unit ninexnine_unit_5004(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C11C)
);

ninexnine_unit ninexnine_unit_5005(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D11C)
);

ninexnine_unit ninexnine_unit_5006(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E11C)
);

ninexnine_unit ninexnine_unit_5007(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F11C)
);

assign C311C=c3011C+c3111C+c3211C+c3311C+c3411C+c3511C+c3611C+c3711C+c3811C+c3911C+c3A11C+c3B11C+c3C11C+c3D11C+c3E11C+c3F11C;
assign A311C=(C311C>=0)?1:0;

assign P411C=A311C;

ninexnine_unit ninexnine_unit_5008(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3012C)
);

ninexnine_unit ninexnine_unit_5009(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3112C)
);

ninexnine_unit ninexnine_unit_5010(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3212C)
);

ninexnine_unit ninexnine_unit_5011(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3312C)
);

ninexnine_unit ninexnine_unit_5012(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3412C)
);

ninexnine_unit ninexnine_unit_5013(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3512C)
);

ninexnine_unit ninexnine_unit_5014(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3612C)
);

ninexnine_unit ninexnine_unit_5015(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3712C)
);

ninexnine_unit ninexnine_unit_5016(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3812C)
);

ninexnine_unit ninexnine_unit_5017(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3912C)
);

ninexnine_unit ninexnine_unit_5018(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A12C)
);

ninexnine_unit ninexnine_unit_5019(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B12C)
);

ninexnine_unit ninexnine_unit_5020(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C12C)
);

ninexnine_unit ninexnine_unit_5021(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D12C)
);

ninexnine_unit ninexnine_unit_5022(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E12C)
);

ninexnine_unit ninexnine_unit_5023(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F12C)
);

assign C312C=c3012C+c3112C+c3212C+c3312C+c3412C+c3512C+c3612C+c3712C+c3812C+c3912C+c3A12C+c3B12C+c3C12C+c3D12C+c3E12C+c3F12C;
assign A312C=(C312C>=0)?1:0;

assign P412C=A312C;

ninexnine_unit ninexnine_unit_5024(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3020C)
);

ninexnine_unit ninexnine_unit_5025(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3120C)
);

ninexnine_unit ninexnine_unit_5026(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3220C)
);

ninexnine_unit ninexnine_unit_5027(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3320C)
);

ninexnine_unit ninexnine_unit_5028(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3420C)
);

ninexnine_unit ninexnine_unit_5029(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3520C)
);

ninexnine_unit ninexnine_unit_5030(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3620C)
);

ninexnine_unit ninexnine_unit_5031(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3720C)
);

ninexnine_unit ninexnine_unit_5032(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3820C)
);

ninexnine_unit ninexnine_unit_5033(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3920C)
);

ninexnine_unit ninexnine_unit_5034(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A20C)
);

ninexnine_unit ninexnine_unit_5035(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B20C)
);

ninexnine_unit ninexnine_unit_5036(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C20C)
);

ninexnine_unit ninexnine_unit_5037(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D20C)
);

ninexnine_unit ninexnine_unit_5038(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E20C)
);

ninexnine_unit ninexnine_unit_5039(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F20C)
);

assign C320C=c3020C+c3120C+c3220C+c3320C+c3420C+c3520C+c3620C+c3720C+c3820C+c3920C+c3A20C+c3B20C+c3C20C+c3D20C+c3E20C+c3F20C;
assign A320C=(C320C>=0)?1:0;

assign P420C=A320C;

ninexnine_unit ninexnine_unit_5040(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3021C)
);

ninexnine_unit ninexnine_unit_5041(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3121C)
);

ninexnine_unit ninexnine_unit_5042(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3221C)
);

ninexnine_unit ninexnine_unit_5043(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3321C)
);

ninexnine_unit ninexnine_unit_5044(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3421C)
);

ninexnine_unit ninexnine_unit_5045(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3521C)
);

ninexnine_unit ninexnine_unit_5046(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3621C)
);

ninexnine_unit ninexnine_unit_5047(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3721C)
);

ninexnine_unit ninexnine_unit_5048(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3821C)
);

ninexnine_unit ninexnine_unit_5049(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3921C)
);

ninexnine_unit ninexnine_unit_5050(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A21C)
);

ninexnine_unit ninexnine_unit_5051(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B21C)
);

ninexnine_unit ninexnine_unit_5052(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C21C)
);

ninexnine_unit ninexnine_unit_5053(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D21C)
);

ninexnine_unit ninexnine_unit_5054(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E21C)
);

ninexnine_unit ninexnine_unit_5055(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F21C)
);

assign C321C=c3021C+c3121C+c3221C+c3321C+c3421C+c3521C+c3621C+c3721C+c3821C+c3921C+c3A21C+c3B21C+c3C21C+c3D21C+c3E21C+c3F21C;
assign A321C=(C321C>=0)?1:0;

assign P421C=A321C;

ninexnine_unit ninexnine_unit_5056(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3C000),
				.b1(W3C010),
				.b2(W3C020),
				.b3(W3C100),
				.b4(W3C110),
				.b5(W3C120),
				.b6(W3C200),
				.b7(W3C210),
				.b8(W3C220),
				.c(c3022C)
);

ninexnine_unit ninexnine_unit_5057(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3C001),
				.b1(W3C011),
				.b2(W3C021),
				.b3(W3C101),
				.b4(W3C111),
				.b5(W3C121),
				.b6(W3C201),
				.b7(W3C211),
				.b8(W3C221),
				.c(c3122C)
);

ninexnine_unit ninexnine_unit_5058(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3C002),
				.b1(W3C012),
				.b2(W3C022),
				.b3(W3C102),
				.b4(W3C112),
				.b5(W3C122),
				.b6(W3C202),
				.b7(W3C212),
				.b8(W3C222),
				.c(c3222C)
);

ninexnine_unit ninexnine_unit_5059(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3C003),
				.b1(W3C013),
				.b2(W3C023),
				.b3(W3C103),
				.b4(W3C113),
				.b5(W3C123),
				.b6(W3C203),
				.b7(W3C213),
				.b8(W3C223),
				.c(c3322C)
);

ninexnine_unit ninexnine_unit_5060(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3C004),
				.b1(W3C014),
				.b2(W3C024),
				.b3(W3C104),
				.b4(W3C114),
				.b5(W3C124),
				.b6(W3C204),
				.b7(W3C214),
				.b8(W3C224),
				.c(c3422C)
);

ninexnine_unit ninexnine_unit_5061(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3C005),
				.b1(W3C015),
				.b2(W3C025),
				.b3(W3C105),
				.b4(W3C115),
				.b5(W3C125),
				.b6(W3C205),
				.b7(W3C215),
				.b8(W3C225),
				.c(c3522C)
);

ninexnine_unit ninexnine_unit_5062(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3C006),
				.b1(W3C016),
				.b2(W3C026),
				.b3(W3C106),
				.b4(W3C116),
				.b5(W3C126),
				.b6(W3C206),
				.b7(W3C216),
				.b8(W3C226),
				.c(c3622C)
);

ninexnine_unit ninexnine_unit_5063(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3C007),
				.b1(W3C017),
				.b2(W3C027),
				.b3(W3C107),
				.b4(W3C117),
				.b5(W3C127),
				.b6(W3C207),
				.b7(W3C217),
				.b8(W3C227),
				.c(c3722C)
);

ninexnine_unit ninexnine_unit_5064(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3C008),
				.b1(W3C018),
				.b2(W3C028),
				.b3(W3C108),
				.b4(W3C118),
				.b5(W3C128),
				.b6(W3C208),
				.b7(W3C218),
				.b8(W3C228),
				.c(c3822C)
);

ninexnine_unit ninexnine_unit_5065(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3C009),
				.b1(W3C019),
				.b2(W3C029),
				.b3(W3C109),
				.b4(W3C119),
				.b5(W3C129),
				.b6(W3C209),
				.b7(W3C219),
				.b8(W3C229),
				.c(c3922C)
);

ninexnine_unit ninexnine_unit_5066(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3C00A),
				.b1(W3C01A),
				.b2(W3C02A),
				.b3(W3C10A),
				.b4(W3C11A),
				.b5(W3C12A),
				.b6(W3C20A),
				.b7(W3C21A),
				.b8(W3C22A),
				.c(c3A22C)
);

ninexnine_unit ninexnine_unit_5067(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3C00B),
				.b1(W3C01B),
				.b2(W3C02B),
				.b3(W3C10B),
				.b4(W3C11B),
				.b5(W3C12B),
				.b6(W3C20B),
				.b7(W3C21B),
				.b8(W3C22B),
				.c(c3B22C)
);

ninexnine_unit ninexnine_unit_5068(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3C00C),
				.b1(W3C01C),
				.b2(W3C02C),
				.b3(W3C10C),
				.b4(W3C11C),
				.b5(W3C12C),
				.b6(W3C20C),
				.b7(W3C21C),
				.b8(W3C22C),
				.c(c3C22C)
);

ninexnine_unit ninexnine_unit_5069(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3C00D),
				.b1(W3C01D),
				.b2(W3C02D),
				.b3(W3C10D),
				.b4(W3C11D),
				.b5(W3C12D),
				.b6(W3C20D),
				.b7(W3C21D),
				.b8(W3C22D),
				.c(c3D22C)
);

ninexnine_unit ninexnine_unit_5070(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3C00E),
				.b1(W3C01E),
				.b2(W3C02E),
				.b3(W3C10E),
				.b4(W3C11E),
				.b5(W3C12E),
				.b6(W3C20E),
				.b7(W3C21E),
				.b8(W3C22E),
				.c(c3E22C)
);

ninexnine_unit ninexnine_unit_5071(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3C00F),
				.b1(W3C01F),
				.b2(W3C02F),
				.b3(W3C10F),
				.b4(W3C11F),
				.b5(W3C12F),
				.b6(W3C20F),
				.b7(W3C21F),
				.b8(W3C22F),
				.c(c3F22C)
);

assign C322C=c3022C+c3122C+c3222C+c3322C+c3422C+c3522C+c3622C+c3722C+c3822C+c3922C+c3A22C+c3B22C+c3C22C+c3D22C+c3E22C+c3F22C;
assign A322C=(C322C>=0)?1:0;

assign P422C=A322C;

ninexnine_unit ninexnine_unit_5072(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3000D)
);

ninexnine_unit ninexnine_unit_5073(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3100D)
);

ninexnine_unit ninexnine_unit_5074(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3200D)
);

ninexnine_unit ninexnine_unit_5075(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3300D)
);

ninexnine_unit ninexnine_unit_5076(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3400D)
);

ninexnine_unit ninexnine_unit_5077(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3500D)
);

ninexnine_unit ninexnine_unit_5078(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3600D)
);

ninexnine_unit ninexnine_unit_5079(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3700D)
);

ninexnine_unit ninexnine_unit_5080(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3800D)
);

ninexnine_unit ninexnine_unit_5081(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3900D)
);

ninexnine_unit ninexnine_unit_5082(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A00D)
);

ninexnine_unit ninexnine_unit_5083(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B00D)
);

ninexnine_unit ninexnine_unit_5084(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C00D)
);

ninexnine_unit ninexnine_unit_5085(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D00D)
);

ninexnine_unit ninexnine_unit_5086(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E00D)
);

ninexnine_unit ninexnine_unit_5087(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F00D)
);

assign C300D=c3000D+c3100D+c3200D+c3300D+c3400D+c3500D+c3600D+c3700D+c3800D+c3900D+c3A00D+c3B00D+c3C00D+c3D00D+c3E00D+c3F00D;
assign A300D=(C300D>=0)?1:0;

assign P400D=A300D;

ninexnine_unit ninexnine_unit_5088(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3001D)
);

ninexnine_unit ninexnine_unit_5089(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3101D)
);

ninexnine_unit ninexnine_unit_5090(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3201D)
);

ninexnine_unit ninexnine_unit_5091(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3301D)
);

ninexnine_unit ninexnine_unit_5092(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3401D)
);

ninexnine_unit ninexnine_unit_5093(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3501D)
);

ninexnine_unit ninexnine_unit_5094(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3601D)
);

ninexnine_unit ninexnine_unit_5095(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3701D)
);

ninexnine_unit ninexnine_unit_5096(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3801D)
);

ninexnine_unit ninexnine_unit_5097(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3901D)
);

ninexnine_unit ninexnine_unit_5098(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A01D)
);

ninexnine_unit ninexnine_unit_5099(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B01D)
);

ninexnine_unit ninexnine_unit_5100(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C01D)
);

ninexnine_unit ninexnine_unit_5101(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D01D)
);

ninexnine_unit ninexnine_unit_5102(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E01D)
);

ninexnine_unit ninexnine_unit_5103(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F01D)
);

assign C301D=c3001D+c3101D+c3201D+c3301D+c3401D+c3501D+c3601D+c3701D+c3801D+c3901D+c3A01D+c3B01D+c3C01D+c3D01D+c3E01D+c3F01D;
assign A301D=(C301D>=0)?1:0;

assign P401D=A301D;

ninexnine_unit ninexnine_unit_5104(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3002D)
);

ninexnine_unit ninexnine_unit_5105(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3102D)
);

ninexnine_unit ninexnine_unit_5106(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3202D)
);

ninexnine_unit ninexnine_unit_5107(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3302D)
);

ninexnine_unit ninexnine_unit_5108(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3402D)
);

ninexnine_unit ninexnine_unit_5109(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3502D)
);

ninexnine_unit ninexnine_unit_5110(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3602D)
);

ninexnine_unit ninexnine_unit_5111(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3702D)
);

ninexnine_unit ninexnine_unit_5112(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3802D)
);

ninexnine_unit ninexnine_unit_5113(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3902D)
);

ninexnine_unit ninexnine_unit_5114(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A02D)
);

ninexnine_unit ninexnine_unit_5115(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B02D)
);

ninexnine_unit ninexnine_unit_5116(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C02D)
);

ninexnine_unit ninexnine_unit_5117(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D02D)
);

ninexnine_unit ninexnine_unit_5118(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E02D)
);

ninexnine_unit ninexnine_unit_5119(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F02D)
);

assign C302D=c3002D+c3102D+c3202D+c3302D+c3402D+c3502D+c3602D+c3702D+c3802D+c3902D+c3A02D+c3B02D+c3C02D+c3D02D+c3E02D+c3F02D;
assign A302D=(C302D>=0)?1:0;

assign P402D=A302D;

ninexnine_unit ninexnine_unit_5120(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3010D)
);

ninexnine_unit ninexnine_unit_5121(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3110D)
);

ninexnine_unit ninexnine_unit_5122(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3210D)
);

ninexnine_unit ninexnine_unit_5123(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3310D)
);

ninexnine_unit ninexnine_unit_5124(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3410D)
);

ninexnine_unit ninexnine_unit_5125(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3510D)
);

ninexnine_unit ninexnine_unit_5126(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3610D)
);

ninexnine_unit ninexnine_unit_5127(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3710D)
);

ninexnine_unit ninexnine_unit_5128(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3810D)
);

ninexnine_unit ninexnine_unit_5129(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3910D)
);

ninexnine_unit ninexnine_unit_5130(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A10D)
);

ninexnine_unit ninexnine_unit_5131(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B10D)
);

ninexnine_unit ninexnine_unit_5132(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C10D)
);

ninexnine_unit ninexnine_unit_5133(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D10D)
);

ninexnine_unit ninexnine_unit_5134(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E10D)
);

ninexnine_unit ninexnine_unit_5135(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F10D)
);

assign C310D=c3010D+c3110D+c3210D+c3310D+c3410D+c3510D+c3610D+c3710D+c3810D+c3910D+c3A10D+c3B10D+c3C10D+c3D10D+c3E10D+c3F10D;
assign A310D=(C310D>=0)?1:0;

assign P410D=A310D;

ninexnine_unit ninexnine_unit_5136(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3011D)
);

ninexnine_unit ninexnine_unit_5137(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3111D)
);

ninexnine_unit ninexnine_unit_5138(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3211D)
);

ninexnine_unit ninexnine_unit_5139(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3311D)
);

ninexnine_unit ninexnine_unit_5140(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3411D)
);

ninexnine_unit ninexnine_unit_5141(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3511D)
);

ninexnine_unit ninexnine_unit_5142(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3611D)
);

ninexnine_unit ninexnine_unit_5143(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3711D)
);

ninexnine_unit ninexnine_unit_5144(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3811D)
);

ninexnine_unit ninexnine_unit_5145(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3911D)
);

ninexnine_unit ninexnine_unit_5146(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A11D)
);

ninexnine_unit ninexnine_unit_5147(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B11D)
);

ninexnine_unit ninexnine_unit_5148(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C11D)
);

ninexnine_unit ninexnine_unit_5149(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D11D)
);

ninexnine_unit ninexnine_unit_5150(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E11D)
);

ninexnine_unit ninexnine_unit_5151(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F11D)
);

assign C311D=c3011D+c3111D+c3211D+c3311D+c3411D+c3511D+c3611D+c3711D+c3811D+c3911D+c3A11D+c3B11D+c3C11D+c3D11D+c3E11D+c3F11D;
assign A311D=(C311D>=0)?1:0;

assign P411D=A311D;

ninexnine_unit ninexnine_unit_5152(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3012D)
);

ninexnine_unit ninexnine_unit_5153(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3112D)
);

ninexnine_unit ninexnine_unit_5154(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3212D)
);

ninexnine_unit ninexnine_unit_5155(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3312D)
);

ninexnine_unit ninexnine_unit_5156(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3412D)
);

ninexnine_unit ninexnine_unit_5157(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3512D)
);

ninexnine_unit ninexnine_unit_5158(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3612D)
);

ninexnine_unit ninexnine_unit_5159(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3712D)
);

ninexnine_unit ninexnine_unit_5160(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3812D)
);

ninexnine_unit ninexnine_unit_5161(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3912D)
);

ninexnine_unit ninexnine_unit_5162(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A12D)
);

ninexnine_unit ninexnine_unit_5163(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B12D)
);

ninexnine_unit ninexnine_unit_5164(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C12D)
);

ninexnine_unit ninexnine_unit_5165(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D12D)
);

ninexnine_unit ninexnine_unit_5166(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E12D)
);

ninexnine_unit ninexnine_unit_5167(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F12D)
);

assign C312D=c3012D+c3112D+c3212D+c3312D+c3412D+c3512D+c3612D+c3712D+c3812D+c3912D+c3A12D+c3B12D+c3C12D+c3D12D+c3E12D+c3F12D;
assign A312D=(C312D>=0)?1:0;

assign P412D=A312D;

ninexnine_unit ninexnine_unit_5168(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3020D)
);

ninexnine_unit ninexnine_unit_5169(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3120D)
);

ninexnine_unit ninexnine_unit_5170(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3220D)
);

ninexnine_unit ninexnine_unit_5171(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3320D)
);

ninexnine_unit ninexnine_unit_5172(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3420D)
);

ninexnine_unit ninexnine_unit_5173(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3520D)
);

ninexnine_unit ninexnine_unit_5174(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3620D)
);

ninexnine_unit ninexnine_unit_5175(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3720D)
);

ninexnine_unit ninexnine_unit_5176(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3820D)
);

ninexnine_unit ninexnine_unit_5177(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3920D)
);

ninexnine_unit ninexnine_unit_5178(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A20D)
);

ninexnine_unit ninexnine_unit_5179(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B20D)
);

ninexnine_unit ninexnine_unit_5180(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C20D)
);

ninexnine_unit ninexnine_unit_5181(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D20D)
);

ninexnine_unit ninexnine_unit_5182(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E20D)
);

ninexnine_unit ninexnine_unit_5183(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F20D)
);

assign C320D=c3020D+c3120D+c3220D+c3320D+c3420D+c3520D+c3620D+c3720D+c3820D+c3920D+c3A20D+c3B20D+c3C20D+c3D20D+c3E20D+c3F20D;
assign A320D=(C320D>=0)?1:0;

assign P420D=A320D;

ninexnine_unit ninexnine_unit_5184(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3021D)
);

ninexnine_unit ninexnine_unit_5185(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3121D)
);

ninexnine_unit ninexnine_unit_5186(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3221D)
);

ninexnine_unit ninexnine_unit_5187(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3321D)
);

ninexnine_unit ninexnine_unit_5188(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3421D)
);

ninexnine_unit ninexnine_unit_5189(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3521D)
);

ninexnine_unit ninexnine_unit_5190(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3621D)
);

ninexnine_unit ninexnine_unit_5191(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3721D)
);

ninexnine_unit ninexnine_unit_5192(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3821D)
);

ninexnine_unit ninexnine_unit_5193(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3921D)
);

ninexnine_unit ninexnine_unit_5194(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A21D)
);

ninexnine_unit ninexnine_unit_5195(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B21D)
);

ninexnine_unit ninexnine_unit_5196(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C21D)
);

ninexnine_unit ninexnine_unit_5197(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D21D)
);

ninexnine_unit ninexnine_unit_5198(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E21D)
);

ninexnine_unit ninexnine_unit_5199(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F21D)
);

assign C321D=c3021D+c3121D+c3221D+c3321D+c3421D+c3521D+c3621D+c3721D+c3821D+c3921D+c3A21D+c3B21D+c3C21D+c3D21D+c3E21D+c3F21D;
assign A321D=(C321D>=0)?1:0;

assign P421D=A321D;

ninexnine_unit ninexnine_unit_5200(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3D000),
				.b1(W3D010),
				.b2(W3D020),
				.b3(W3D100),
				.b4(W3D110),
				.b5(W3D120),
				.b6(W3D200),
				.b7(W3D210),
				.b8(W3D220),
				.c(c3022D)
);

ninexnine_unit ninexnine_unit_5201(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3D001),
				.b1(W3D011),
				.b2(W3D021),
				.b3(W3D101),
				.b4(W3D111),
				.b5(W3D121),
				.b6(W3D201),
				.b7(W3D211),
				.b8(W3D221),
				.c(c3122D)
);

ninexnine_unit ninexnine_unit_5202(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3D002),
				.b1(W3D012),
				.b2(W3D022),
				.b3(W3D102),
				.b4(W3D112),
				.b5(W3D122),
				.b6(W3D202),
				.b7(W3D212),
				.b8(W3D222),
				.c(c3222D)
);

ninexnine_unit ninexnine_unit_5203(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3D003),
				.b1(W3D013),
				.b2(W3D023),
				.b3(W3D103),
				.b4(W3D113),
				.b5(W3D123),
				.b6(W3D203),
				.b7(W3D213),
				.b8(W3D223),
				.c(c3322D)
);

ninexnine_unit ninexnine_unit_5204(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3D004),
				.b1(W3D014),
				.b2(W3D024),
				.b3(W3D104),
				.b4(W3D114),
				.b5(W3D124),
				.b6(W3D204),
				.b7(W3D214),
				.b8(W3D224),
				.c(c3422D)
);

ninexnine_unit ninexnine_unit_5205(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3D005),
				.b1(W3D015),
				.b2(W3D025),
				.b3(W3D105),
				.b4(W3D115),
				.b5(W3D125),
				.b6(W3D205),
				.b7(W3D215),
				.b8(W3D225),
				.c(c3522D)
);

ninexnine_unit ninexnine_unit_5206(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3D006),
				.b1(W3D016),
				.b2(W3D026),
				.b3(W3D106),
				.b4(W3D116),
				.b5(W3D126),
				.b6(W3D206),
				.b7(W3D216),
				.b8(W3D226),
				.c(c3622D)
);

ninexnine_unit ninexnine_unit_5207(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3D007),
				.b1(W3D017),
				.b2(W3D027),
				.b3(W3D107),
				.b4(W3D117),
				.b5(W3D127),
				.b6(W3D207),
				.b7(W3D217),
				.b8(W3D227),
				.c(c3722D)
);

ninexnine_unit ninexnine_unit_5208(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3D008),
				.b1(W3D018),
				.b2(W3D028),
				.b3(W3D108),
				.b4(W3D118),
				.b5(W3D128),
				.b6(W3D208),
				.b7(W3D218),
				.b8(W3D228),
				.c(c3822D)
);

ninexnine_unit ninexnine_unit_5209(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3D009),
				.b1(W3D019),
				.b2(W3D029),
				.b3(W3D109),
				.b4(W3D119),
				.b5(W3D129),
				.b6(W3D209),
				.b7(W3D219),
				.b8(W3D229),
				.c(c3922D)
);

ninexnine_unit ninexnine_unit_5210(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3D00A),
				.b1(W3D01A),
				.b2(W3D02A),
				.b3(W3D10A),
				.b4(W3D11A),
				.b5(W3D12A),
				.b6(W3D20A),
				.b7(W3D21A),
				.b8(W3D22A),
				.c(c3A22D)
);

ninexnine_unit ninexnine_unit_5211(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3D00B),
				.b1(W3D01B),
				.b2(W3D02B),
				.b3(W3D10B),
				.b4(W3D11B),
				.b5(W3D12B),
				.b6(W3D20B),
				.b7(W3D21B),
				.b8(W3D22B),
				.c(c3B22D)
);

ninexnine_unit ninexnine_unit_5212(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3D00C),
				.b1(W3D01C),
				.b2(W3D02C),
				.b3(W3D10C),
				.b4(W3D11C),
				.b5(W3D12C),
				.b6(W3D20C),
				.b7(W3D21C),
				.b8(W3D22C),
				.c(c3C22D)
);

ninexnine_unit ninexnine_unit_5213(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3D00D),
				.b1(W3D01D),
				.b2(W3D02D),
				.b3(W3D10D),
				.b4(W3D11D),
				.b5(W3D12D),
				.b6(W3D20D),
				.b7(W3D21D),
				.b8(W3D22D),
				.c(c3D22D)
);

ninexnine_unit ninexnine_unit_5214(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3D00E),
				.b1(W3D01E),
				.b2(W3D02E),
				.b3(W3D10E),
				.b4(W3D11E),
				.b5(W3D12E),
				.b6(W3D20E),
				.b7(W3D21E),
				.b8(W3D22E),
				.c(c3E22D)
);

ninexnine_unit ninexnine_unit_5215(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3D00F),
				.b1(W3D01F),
				.b2(W3D02F),
				.b3(W3D10F),
				.b4(W3D11F),
				.b5(W3D12F),
				.b6(W3D20F),
				.b7(W3D21F),
				.b8(W3D22F),
				.c(c3F22D)
);

assign C322D=c3022D+c3122D+c3222D+c3322D+c3422D+c3522D+c3622D+c3722D+c3822D+c3922D+c3A22D+c3B22D+c3C22D+c3D22D+c3E22D+c3F22D;
assign A322D=(C322D>=0)?1:0;

assign P422D=A322D;

ninexnine_unit ninexnine_unit_5216(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3000E)
);

ninexnine_unit ninexnine_unit_5217(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3100E)
);

ninexnine_unit ninexnine_unit_5218(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3200E)
);

ninexnine_unit ninexnine_unit_5219(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3300E)
);

ninexnine_unit ninexnine_unit_5220(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3400E)
);

ninexnine_unit ninexnine_unit_5221(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3500E)
);

ninexnine_unit ninexnine_unit_5222(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3600E)
);

ninexnine_unit ninexnine_unit_5223(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3700E)
);

ninexnine_unit ninexnine_unit_5224(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3800E)
);

ninexnine_unit ninexnine_unit_5225(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3900E)
);

ninexnine_unit ninexnine_unit_5226(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A00E)
);

ninexnine_unit ninexnine_unit_5227(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B00E)
);

ninexnine_unit ninexnine_unit_5228(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C00E)
);

ninexnine_unit ninexnine_unit_5229(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D00E)
);

ninexnine_unit ninexnine_unit_5230(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E00E)
);

ninexnine_unit ninexnine_unit_5231(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F00E)
);

assign C300E=c3000E+c3100E+c3200E+c3300E+c3400E+c3500E+c3600E+c3700E+c3800E+c3900E+c3A00E+c3B00E+c3C00E+c3D00E+c3E00E+c3F00E;
assign A300E=(C300E>=0)?1:0;

assign P400E=A300E;

ninexnine_unit ninexnine_unit_5232(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3001E)
);

ninexnine_unit ninexnine_unit_5233(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3101E)
);

ninexnine_unit ninexnine_unit_5234(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3201E)
);

ninexnine_unit ninexnine_unit_5235(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3301E)
);

ninexnine_unit ninexnine_unit_5236(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3401E)
);

ninexnine_unit ninexnine_unit_5237(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3501E)
);

ninexnine_unit ninexnine_unit_5238(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3601E)
);

ninexnine_unit ninexnine_unit_5239(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3701E)
);

ninexnine_unit ninexnine_unit_5240(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3801E)
);

ninexnine_unit ninexnine_unit_5241(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3901E)
);

ninexnine_unit ninexnine_unit_5242(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A01E)
);

ninexnine_unit ninexnine_unit_5243(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B01E)
);

ninexnine_unit ninexnine_unit_5244(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C01E)
);

ninexnine_unit ninexnine_unit_5245(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D01E)
);

ninexnine_unit ninexnine_unit_5246(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E01E)
);

ninexnine_unit ninexnine_unit_5247(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F01E)
);

assign C301E=c3001E+c3101E+c3201E+c3301E+c3401E+c3501E+c3601E+c3701E+c3801E+c3901E+c3A01E+c3B01E+c3C01E+c3D01E+c3E01E+c3F01E;
assign A301E=(C301E>=0)?1:0;

assign P401E=A301E;

ninexnine_unit ninexnine_unit_5248(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3002E)
);

ninexnine_unit ninexnine_unit_5249(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3102E)
);

ninexnine_unit ninexnine_unit_5250(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3202E)
);

ninexnine_unit ninexnine_unit_5251(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3302E)
);

ninexnine_unit ninexnine_unit_5252(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3402E)
);

ninexnine_unit ninexnine_unit_5253(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3502E)
);

ninexnine_unit ninexnine_unit_5254(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3602E)
);

ninexnine_unit ninexnine_unit_5255(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3702E)
);

ninexnine_unit ninexnine_unit_5256(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3802E)
);

ninexnine_unit ninexnine_unit_5257(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3902E)
);

ninexnine_unit ninexnine_unit_5258(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A02E)
);

ninexnine_unit ninexnine_unit_5259(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B02E)
);

ninexnine_unit ninexnine_unit_5260(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C02E)
);

ninexnine_unit ninexnine_unit_5261(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D02E)
);

ninexnine_unit ninexnine_unit_5262(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E02E)
);

ninexnine_unit ninexnine_unit_5263(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F02E)
);

assign C302E=c3002E+c3102E+c3202E+c3302E+c3402E+c3502E+c3602E+c3702E+c3802E+c3902E+c3A02E+c3B02E+c3C02E+c3D02E+c3E02E+c3F02E;
assign A302E=(C302E>=0)?1:0;

assign P402E=A302E;

ninexnine_unit ninexnine_unit_5264(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3010E)
);

ninexnine_unit ninexnine_unit_5265(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3110E)
);

ninexnine_unit ninexnine_unit_5266(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3210E)
);

ninexnine_unit ninexnine_unit_5267(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3310E)
);

ninexnine_unit ninexnine_unit_5268(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3410E)
);

ninexnine_unit ninexnine_unit_5269(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3510E)
);

ninexnine_unit ninexnine_unit_5270(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3610E)
);

ninexnine_unit ninexnine_unit_5271(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3710E)
);

ninexnine_unit ninexnine_unit_5272(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3810E)
);

ninexnine_unit ninexnine_unit_5273(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3910E)
);

ninexnine_unit ninexnine_unit_5274(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A10E)
);

ninexnine_unit ninexnine_unit_5275(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B10E)
);

ninexnine_unit ninexnine_unit_5276(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C10E)
);

ninexnine_unit ninexnine_unit_5277(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D10E)
);

ninexnine_unit ninexnine_unit_5278(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E10E)
);

ninexnine_unit ninexnine_unit_5279(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F10E)
);

assign C310E=c3010E+c3110E+c3210E+c3310E+c3410E+c3510E+c3610E+c3710E+c3810E+c3910E+c3A10E+c3B10E+c3C10E+c3D10E+c3E10E+c3F10E;
assign A310E=(C310E>=0)?1:0;

assign P410E=A310E;

ninexnine_unit ninexnine_unit_5280(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3011E)
);

ninexnine_unit ninexnine_unit_5281(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3111E)
);

ninexnine_unit ninexnine_unit_5282(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3211E)
);

ninexnine_unit ninexnine_unit_5283(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3311E)
);

ninexnine_unit ninexnine_unit_5284(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3411E)
);

ninexnine_unit ninexnine_unit_5285(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3511E)
);

ninexnine_unit ninexnine_unit_5286(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3611E)
);

ninexnine_unit ninexnine_unit_5287(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3711E)
);

ninexnine_unit ninexnine_unit_5288(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3811E)
);

ninexnine_unit ninexnine_unit_5289(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3911E)
);

ninexnine_unit ninexnine_unit_5290(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A11E)
);

ninexnine_unit ninexnine_unit_5291(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B11E)
);

ninexnine_unit ninexnine_unit_5292(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C11E)
);

ninexnine_unit ninexnine_unit_5293(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D11E)
);

ninexnine_unit ninexnine_unit_5294(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E11E)
);

ninexnine_unit ninexnine_unit_5295(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F11E)
);

assign C311E=c3011E+c3111E+c3211E+c3311E+c3411E+c3511E+c3611E+c3711E+c3811E+c3911E+c3A11E+c3B11E+c3C11E+c3D11E+c3E11E+c3F11E;
assign A311E=(C311E>=0)?1:0;

assign P411E=A311E;

ninexnine_unit ninexnine_unit_5296(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3012E)
);

ninexnine_unit ninexnine_unit_5297(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3112E)
);

ninexnine_unit ninexnine_unit_5298(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3212E)
);

ninexnine_unit ninexnine_unit_5299(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3312E)
);

ninexnine_unit ninexnine_unit_5300(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3412E)
);

ninexnine_unit ninexnine_unit_5301(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3512E)
);

ninexnine_unit ninexnine_unit_5302(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3612E)
);

ninexnine_unit ninexnine_unit_5303(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3712E)
);

ninexnine_unit ninexnine_unit_5304(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3812E)
);

ninexnine_unit ninexnine_unit_5305(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3912E)
);

ninexnine_unit ninexnine_unit_5306(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A12E)
);

ninexnine_unit ninexnine_unit_5307(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B12E)
);

ninexnine_unit ninexnine_unit_5308(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C12E)
);

ninexnine_unit ninexnine_unit_5309(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D12E)
);

ninexnine_unit ninexnine_unit_5310(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E12E)
);

ninexnine_unit ninexnine_unit_5311(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F12E)
);

assign C312E=c3012E+c3112E+c3212E+c3312E+c3412E+c3512E+c3612E+c3712E+c3812E+c3912E+c3A12E+c3B12E+c3C12E+c3D12E+c3E12E+c3F12E;
assign A312E=(C312E>=0)?1:0;

assign P412E=A312E;

ninexnine_unit ninexnine_unit_5312(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3020E)
);

ninexnine_unit ninexnine_unit_5313(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3120E)
);

ninexnine_unit ninexnine_unit_5314(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3220E)
);

ninexnine_unit ninexnine_unit_5315(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3320E)
);

ninexnine_unit ninexnine_unit_5316(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3420E)
);

ninexnine_unit ninexnine_unit_5317(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3520E)
);

ninexnine_unit ninexnine_unit_5318(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3620E)
);

ninexnine_unit ninexnine_unit_5319(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3720E)
);

ninexnine_unit ninexnine_unit_5320(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3820E)
);

ninexnine_unit ninexnine_unit_5321(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3920E)
);

ninexnine_unit ninexnine_unit_5322(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A20E)
);

ninexnine_unit ninexnine_unit_5323(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B20E)
);

ninexnine_unit ninexnine_unit_5324(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C20E)
);

ninexnine_unit ninexnine_unit_5325(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D20E)
);

ninexnine_unit ninexnine_unit_5326(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E20E)
);

ninexnine_unit ninexnine_unit_5327(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F20E)
);

assign C320E=c3020E+c3120E+c3220E+c3320E+c3420E+c3520E+c3620E+c3720E+c3820E+c3920E+c3A20E+c3B20E+c3C20E+c3D20E+c3E20E+c3F20E;
assign A320E=(C320E>=0)?1:0;

assign P420E=A320E;

ninexnine_unit ninexnine_unit_5328(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3021E)
);

ninexnine_unit ninexnine_unit_5329(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3121E)
);

ninexnine_unit ninexnine_unit_5330(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3221E)
);

ninexnine_unit ninexnine_unit_5331(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3321E)
);

ninexnine_unit ninexnine_unit_5332(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3421E)
);

ninexnine_unit ninexnine_unit_5333(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3521E)
);

ninexnine_unit ninexnine_unit_5334(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3621E)
);

ninexnine_unit ninexnine_unit_5335(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3721E)
);

ninexnine_unit ninexnine_unit_5336(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3821E)
);

ninexnine_unit ninexnine_unit_5337(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3921E)
);

ninexnine_unit ninexnine_unit_5338(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A21E)
);

ninexnine_unit ninexnine_unit_5339(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B21E)
);

ninexnine_unit ninexnine_unit_5340(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C21E)
);

ninexnine_unit ninexnine_unit_5341(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D21E)
);

ninexnine_unit ninexnine_unit_5342(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E21E)
);

ninexnine_unit ninexnine_unit_5343(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F21E)
);

assign C321E=c3021E+c3121E+c3221E+c3321E+c3421E+c3521E+c3621E+c3721E+c3821E+c3921E+c3A21E+c3B21E+c3C21E+c3D21E+c3E21E+c3F21E;
assign A321E=(C321E>=0)?1:0;

assign P421E=A321E;

ninexnine_unit ninexnine_unit_5344(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3E000),
				.b1(W3E010),
				.b2(W3E020),
				.b3(W3E100),
				.b4(W3E110),
				.b5(W3E120),
				.b6(W3E200),
				.b7(W3E210),
				.b8(W3E220),
				.c(c3022E)
);

ninexnine_unit ninexnine_unit_5345(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3E001),
				.b1(W3E011),
				.b2(W3E021),
				.b3(W3E101),
				.b4(W3E111),
				.b5(W3E121),
				.b6(W3E201),
				.b7(W3E211),
				.b8(W3E221),
				.c(c3122E)
);

ninexnine_unit ninexnine_unit_5346(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3E002),
				.b1(W3E012),
				.b2(W3E022),
				.b3(W3E102),
				.b4(W3E112),
				.b5(W3E122),
				.b6(W3E202),
				.b7(W3E212),
				.b8(W3E222),
				.c(c3222E)
);

ninexnine_unit ninexnine_unit_5347(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3E003),
				.b1(W3E013),
				.b2(W3E023),
				.b3(W3E103),
				.b4(W3E113),
				.b5(W3E123),
				.b6(W3E203),
				.b7(W3E213),
				.b8(W3E223),
				.c(c3322E)
);

ninexnine_unit ninexnine_unit_5348(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3E004),
				.b1(W3E014),
				.b2(W3E024),
				.b3(W3E104),
				.b4(W3E114),
				.b5(W3E124),
				.b6(W3E204),
				.b7(W3E214),
				.b8(W3E224),
				.c(c3422E)
);

ninexnine_unit ninexnine_unit_5349(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3E005),
				.b1(W3E015),
				.b2(W3E025),
				.b3(W3E105),
				.b4(W3E115),
				.b5(W3E125),
				.b6(W3E205),
				.b7(W3E215),
				.b8(W3E225),
				.c(c3522E)
);

ninexnine_unit ninexnine_unit_5350(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3E006),
				.b1(W3E016),
				.b2(W3E026),
				.b3(W3E106),
				.b4(W3E116),
				.b5(W3E126),
				.b6(W3E206),
				.b7(W3E216),
				.b8(W3E226),
				.c(c3622E)
);

ninexnine_unit ninexnine_unit_5351(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3E007),
				.b1(W3E017),
				.b2(W3E027),
				.b3(W3E107),
				.b4(W3E117),
				.b5(W3E127),
				.b6(W3E207),
				.b7(W3E217),
				.b8(W3E227),
				.c(c3722E)
);

ninexnine_unit ninexnine_unit_5352(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3E008),
				.b1(W3E018),
				.b2(W3E028),
				.b3(W3E108),
				.b4(W3E118),
				.b5(W3E128),
				.b6(W3E208),
				.b7(W3E218),
				.b8(W3E228),
				.c(c3822E)
);

ninexnine_unit ninexnine_unit_5353(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3E009),
				.b1(W3E019),
				.b2(W3E029),
				.b3(W3E109),
				.b4(W3E119),
				.b5(W3E129),
				.b6(W3E209),
				.b7(W3E219),
				.b8(W3E229),
				.c(c3922E)
);

ninexnine_unit ninexnine_unit_5354(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3E00A),
				.b1(W3E01A),
				.b2(W3E02A),
				.b3(W3E10A),
				.b4(W3E11A),
				.b5(W3E12A),
				.b6(W3E20A),
				.b7(W3E21A),
				.b8(W3E22A),
				.c(c3A22E)
);

ninexnine_unit ninexnine_unit_5355(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3E00B),
				.b1(W3E01B),
				.b2(W3E02B),
				.b3(W3E10B),
				.b4(W3E11B),
				.b5(W3E12B),
				.b6(W3E20B),
				.b7(W3E21B),
				.b8(W3E22B),
				.c(c3B22E)
);

ninexnine_unit ninexnine_unit_5356(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3E00C),
				.b1(W3E01C),
				.b2(W3E02C),
				.b3(W3E10C),
				.b4(W3E11C),
				.b5(W3E12C),
				.b6(W3E20C),
				.b7(W3E21C),
				.b8(W3E22C),
				.c(c3C22E)
);

ninexnine_unit ninexnine_unit_5357(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3E00D),
				.b1(W3E01D),
				.b2(W3E02D),
				.b3(W3E10D),
				.b4(W3E11D),
				.b5(W3E12D),
				.b6(W3E20D),
				.b7(W3E21D),
				.b8(W3E22D),
				.c(c3D22E)
);

ninexnine_unit ninexnine_unit_5358(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3E00E),
				.b1(W3E01E),
				.b2(W3E02E),
				.b3(W3E10E),
				.b4(W3E11E),
				.b5(W3E12E),
				.b6(W3E20E),
				.b7(W3E21E),
				.b8(W3E22E),
				.c(c3E22E)
);

ninexnine_unit ninexnine_unit_5359(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3E00F),
				.b1(W3E01F),
				.b2(W3E02F),
				.b3(W3E10F),
				.b4(W3E11F),
				.b5(W3E12F),
				.b6(W3E20F),
				.b7(W3E21F),
				.b8(W3E22F),
				.c(c3F22E)
);

assign C322E=c3022E+c3122E+c3222E+c3322E+c3422E+c3522E+c3622E+c3722E+c3822E+c3922E+c3A22E+c3B22E+c3C22E+c3D22E+c3E22E+c3F22E;
assign A322E=(C322E>=0)?1:0;

assign P422E=A322E;

ninexnine_unit ninexnine_unit_5360(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3000F)
);

ninexnine_unit ninexnine_unit_5361(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3100F)
);

ninexnine_unit ninexnine_unit_5362(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3200F)
);

ninexnine_unit ninexnine_unit_5363(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3300F)
);

ninexnine_unit ninexnine_unit_5364(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3400F)
);

ninexnine_unit ninexnine_unit_5365(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3500F)
);

ninexnine_unit ninexnine_unit_5366(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3600F)
);

ninexnine_unit ninexnine_unit_5367(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3700F)
);

ninexnine_unit ninexnine_unit_5368(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3800F)
);

ninexnine_unit ninexnine_unit_5369(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3900F)
);

ninexnine_unit ninexnine_unit_5370(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A00F)
);

ninexnine_unit ninexnine_unit_5371(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B00F)
);

ninexnine_unit ninexnine_unit_5372(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C00F)
);

ninexnine_unit ninexnine_unit_5373(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D00F)
);

ninexnine_unit ninexnine_unit_5374(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E00F)
);

ninexnine_unit ninexnine_unit_5375(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F00F)
);

assign C300F=c3000F+c3100F+c3200F+c3300F+c3400F+c3500F+c3600F+c3700F+c3800F+c3900F+c3A00F+c3B00F+c3C00F+c3D00F+c3E00F+c3F00F;
assign A300F=(C300F>=0)?1:0;

assign P400F=A300F;

ninexnine_unit ninexnine_unit_5376(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3001F)
);

ninexnine_unit ninexnine_unit_5377(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3101F)
);

ninexnine_unit ninexnine_unit_5378(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3201F)
);

ninexnine_unit ninexnine_unit_5379(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3301F)
);

ninexnine_unit ninexnine_unit_5380(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3401F)
);

ninexnine_unit ninexnine_unit_5381(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3501F)
);

ninexnine_unit ninexnine_unit_5382(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3601F)
);

ninexnine_unit ninexnine_unit_5383(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3701F)
);

ninexnine_unit ninexnine_unit_5384(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3801F)
);

ninexnine_unit ninexnine_unit_5385(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3901F)
);

ninexnine_unit ninexnine_unit_5386(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A01F)
);

ninexnine_unit ninexnine_unit_5387(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B01F)
);

ninexnine_unit ninexnine_unit_5388(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C01F)
);

ninexnine_unit ninexnine_unit_5389(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D01F)
);

ninexnine_unit ninexnine_unit_5390(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E01F)
);

ninexnine_unit ninexnine_unit_5391(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F01F)
);

assign C301F=c3001F+c3101F+c3201F+c3301F+c3401F+c3501F+c3601F+c3701F+c3801F+c3901F+c3A01F+c3B01F+c3C01F+c3D01F+c3E01F+c3F01F;
assign A301F=(C301F>=0)?1:0;

assign P401F=A301F;

ninexnine_unit ninexnine_unit_5392(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3002F)
);

ninexnine_unit ninexnine_unit_5393(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3102F)
);

ninexnine_unit ninexnine_unit_5394(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3202F)
);

ninexnine_unit ninexnine_unit_5395(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3302F)
);

ninexnine_unit ninexnine_unit_5396(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3402F)
);

ninexnine_unit ninexnine_unit_5397(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3502F)
);

ninexnine_unit ninexnine_unit_5398(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3602F)
);

ninexnine_unit ninexnine_unit_5399(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3702F)
);

ninexnine_unit ninexnine_unit_5400(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3802F)
);

ninexnine_unit ninexnine_unit_5401(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3902F)
);

ninexnine_unit ninexnine_unit_5402(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A02F)
);

ninexnine_unit ninexnine_unit_5403(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B02F)
);

ninexnine_unit ninexnine_unit_5404(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C02F)
);

ninexnine_unit ninexnine_unit_5405(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D02F)
);

ninexnine_unit ninexnine_unit_5406(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E02F)
);

ninexnine_unit ninexnine_unit_5407(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F02F)
);

assign C302F=c3002F+c3102F+c3202F+c3302F+c3402F+c3502F+c3602F+c3702F+c3802F+c3902F+c3A02F+c3B02F+c3C02F+c3D02F+c3E02F+c3F02F;
assign A302F=(C302F>=0)?1:0;

assign P402F=A302F;

ninexnine_unit ninexnine_unit_5408(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3010F)
);

ninexnine_unit ninexnine_unit_5409(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3110F)
);

ninexnine_unit ninexnine_unit_5410(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3210F)
);

ninexnine_unit ninexnine_unit_5411(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3310F)
);

ninexnine_unit ninexnine_unit_5412(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3410F)
);

ninexnine_unit ninexnine_unit_5413(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3510F)
);

ninexnine_unit ninexnine_unit_5414(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3610F)
);

ninexnine_unit ninexnine_unit_5415(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3710F)
);

ninexnine_unit ninexnine_unit_5416(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3810F)
);

ninexnine_unit ninexnine_unit_5417(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3910F)
);

ninexnine_unit ninexnine_unit_5418(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A10F)
);

ninexnine_unit ninexnine_unit_5419(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B10F)
);

ninexnine_unit ninexnine_unit_5420(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C10F)
);

ninexnine_unit ninexnine_unit_5421(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D10F)
);

ninexnine_unit ninexnine_unit_5422(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E10F)
);

ninexnine_unit ninexnine_unit_5423(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F10F)
);

assign C310F=c3010F+c3110F+c3210F+c3310F+c3410F+c3510F+c3610F+c3710F+c3810F+c3910F+c3A10F+c3B10F+c3C10F+c3D10F+c3E10F+c3F10F;
assign A310F=(C310F>=0)?1:0;

assign P410F=A310F;

ninexnine_unit ninexnine_unit_5424(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3011F)
);

ninexnine_unit ninexnine_unit_5425(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3111F)
);

ninexnine_unit ninexnine_unit_5426(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3211F)
);

ninexnine_unit ninexnine_unit_5427(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3311F)
);

ninexnine_unit ninexnine_unit_5428(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3411F)
);

ninexnine_unit ninexnine_unit_5429(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3511F)
);

ninexnine_unit ninexnine_unit_5430(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3611F)
);

ninexnine_unit ninexnine_unit_5431(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3711F)
);

ninexnine_unit ninexnine_unit_5432(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3811F)
);

ninexnine_unit ninexnine_unit_5433(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3911F)
);

ninexnine_unit ninexnine_unit_5434(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A11F)
);

ninexnine_unit ninexnine_unit_5435(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B11F)
);

ninexnine_unit ninexnine_unit_5436(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C11F)
);

ninexnine_unit ninexnine_unit_5437(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D11F)
);

ninexnine_unit ninexnine_unit_5438(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E11F)
);

ninexnine_unit ninexnine_unit_5439(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F11F)
);

assign C311F=c3011F+c3111F+c3211F+c3311F+c3411F+c3511F+c3611F+c3711F+c3811F+c3911F+c3A11F+c3B11F+c3C11F+c3D11F+c3E11F+c3F11F;
assign A311F=(C311F>=0)?1:0;

assign P411F=A311F;

ninexnine_unit ninexnine_unit_5440(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3012F)
);

ninexnine_unit ninexnine_unit_5441(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3112F)
);

ninexnine_unit ninexnine_unit_5442(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3212F)
);

ninexnine_unit ninexnine_unit_5443(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3312F)
);

ninexnine_unit ninexnine_unit_5444(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3412F)
);

ninexnine_unit ninexnine_unit_5445(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3512F)
);

ninexnine_unit ninexnine_unit_5446(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3612F)
);

ninexnine_unit ninexnine_unit_5447(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3712F)
);

ninexnine_unit ninexnine_unit_5448(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3812F)
);

ninexnine_unit ninexnine_unit_5449(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3912F)
);

ninexnine_unit ninexnine_unit_5450(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A12F)
);

ninexnine_unit ninexnine_unit_5451(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B12F)
);

ninexnine_unit ninexnine_unit_5452(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C12F)
);

ninexnine_unit ninexnine_unit_5453(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D12F)
);

ninexnine_unit ninexnine_unit_5454(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E12F)
);

ninexnine_unit ninexnine_unit_5455(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F12F)
);

assign C312F=c3012F+c3112F+c3212F+c3312F+c3412F+c3512F+c3612F+c3712F+c3812F+c3912F+c3A12F+c3B12F+c3C12F+c3D12F+c3E12F+c3F12F;
assign A312F=(C312F>=0)?1:0;

assign P412F=A312F;

ninexnine_unit ninexnine_unit_5456(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3020F)
);

ninexnine_unit ninexnine_unit_5457(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3120F)
);

ninexnine_unit ninexnine_unit_5458(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3220F)
);

ninexnine_unit ninexnine_unit_5459(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3320F)
);

ninexnine_unit ninexnine_unit_5460(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3420F)
);

ninexnine_unit ninexnine_unit_5461(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3520F)
);

ninexnine_unit ninexnine_unit_5462(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3620F)
);

ninexnine_unit ninexnine_unit_5463(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3720F)
);

ninexnine_unit ninexnine_unit_5464(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3820F)
);

ninexnine_unit ninexnine_unit_5465(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3920F)
);

ninexnine_unit ninexnine_unit_5466(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A20F)
);

ninexnine_unit ninexnine_unit_5467(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B20F)
);

ninexnine_unit ninexnine_unit_5468(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C20F)
);

ninexnine_unit ninexnine_unit_5469(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D20F)
);

ninexnine_unit ninexnine_unit_5470(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E20F)
);

ninexnine_unit ninexnine_unit_5471(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F20F)
);

assign C320F=c3020F+c3120F+c3220F+c3320F+c3420F+c3520F+c3620F+c3720F+c3820F+c3920F+c3A20F+c3B20F+c3C20F+c3D20F+c3E20F+c3F20F;
assign A320F=(C320F>=0)?1:0;

assign P420F=A320F;

ninexnine_unit ninexnine_unit_5472(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3021F)
);

ninexnine_unit ninexnine_unit_5473(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3121F)
);

ninexnine_unit ninexnine_unit_5474(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3221F)
);

ninexnine_unit ninexnine_unit_5475(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3321F)
);

ninexnine_unit ninexnine_unit_5476(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3421F)
);

ninexnine_unit ninexnine_unit_5477(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3521F)
);

ninexnine_unit ninexnine_unit_5478(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3621F)
);

ninexnine_unit ninexnine_unit_5479(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3721F)
);

ninexnine_unit ninexnine_unit_5480(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3821F)
);

ninexnine_unit ninexnine_unit_5481(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3921F)
);

ninexnine_unit ninexnine_unit_5482(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A21F)
);

ninexnine_unit ninexnine_unit_5483(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B21F)
);

ninexnine_unit ninexnine_unit_5484(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C21F)
);

ninexnine_unit ninexnine_unit_5485(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D21F)
);

ninexnine_unit ninexnine_unit_5486(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E21F)
);

ninexnine_unit ninexnine_unit_5487(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F21F)
);

assign C321F=c3021F+c3121F+c3221F+c3321F+c3421F+c3521F+c3621F+c3721F+c3821F+c3921F+c3A21F+c3B21F+c3C21F+c3D21F+c3E21F+c3F21F;
assign A321F=(C321F>=0)?1:0;

assign P421F=A321F;

ninexnine_unit ninexnine_unit_5488(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3F000),
				.b1(W3F010),
				.b2(W3F020),
				.b3(W3F100),
				.b4(W3F110),
				.b5(W3F120),
				.b6(W3F200),
				.b7(W3F210),
				.b8(W3F220),
				.c(c3022F)
);

ninexnine_unit ninexnine_unit_5489(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3F001),
				.b1(W3F011),
				.b2(W3F021),
				.b3(W3F101),
				.b4(W3F111),
				.b5(W3F121),
				.b6(W3F201),
				.b7(W3F211),
				.b8(W3F221),
				.c(c3122F)
);

ninexnine_unit ninexnine_unit_5490(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3F002),
				.b1(W3F012),
				.b2(W3F022),
				.b3(W3F102),
				.b4(W3F112),
				.b5(W3F122),
				.b6(W3F202),
				.b7(W3F212),
				.b8(W3F222),
				.c(c3222F)
);

ninexnine_unit ninexnine_unit_5491(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3F003),
				.b1(W3F013),
				.b2(W3F023),
				.b3(W3F103),
				.b4(W3F113),
				.b5(W3F123),
				.b6(W3F203),
				.b7(W3F213),
				.b8(W3F223),
				.c(c3322F)
);

ninexnine_unit ninexnine_unit_5492(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3F004),
				.b1(W3F014),
				.b2(W3F024),
				.b3(W3F104),
				.b4(W3F114),
				.b5(W3F124),
				.b6(W3F204),
				.b7(W3F214),
				.b8(W3F224),
				.c(c3422F)
);

ninexnine_unit ninexnine_unit_5493(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3F005),
				.b1(W3F015),
				.b2(W3F025),
				.b3(W3F105),
				.b4(W3F115),
				.b5(W3F125),
				.b6(W3F205),
				.b7(W3F215),
				.b8(W3F225),
				.c(c3522F)
);

ninexnine_unit ninexnine_unit_5494(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3F006),
				.b1(W3F016),
				.b2(W3F026),
				.b3(W3F106),
				.b4(W3F116),
				.b5(W3F126),
				.b6(W3F206),
				.b7(W3F216),
				.b8(W3F226),
				.c(c3622F)
);

ninexnine_unit ninexnine_unit_5495(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3F007),
				.b1(W3F017),
				.b2(W3F027),
				.b3(W3F107),
				.b4(W3F117),
				.b5(W3F127),
				.b6(W3F207),
				.b7(W3F217),
				.b8(W3F227),
				.c(c3722F)
);

ninexnine_unit ninexnine_unit_5496(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3F008),
				.b1(W3F018),
				.b2(W3F028),
				.b3(W3F108),
				.b4(W3F118),
				.b5(W3F128),
				.b6(W3F208),
				.b7(W3F218),
				.b8(W3F228),
				.c(c3822F)
);

ninexnine_unit ninexnine_unit_5497(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3F009),
				.b1(W3F019),
				.b2(W3F029),
				.b3(W3F109),
				.b4(W3F119),
				.b5(W3F129),
				.b6(W3F209),
				.b7(W3F219),
				.b8(W3F229),
				.c(c3922F)
);

ninexnine_unit ninexnine_unit_5498(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3F00A),
				.b1(W3F01A),
				.b2(W3F02A),
				.b3(W3F10A),
				.b4(W3F11A),
				.b5(W3F12A),
				.b6(W3F20A),
				.b7(W3F21A),
				.b8(W3F22A),
				.c(c3A22F)
);

ninexnine_unit ninexnine_unit_5499(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3F00B),
				.b1(W3F01B),
				.b2(W3F02B),
				.b3(W3F10B),
				.b4(W3F11B),
				.b5(W3F12B),
				.b6(W3F20B),
				.b7(W3F21B),
				.b8(W3F22B),
				.c(c3B22F)
);

ninexnine_unit ninexnine_unit_5500(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3F00C),
				.b1(W3F01C),
				.b2(W3F02C),
				.b3(W3F10C),
				.b4(W3F11C),
				.b5(W3F12C),
				.b6(W3F20C),
				.b7(W3F21C),
				.b8(W3F22C),
				.c(c3C22F)
);

ninexnine_unit ninexnine_unit_5501(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3F00D),
				.b1(W3F01D),
				.b2(W3F02D),
				.b3(W3F10D),
				.b4(W3F11D),
				.b5(W3F12D),
				.b6(W3F20D),
				.b7(W3F21D),
				.b8(W3F22D),
				.c(c3D22F)
);

ninexnine_unit ninexnine_unit_5502(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3F00E),
				.b1(W3F01E),
				.b2(W3F02E),
				.b3(W3F10E),
				.b4(W3F11E),
				.b5(W3F12E),
				.b6(W3F20E),
				.b7(W3F21E),
				.b8(W3F22E),
				.c(c3E22F)
);

ninexnine_unit ninexnine_unit_5503(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3F00F),
				.b1(W3F01F),
				.b2(W3F02F),
				.b3(W3F10F),
				.b4(W3F11F),
				.b5(W3F12F),
				.b6(W3F20F),
				.b7(W3F21F),
				.b8(W3F22F),
				.c(c3F22F)
);

assign C322F=c3022F+c3122F+c3222F+c3322F+c3422F+c3522F+c3622F+c3722F+c3822F+c3922F+c3A22F+c3B22F+c3C22F+c3D22F+c3E22F+c3F22F;
assign A322F=(C322F>=0)?1:0;

assign P422F=A322F;

ninexnine_unit ninexnine_unit_5504(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3000G)
);

ninexnine_unit ninexnine_unit_5505(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3100G)
);

ninexnine_unit ninexnine_unit_5506(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3200G)
);

ninexnine_unit ninexnine_unit_5507(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3300G)
);

ninexnine_unit ninexnine_unit_5508(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3400G)
);

ninexnine_unit ninexnine_unit_5509(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3500G)
);

ninexnine_unit ninexnine_unit_5510(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3600G)
);

ninexnine_unit ninexnine_unit_5511(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3700G)
);

ninexnine_unit ninexnine_unit_5512(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3800G)
);

ninexnine_unit ninexnine_unit_5513(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3900G)
);

ninexnine_unit ninexnine_unit_5514(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A00G)
);

ninexnine_unit ninexnine_unit_5515(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B00G)
);

ninexnine_unit ninexnine_unit_5516(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C00G)
);

ninexnine_unit ninexnine_unit_5517(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D00G)
);

ninexnine_unit ninexnine_unit_5518(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E00G)
);

ninexnine_unit ninexnine_unit_5519(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F00G)
);

assign C300G=c3000G+c3100G+c3200G+c3300G+c3400G+c3500G+c3600G+c3700G+c3800G+c3900G+c3A00G+c3B00G+c3C00G+c3D00G+c3E00G+c3F00G;
assign A300G=(C300G>=0)?1:0;

assign P400G=A300G;

ninexnine_unit ninexnine_unit_5520(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3001G)
);

ninexnine_unit ninexnine_unit_5521(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3101G)
);

ninexnine_unit ninexnine_unit_5522(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3201G)
);

ninexnine_unit ninexnine_unit_5523(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3301G)
);

ninexnine_unit ninexnine_unit_5524(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3401G)
);

ninexnine_unit ninexnine_unit_5525(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3501G)
);

ninexnine_unit ninexnine_unit_5526(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3601G)
);

ninexnine_unit ninexnine_unit_5527(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3701G)
);

ninexnine_unit ninexnine_unit_5528(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3801G)
);

ninexnine_unit ninexnine_unit_5529(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3901G)
);

ninexnine_unit ninexnine_unit_5530(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A01G)
);

ninexnine_unit ninexnine_unit_5531(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B01G)
);

ninexnine_unit ninexnine_unit_5532(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C01G)
);

ninexnine_unit ninexnine_unit_5533(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D01G)
);

ninexnine_unit ninexnine_unit_5534(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E01G)
);

ninexnine_unit ninexnine_unit_5535(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F01G)
);

assign C301G=c3001G+c3101G+c3201G+c3301G+c3401G+c3501G+c3601G+c3701G+c3801G+c3901G+c3A01G+c3B01G+c3C01G+c3D01G+c3E01G+c3F01G;
assign A301G=(C301G>=0)?1:0;

assign P401G=A301G;

ninexnine_unit ninexnine_unit_5536(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3002G)
);

ninexnine_unit ninexnine_unit_5537(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3102G)
);

ninexnine_unit ninexnine_unit_5538(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3202G)
);

ninexnine_unit ninexnine_unit_5539(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3302G)
);

ninexnine_unit ninexnine_unit_5540(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3402G)
);

ninexnine_unit ninexnine_unit_5541(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3502G)
);

ninexnine_unit ninexnine_unit_5542(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3602G)
);

ninexnine_unit ninexnine_unit_5543(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3702G)
);

ninexnine_unit ninexnine_unit_5544(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3802G)
);

ninexnine_unit ninexnine_unit_5545(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3902G)
);

ninexnine_unit ninexnine_unit_5546(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A02G)
);

ninexnine_unit ninexnine_unit_5547(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B02G)
);

ninexnine_unit ninexnine_unit_5548(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C02G)
);

ninexnine_unit ninexnine_unit_5549(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D02G)
);

ninexnine_unit ninexnine_unit_5550(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E02G)
);

ninexnine_unit ninexnine_unit_5551(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F02G)
);

assign C302G=c3002G+c3102G+c3202G+c3302G+c3402G+c3502G+c3602G+c3702G+c3802G+c3902G+c3A02G+c3B02G+c3C02G+c3D02G+c3E02G+c3F02G;
assign A302G=(C302G>=0)?1:0;

assign P402G=A302G;

ninexnine_unit ninexnine_unit_5552(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3010G)
);

ninexnine_unit ninexnine_unit_5553(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3110G)
);

ninexnine_unit ninexnine_unit_5554(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3210G)
);

ninexnine_unit ninexnine_unit_5555(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3310G)
);

ninexnine_unit ninexnine_unit_5556(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3410G)
);

ninexnine_unit ninexnine_unit_5557(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3510G)
);

ninexnine_unit ninexnine_unit_5558(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3610G)
);

ninexnine_unit ninexnine_unit_5559(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3710G)
);

ninexnine_unit ninexnine_unit_5560(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3810G)
);

ninexnine_unit ninexnine_unit_5561(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3910G)
);

ninexnine_unit ninexnine_unit_5562(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A10G)
);

ninexnine_unit ninexnine_unit_5563(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B10G)
);

ninexnine_unit ninexnine_unit_5564(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C10G)
);

ninexnine_unit ninexnine_unit_5565(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D10G)
);

ninexnine_unit ninexnine_unit_5566(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E10G)
);

ninexnine_unit ninexnine_unit_5567(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F10G)
);

assign C310G=c3010G+c3110G+c3210G+c3310G+c3410G+c3510G+c3610G+c3710G+c3810G+c3910G+c3A10G+c3B10G+c3C10G+c3D10G+c3E10G+c3F10G;
assign A310G=(C310G>=0)?1:0;

assign P410G=A310G;

ninexnine_unit ninexnine_unit_5568(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3011G)
);

ninexnine_unit ninexnine_unit_5569(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3111G)
);

ninexnine_unit ninexnine_unit_5570(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3211G)
);

ninexnine_unit ninexnine_unit_5571(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3311G)
);

ninexnine_unit ninexnine_unit_5572(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3411G)
);

ninexnine_unit ninexnine_unit_5573(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3511G)
);

ninexnine_unit ninexnine_unit_5574(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3611G)
);

ninexnine_unit ninexnine_unit_5575(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3711G)
);

ninexnine_unit ninexnine_unit_5576(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3811G)
);

ninexnine_unit ninexnine_unit_5577(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3911G)
);

ninexnine_unit ninexnine_unit_5578(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A11G)
);

ninexnine_unit ninexnine_unit_5579(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B11G)
);

ninexnine_unit ninexnine_unit_5580(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C11G)
);

ninexnine_unit ninexnine_unit_5581(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D11G)
);

ninexnine_unit ninexnine_unit_5582(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E11G)
);

ninexnine_unit ninexnine_unit_5583(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F11G)
);

assign C311G=c3011G+c3111G+c3211G+c3311G+c3411G+c3511G+c3611G+c3711G+c3811G+c3911G+c3A11G+c3B11G+c3C11G+c3D11G+c3E11G+c3F11G;
assign A311G=(C311G>=0)?1:0;

assign P411G=A311G;

ninexnine_unit ninexnine_unit_5584(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3012G)
);

ninexnine_unit ninexnine_unit_5585(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3112G)
);

ninexnine_unit ninexnine_unit_5586(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3212G)
);

ninexnine_unit ninexnine_unit_5587(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3312G)
);

ninexnine_unit ninexnine_unit_5588(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3412G)
);

ninexnine_unit ninexnine_unit_5589(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3512G)
);

ninexnine_unit ninexnine_unit_5590(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3612G)
);

ninexnine_unit ninexnine_unit_5591(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3712G)
);

ninexnine_unit ninexnine_unit_5592(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3812G)
);

ninexnine_unit ninexnine_unit_5593(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3912G)
);

ninexnine_unit ninexnine_unit_5594(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A12G)
);

ninexnine_unit ninexnine_unit_5595(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B12G)
);

ninexnine_unit ninexnine_unit_5596(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C12G)
);

ninexnine_unit ninexnine_unit_5597(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D12G)
);

ninexnine_unit ninexnine_unit_5598(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E12G)
);

ninexnine_unit ninexnine_unit_5599(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F12G)
);

assign C312G=c3012G+c3112G+c3212G+c3312G+c3412G+c3512G+c3612G+c3712G+c3812G+c3912G+c3A12G+c3B12G+c3C12G+c3D12G+c3E12G+c3F12G;
assign A312G=(C312G>=0)?1:0;

assign P412G=A312G;

ninexnine_unit ninexnine_unit_5600(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3020G)
);

ninexnine_unit ninexnine_unit_5601(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3120G)
);

ninexnine_unit ninexnine_unit_5602(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3220G)
);

ninexnine_unit ninexnine_unit_5603(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3320G)
);

ninexnine_unit ninexnine_unit_5604(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3420G)
);

ninexnine_unit ninexnine_unit_5605(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3520G)
);

ninexnine_unit ninexnine_unit_5606(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3620G)
);

ninexnine_unit ninexnine_unit_5607(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3720G)
);

ninexnine_unit ninexnine_unit_5608(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3820G)
);

ninexnine_unit ninexnine_unit_5609(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3920G)
);

ninexnine_unit ninexnine_unit_5610(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A20G)
);

ninexnine_unit ninexnine_unit_5611(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B20G)
);

ninexnine_unit ninexnine_unit_5612(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C20G)
);

ninexnine_unit ninexnine_unit_5613(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D20G)
);

ninexnine_unit ninexnine_unit_5614(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E20G)
);

ninexnine_unit ninexnine_unit_5615(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F20G)
);

assign C320G=c3020G+c3120G+c3220G+c3320G+c3420G+c3520G+c3620G+c3720G+c3820G+c3920G+c3A20G+c3B20G+c3C20G+c3D20G+c3E20G+c3F20G;
assign A320G=(C320G>=0)?1:0;

assign P420G=A320G;

ninexnine_unit ninexnine_unit_5616(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3021G)
);

ninexnine_unit ninexnine_unit_5617(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3121G)
);

ninexnine_unit ninexnine_unit_5618(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3221G)
);

ninexnine_unit ninexnine_unit_5619(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3321G)
);

ninexnine_unit ninexnine_unit_5620(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3421G)
);

ninexnine_unit ninexnine_unit_5621(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3521G)
);

ninexnine_unit ninexnine_unit_5622(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3621G)
);

ninexnine_unit ninexnine_unit_5623(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3721G)
);

ninexnine_unit ninexnine_unit_5624(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3821G)
);

ninexnine_unit ninexnine_unit_5625(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3921G)
);

ninexnine_unit ninexnine_unit_5626(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A21G)
);

ninexnine_unit ninexnine_unit_5627(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B21G)
);

ninexnine_unit ninexnine_unit_5628(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C21G)
);

ninexnine_unit ninexnine_unit_5629(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D21G)
);

ninexnine_unit ninexnine_unit_5630(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E21G)
);

ninexnine_unit ninexnine_unit_5631(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F21G)
);

assign C321G=c3021G+c3121G+c3221G+c3321G+c3421G+c3521G+c3621G+c3721G+c3821G+c3921G+c3A21G+c3B21G+c3C21G+c3D21G+c3E21G+c3F21G;
assign A321G=(C321G>=0)?1:0;

assign P421G=A321G;

ninexnine_unit ninexnine_unit_5632(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3G000),
				.b1(W3G010),
				.b2(W3G020),
				.b3(W3G100),
				.b4(W3G110),
				.b5(W3G120),
				.b6(W3G200),
				.b7(W3G210),
				.b8(W3G220),
				.c(c3022G)
);

ninexnine_unit ninexnine_unit_5633(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3G001),
				.b1(W3G011),
				.b2(W3G021),
				.b3(W3G101),
				.b4(W3G111),
				.b5(W3G121),
				.b6(W3G201),
				.b7(W3G211),
				.b8(W3G221),
				.c(c3122G)
);

ninexnine_unit ninexnine_unit_5634(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3G002),
				.b1(W3G012),
				.b2(W3G022),
				.b3(W3G102),
				.b4(W3G112),
				.b5(W3G122),
				.b6(W3G202),
				.b7(W3G212),
				.b8(W3G222),
				.c(c3222G)
);

ninexnine_unit ninexnine_unit_5635(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3G003),
				.b1(W3G013),
				.b2(W3G023),
				.b3(W3G103),
				.b4(W3G113),
				.b5(W3G123),
				.b6(W3G203),
				.b7(W3G213),
				.b8(W3G223),
				.c(c3322G)
);

ninexnine_unit ninexnine_unit_5636(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3G004),
				.b1(W3G014),
				.b2(W3G024),
				.b3(W3G104),
				.b4(W3G114),
				.b5(W3G124),
				.b6(W3G204),
				.b7(W3G214),
				.b8(W3G224),
				.c(c3422G)
);

ninexnine_unit ninexnine_unit_5637(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3G005),
				.b1(W3G015),
				.b2(W3G025),
				.b3(W3G105),
				.b4(W3G115),
				.b5(W3G125),
				.b6(W3G205),
				.b7(W3G215),
				.b8(W3G225),
				.c(c3522G)
);

ninexnine_unit ninexnine_unit_5638(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3G006),
				.b1(W3G016),
				.b2(W3G026),
				.b3(W3G106),
				.b4(W3G116),
				.b5(W3G126),
				.b6(W3G206),
				.b7(W3G216),
				.b8(W3G226),
				.c(c3622G)
);

ninexnine_unit ninexnine_unit_5639(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3G007),
				.b1(W3G017),
				.b2(W3G027),
				.b3(W3G107),
				.b4(W3G117),
				.b5(W3G127),
				.b6(W3G207),
				.b7(W3G217),
				.b8(W3G227),
				.c(c3722G)
);

ninexnine_unit ninexnine_unit_5640(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3G008),
				.b1(W3G018),
				.b2(W3G028),
				.b3(W3G108),
				.b4(W3G118),
				.b5(W3G128),
				.b6(W3G208),
				.b7(W3G218),
				.b8(W3G228),
				.c(c3822G)
);

ninexnine_unit ninexnine_unit_5641(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3G009),
				.b1(W3G019),
				.b2(W3G029),
				.b3(W3G109),
				.b4(W3G119),
				.b5(W3G129),
				.b6(W3G209),
				.b7(W3G219),
				.b8(W3G229),
				.c(c3922G)
);

ninexnine_unit ninexnine_unit_5642(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3G00A),
				.b1(W3G01A),
				.b2(W3G02A),
				.b3(W3G10A),
				.b4(W3G11A),
				.b5(W3G12A),
				.b6(W3G20A),
				.b7(W3G21A),
				.b8(W3G22A),
				.c(c3A22G)
);

ninexnine_unit ninexnine_unit_5643(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3G00B),
				.b1(W3G01B),
				.b2(W3G02B),
				.b3(W3G10B),
				.b4(W3G11B),
				.b5(W3G12B),
				.b6(W3G20B),
				.b7(W3G21B),
				.b8(W3G22B),
				.c(c3B22G)
);

ninexnine_unit ninexnine_unit_5644(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3G00C),
				.b1(W3G01C),
				.b2(W3G02C),
				.b3(W3G10C),
				.b4(W3G11C),
				.b5(W3G12C),
				.b6(W3G20C),
				.b7(W3G21C),
				.b8(W3G22C),
				.c(c3C22G)
);

ninexnine_unit ninexnine_unit_5645(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3G00D),
				.b1(W3G01D),
				.b2(W3G02D),
				.b3(W3G10D),
				.b4(W3G11D),
				.b5(W3G12D),
				.b6(W3G20D),
				.b7(W3G21D),
				.b8(W3G22D),
				.c(c3D22G)
);

ninexnine_unit ninexnine_unit_5646(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3G00E),
				.b1(W3G01E),
				.b2(W3G02E),
				.b3(W3G10E),
				.b4(W3G11E),
				.b5(W3G12E),
				.b6(W3G20E),
				.b7(W3G21E),
				.b8(W3G22E),
				.c(c3E22G)
);

ninexnine_unit ninexnine_unit_5647(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3G00F),
				.b1(W3G01F),
				.b2(W3G02F),
				.b3(W3G10F),
				.b4(W3G11F),
				.b5(W3G12F),
				.b6(W3G20F),
				.b7(W3G21F),
				.b8(W3G22F),
				.c(c3F22G)
);

assign C322G=c3022G+c3122G+c3222G+c3322G+c3422G+c3522G+c3622G+c3722G+c3822G+c3922G+c3A22G+c3B22G+c3C22G+c3D22G+c3E22G+c3F22G;
assign A322G=(C322G>=0)?1:0;

assign P422G=A322G;

ninexnine_unit ninexnine_unit_5648(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3000H)
);

ninexnine_unit ninexnine_unit_5649(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3100H)
);

ninexnine_unit ninexnine_unit_5650(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3200H)
);

ninexnine_unit ninexnine_unit_5651(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3300H)
);

ninexnine_unit ninexnine_unit_5652(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3400H)
);

ninexnine_unit ninexnine_unit_5653(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3500H)
);

ninexnine_unit ninexnine_unit_5654(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3600H)
);

ninexnine_unit ninexnine_unit_5655(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3700H)
);

ninexnine_unit ninexnine_unit_5656(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3800H)
);

ninexnine_unit ninexnine_unit_5657(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3900H)
);

ninexnine_unit ninexnine_unit_5658(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A00H)
);

ninexnine_unit ninexnine_unit_5659(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B00H)
);

ninexnine_unit ninexnine_unit_5660(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C00H)
);

ninexnine_unit ninexnine_unit_5661(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D00H)
);

ninexnine_unit ninexnine_unit_5662(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E00H)
);

ninexnine_unit ninexnine_unit_5663(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F00H)
);

assign C300H=c3000H+c3100H+c3200H+c3300H+c3400H+c3500H+c3600H+c3700H+c3800H+c3900H+c3A00H+c3B00H+c3C00H+c3D00H+c3E00H+c3F00H;
assign A300H=(C300H>=0)?1:0;

assign P400H=A300H;

ninexnine_unit ninexnine_unit_5664(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3001H)
);

ninexnine_unit ninexnine_unit_5665(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3101H)
);

ninexnine_unit ninexnine_unit_5666(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3201H)
);

ninexnine_unit ninexnine_unit_5667(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3301H)
);

ninexnine_unit ninexnine_unit_5668(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3401H)
);

ninexnine_unit ninexnine_unit_5669(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3501H)
);

ninexnine_unit ninexnine_unit_5670(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3601H)
);

ninexnine_unit ninexnine_unit_5671(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3701H)
);

ninexnine_unit ninexnine_unit_5672(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3801H)
);

ninexnine_unit ninexnine_unit_5673(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3901H)
);

ninexnine_unit ninexnine_unit_5674(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A01H)
);

ninexnine_unit ninexnine_unit_5675(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B01H)
);

ninexnine_unit ninexnine_unit_5676(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C01H)
);

ninexnine_unit ninexnine_unit_5677(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D01H)
);

ninexnine_unit ninexnine_unit_5678(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E01H)
);

ninexnine_unit ninexnine_unit_5679(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F01H)
);

assign C301H=c3001H+c3101H+c3201H+c3301H+c3401H+c3501H+c3601H+c3701H+c3801H+c3901H+c3A01H+c3B01H+c3C01H+c3D01H+c3E01H+c3F01H;
assign A301H=(C301H>=0)?1:0;

assign P401H=A301H;

ninexnine_unit ninexnine_unit_5680(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3002H)
);

ninexnine_unit ninexnine_unit_5681(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3102H)
);

ninexnine_unit ninexnine_unit_5682(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3202H)
);

ninexnine_unit ninexnine_unit_5683(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3302H)
);

ninexnine_unit ninexnine_unit_5684(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3402H)
);

ninexnine_unit ninexnine_unit_5685(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3502H)
);

ninexnine_unit ninexnine_unit_5686(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3602H)
);

ninexnine_unit ninexnine_unit_5687(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3702H)
);

ninexnine_unit ninexnine_unit_5688(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3802H)
);

ninexnine_unit ninexnine_unit_5689(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3902H)
);

ninexnine_unit ninexnine_unit_5690(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A02H)
);

ninexnine_unit ninexnine_unit_5691(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B02H)
);

ninexnine_unit ninexnine_unit_5692(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C02H)
);

ninexnine_unit ninexnine_unit_5693(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D02H)
);

ninexnine_unit ninexnine_unit_5694(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E02H)
);

ninexnine_unit ninexnine_unit_5695(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F02H)
);

assign C302H=c3002H+c3102H+c3202H+c3302H+c3402H+c3502H+c3602H+c3702H+c3802H+c3902H+c3A02H+c3B02H+c3C02H+c3D02H+c3E02H+c3F02H;
assign A302H=(C302H>=0)?1:0;

assign P402H=A302H;

ninexnine_unit ninexnine_unit_5696(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3010H)
);

ninexnine_unit ninexnine_unit_5697(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3110H)
);

ninexnine_unit ninexnine_unit_5698(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3210H)
);

ninexnine_unit ninexnine_unit_5699(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3310H)
);

ninexnine_unit ninexnine_unit_5700(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3410H)
);

ninexnine_unit ninexnine_unit_5701(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3510H)
);

ninexnine_unit ninexnine_unit_5702(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3610H)
);

ninexnine_unit ninexnine_unit_5703(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3710H)
);

ninexnine_unit ninexnine_unit_5704(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3810H)
);

ninexnine_unit ninexnine_unit_5705(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3910H)
);

ninexnine_unit ninexnine_unit_5706(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A10H)
);

ninexnine_unit ninexnine_unit_5707(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B10H)
);

ninexnine_unit ninexnine_unit_5708(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C10H)
);

ninexnine_unit ninexnine_unit_5709(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D10H)
);

ninexnine_unit ninexnine_unit_5710(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E10H)
);

ninexnine_unit ninexnine_unit_5711(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F10H)
);

assign C310H=c3010H+c3110H+c3210H+c3310H+c3410H+c3510H+c3610H+c3710H+c3810H+c3910H+c3A10H+c3B10H+c3C10H+c3D10H+c3E10H+c3F10H;
assign A310H=(C310H>=0)?1:0;

assign P410H=A310H;

ninexnine_unit ninexnine_unit_5712(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3011H)
);

ninexnine_unit ninexnine_unit_5713(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3111H)
);

ninexnine_unit ninexnine_unit_5714(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3211H)
);

ninexnine_unit ninexnine_unit_5715(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3311H)
);

ninexnine_unit ninexnine_unit_5716(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3411H)
);

ninexnine_unit ninexnine_unit_5717(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3511H)
);

ninexnine_unit ninexnine_unit_5718(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3611H)
);

ninexnine_unit ninexnine_unit_5719(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3711H)
);

ninexnine_unit ninexnine_unit_5720(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3811H)
);

ninexnine_unit ninexnine_unit_5721(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3911H)
);

ninexnine_unit ninexnine_unit_5722(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A11H)
);

ninexnine_unit ninexnine_unit_5723(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B11H)
);

ninexnine_unit ninexnine_unit_5724(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C11H)
);

ninexnine_unit ninexnine_unit_5725(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D11H)
);

ninexnine_unit ninexnine_unit_5726(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E11H)
);

ninexnine_unit ninexnine_unit_5727(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F11H)
);

assign C311H=c3011H+c3111H+c3211H+c3311H+c3411H+c3511H+c3611H+c3711H+c3811H+c3911H+c3A11H+c3B11H+c3C11H+c3D11H+c3E11H+c3F11H;
assign A311H=(C311H>=0)?1:0;

assign P411H=A311H;

ninexnine_unit ninexnine_unit_5728(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3012H)
);

ninexnine_unit ninexnine_unit_5729(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3112H)
);

ninexnine_unit ninexnine_unit_5730(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3212H)
);

ninexnine_unit ninexnine_unit_5731(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3312H)
);

ninexnine_unit ninexnine_unit_5732(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3412H)
);

ninexnine_unit ninexnine_unit_5733(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3512H)
);

ninexnine_unit ninexnine_unit_5734(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3612H)
);

ninexnine_unit ninexnine_unit_5735(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3712H)
);

ninexnine_unit ninexnine_unit_5736(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3812H)
);

ninexnine_unit ninexnine_unit_5737(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3912H)
);

ninexnine_unit ninexnine_unit_5738(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A12H)
);

ninexnine_unit ninexnine_unit_5739(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B12H)
);

ninexnine_unit ninexnine_unit_5740(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C12H)
);

ninexnine_unit ninexnine_unit_5741(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D12H)
);

ninexnine_unit ninexnine_unit_5742(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E12H)
);

ninexnine_unit ninexnine_unit_5743(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F12H)
);

assign C312H=c3012H+c3112H+c3212H+c3312H+c3412H+c3512H+c3612H+c3712H+c3812H+c3912H+c3A12H+c3B12H+c3C12H+c3D12H+c3E12H+c3F12H;
assign A312H=(C312H>=0)?1:0;

assign P412H=A312H;

ninexnine_unit ninexnine_unit_5744(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3020H)
);

ninexnine_unit ninexnine_unit_5745(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3120H)
);

ninexnine_unit ninexnine_unit_5746(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3220H)
);

ninexnine_unit ninexnine_unit_5747(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3320H)
);

ninexnine_unit ninexnine_unit_5748(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3420H)
);

ninexnine_unit ninexnine_unit_5749(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3520H)
);

ninexnine_unit ninexnine_unit_5750(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3620H)
);

ninexnine_unit ninexnine_unit_5751(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3720H)
);

ninexnine_unit ninexnine_unit_5752(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3820H)
);

ninexnine_unit ninexnine_unit_5753(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3920H)
);

ninexnine_unit ninexnine_unit_5754(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A20H)
);

ninexnine_unit ninexnine_unit_5755(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B20H)
);

ninexnine_unit ninexnine_unit_5756(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C20H)
);

ninexnine_unit ninexnine_unit_5757(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D20H)
);

ninexnine_unit ninexnine_unit_5758(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E20H)
);

ninexnine_unit ninexnine_unit_5759(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F20H)
);

assign C320H=c3020H+c3120H+c3220H+c3320H+c3420H+c3520H+c3620H+c3720H+c3820H+c3920H+c3A20H+c3B20H+c3C20H+c3D20H+c3E20H+c3F20H;
assign A320H=(C320H>=0)?1:0;

assign P420H=A320H;

ninexnine_unit ninexnine_unit_5760(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3021H)
);

ninexnine_unit ninexnine_unit_5761(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3121H)
);

ninexnine_unit ninexnine_unit_5762(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3221H)
);

ninexnine_unit ninexnine_unit_5763(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3321H)
);

ninexnine_unit ninexnine_unit_5764(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3421H)
);

ninexnine_unit ninexnine_unit_5765(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3521H)
);

ninexnine_unit ninexnine_unit_5766(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3621H)
);

ninexnine_unit ninexnine_unit_5767(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3721H)
);

ninexnine_unit ninexnine_unit_5768(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3821H)
);

ninexnine_unit ninexnine_unit_5769(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3921H)
);

ninexnine_unit ninexnine_unit_5770(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A21H)
);

ninexnine_unit ninexnine_unit_5771(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B21H)
);

ninexnine_unit ninexnine_unit_5772(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C21H)
);

ninexnine_unit ninexnine_unit_5773(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D21H)
);

ninexnine_unit ninexnine_unit_5774(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E21H)
);

ninexnine_unit ninexnine_unit_5775(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F21H)
);

assign C321H=c3021H+c3121H+c3221H+c3321H+c3421H+c3521H+c3621H+c3721H+c3821H+c3921H+c3A21H+c3B21H+c3C21H+c3D21H+c3E21H+c3F21H;
assign A321H=(C321H>=0)?1:0;

assign P421H=A321H;

ninexnine_unit ninexnine_unit_5776(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3H000),
				.b1(W3H010),
				.b2(W3H020),
				.b3(W3H100),
				.b4(W3H110),
				.b5(W3H120),
				.b6(W3H200),
				.b7(W3H210),
				.b8(W3H220),
				.c(c3022H)
);

ninexnine_unit ninexnine_unit_5777(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3H001),
				.b1(W3H011),
				.b2(W3H021),
				.b3(W3H101),
				.b4(W3H111),
				.b5(W3H121),
				.b6(W3H201),
				.b7(W3H211),
				.b8(W3H221),
				.c(c3122H)
);

ninexnine_unit ninexnine_unit_5778(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3H002),
				.b1(W3H012),
				.b2(W3H022),
				.b3(W3H102),
				.b4(W3H112),
				.b5(W3H122),
				.b6(W3H202),
				.b7(W3H212),
				.b8(W3H222),
				.c(c3222H)
);

ninexnine_unit ninexnine_unit_5779(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3H003),
				.b1(W3H013),
				.b2(W3H023),
				.b3(W3H103),
				.b4(W3H113),
				.b5(W3H123),
				.b6(W3H203),
				.b7(W3H213),
				.b8(W3H223),
				.c(c3322H)
);

ninexnine_unit ninexnine_unit_5780(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3H004),
				.b1(W3H014),
				.b2(W3H024),
				.b3(W3H104),
				.b4(W3H114),
				.b5(W3H124),
				.b6(W3H204),
				.b7(W3H214),
				.b8(W3H224),
				.c(c3422H)
);

ninexnine_unit ninexnine_unit_5781(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3H005),
				.b1(W3H015),
				.b2(W3H025),
				.b3(W3H105),
				.b4(W3H115),
				.b5(W3H125),
				.b6(W3H205),
				.b7(W3H215),
				.b8(W3H225),
				.c(c3522H)
);

ninexnine_unit ninexnine_unit_5782(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3H006),
				.b1(W3H016),
				.b2(W3H026),
				.b3(W3H106),
				.b4(W3H116),
				.b5(W3H126),
				.b6(W3H206),
				.b7(W3H216),
				.b8(W3H226),
				.c(c3622H)
);

ninexnine_unit ninexnine_unit_5783(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3H007),
				.b1(W3H017),
				.b2(W3H027),
				.b3(W3H107),
				.b4(W3H117),
				.b5(W3H127),
				.b6(W3H207),
				.b7(W3H217),
				.b8(W3H227),
				.c(c3722H)
);

ninexnine_unit ninexnine_unit_5784(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3H008),
				.b1(W3H018),
				.b2(W3H028),
				.b3(W3H108),
				.b4(W3H118),
				.b5(W3H128),
				.b6(W3H208),
				.b7(W3H218),
				.b8(W3H228),
				.c(c3822H)
);

ninexnine_unit ninexnine_unit_5785(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3H009),
				.b1(W3H019),
				.b2(W3H029),
				.b3(W3H109),
				.b4(W3H119),
				.b5(W3H129),
				.b6(W3H209),
				.b7(W3H219),
				.b8(W3H229),
				.c(c3922H)
);

ninexnine_unit ninexnine_unit_5786(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3H00A),
				.b1(W3H01A),
				.b2(W3H02A),
				.b3(W3H10A),
				.b4(W3H11A),
				.b5(W3H12A),
				.b6(W3H20A),
				.b7(W3H21A),
				.b8(W3H22A),
				.c(c3A22H)
);

ninexnine_unit ninexnine_unit_5787(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3H00B),
				.b1(W3H01B),
				.b2(W3H02B),
				.b3(W3H10B),
				.b4(W3H11B),
				.b5(W3H12B),
				.b6(W3H20B),
				.b7(W3H21B),
				.b8(W3H22B),
				.c(c3B22H)
);

ninexnine_unit ninexnine_unit_5788(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3H00C),
				.b1(W3H01C),
				.b2(W3H02C),
				.b3(W3H10C),
				.b4(W3H11C),
				.b5(W3H12C),
				.b6(W3H20C),
				.b7(W3H21C),
				.b8(W3H22C),
				.c(c3C22H)
);

ninexnine_unit ninexnine_unit_5789(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3H00D),
				.b1(W3H01D),
				.b2(W3H02D),
				.b3(W3H10D),
				.b4(W3H11D),
				.b5(W3H12D),
				.b6(W3H20D),
				.b7(W3H21D),
				.b8(W3H22D),
				.c(c3D22H)
);

ninexnine_unit ninexnine_unit_5790(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3H00E),
				.b1(W3H01E),
				.b2(W3H02E),
				.b3(W3H10E),
				.b4(W3H11E),
				.b5(W3H12E),
				.b6(W3H20E),
				.b7(W3H21E),
				.b8(W3H22E),
				.c(c3E22H)
);

ninexnine_unit ninexnine_unit_5791(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3H00F),
				.b1(W3H01F),
				.b2(W3H02F),
				.b3(W3H10F),
				.b4(W3H11F),
				.b5(W3H12F),
				.b6(W3H20F),
				.b7(W3H21F),
				.b8(W3H22F),
				.c(c3F22H)
);

assign C322H=c3022H+c3122H+c3222H+c3322H+c3422H+c3522H+c3622H+c3722H+c3822H+c3922H+c3A22H+c3B22H+c3C22H+c3D22H+c3E22H+c3F22H;
assign A322H=(C322H>=0)?1:0;

assign P422H=A322H;

ninexnine_unit ninexnine_unit_5792(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3000I)
);

ninexnine_unit ninexnine_unit_5793(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3100I)
);

ninexnine_unit ninexnine_unit_5794(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3200I)
);

ninexnine_unit ninexnine_unit_5795(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3300I)
);

ninexnine_unit ninexnine_unit_5796(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3400I)
);

ninexnine_unit ninexnine_unit_5797(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3500I)
);

ninexnine_unit ninexnine_unit_5798(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3600I)
);

ninexnine_unit ninexnine_unit_5799(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3700I)
);

ninexnine_unit ninexnine_unit_5800(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3800I)
);

ninexnine_unit ninexnine_unit_5801(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3900I)
);

ninexnine_unit ninexnine_unit_5802(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A00I)
);

ninexnine_unit ninexnine_unit_5803(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B00I)
);

ninexnine_unit ninexnine_unit_5804(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C00I)
);

ninexnine_unit ninexnine_unit_5805(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D00I)
);

ninexnine_unit ninexnine_unit_5806(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E00I)
);

ninexnine_unit ninexnine_unit_5807(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F00I)
);

assign C300I=c3000I+c3100I+c3200I+c3300I+c3400I+c3500I+c3600I+c3700I+c3800I+c3900I+c3A00I+c3B00I+c3C00I+c3D00I+c3E00I+c3F00I;
assign A300I=(C300I>=0)?1:0;

assign P400I=A300I;

ninexnine_unit ninexnine_unit_5808(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3001I)
);

ninexnine_unit ninexnine_unit_5809(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3101I)
);

ninexnine_unit ninexnine_unit_5810(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3201I)
);

ninexnine_unit ninexnine_unit_5811(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3301I)
);

ninexnine_unit ninexnine_unit_5812(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3401I)
);

ninexnine_unit ninexnine_unit_5813(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3501I)
);

ninexnine_unit ninexnine_unit_5814(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3601I)
);

ninexnine_unit ninexnine_unit_5815(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3701I)
);

ninexnine_unit ninexnine_unit_5816(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3801I)
);

ninexnine_unit ninexnine_unit_5817(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3901I)
);

ninexnine_unit ninexnine_unit_5818(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A01I)
);

ninexnine_unit ninexnine_unit_5819(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B01I)
);

ninexnine_unit ninexnine_unit_5820(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C01I)
);

ninexnine_unit ninexnine_unit_5821(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D01I)
);

ninexnine_unit ninexnine_unit_5822(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E01I)
);

ninexnine_unit ninexnine_unit_5823(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F01I)
);

assign C301I=c3001I+c3101I+c3201I+c3301I+c3401I+c3501I+c3601I+c3701I+c3801I+c3901I+c3A01I+c3B01I+c3C01I+c3D01I+c3E01I+c3F01I;
assign A301I=(C301I>=0)?1:0;

assign P401I=A301I;

ninexnine_unit ninexnine_unit_5824(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3002I)
);

ninexnine_unit ninexnine_unit_5825(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3102I)
);

ninexnine_unit ninexnine_unit_5826(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3202I)
);

ninexnine_unit ninexnine_unit_5827(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3302I)
);

ninexnine_unit ninexnine_unit_5828(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3402I)
);

ninexnine_unit ninexnine_unit_5829(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3502I)
);

ninexnine_unit ninexnine_unit_5830(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3602I)
);

ninexnine_unit ninexnine_unit_5831(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3702I)
);

ninexnine_unit ninexnine_unit_5832(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3802I)
);

ninexnine_unit ninexnine_unit_5833(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3902I)
);

ninexnine_unit ninexnine_unit_5834(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A02I)
);

ninexnine_unit ninexnine_unit_5835(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B02I)
);

ninexnine_unit ninexnine_unit_5836(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C02I)
);

ninexnine_unit ninexnine_unit_5837(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D02I)
);

ninexnine_unit ninexnine_unit_5838(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E02I)
);

ninexnine_unit ninexnine_unit_5839(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F02I)
);

assign C302I=c3002I+c3102I+c3202I+c3302I+c3402I+c3502I+c3602I+c3702I+c3802I+c3902I+c3A02I+c3B02I+c3C02I+c3D02I+c3E02I+c3F02I;
assign A302I=(C302I>=0)?1:0;

assign P402I=A302I;

ninexnine_unit ninexnine_unit_5840(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3010I)
);

ninexnine_unit ninexnine_unit_5841(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3110I)
);

ninexnine_unit ninexnine_unit_5842(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3210I)
);

ninexnine_unit ninexnine_unit_5843(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3310I)
);

ninexnine_unit ninexnine_unit_5844(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3410I)
);

ninexnine_unit ninexnine_unit_5845(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3510I)
);

ninexnine_unit ninexnine_unit_5846(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3610I)
);

ninexnine_unit ninexnine_unit_5847(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3710I)
);

ninexnine_unit ninexnine_unit_5848(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3810I)
);

ninexnine_unit ninexnine_unit_5849(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3910I)
);

ninexnine_unit ninexnine_unit_5850(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A10I)
);

ninexnine_unit ninexnine_unit_5851(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B10I)
);

ninexnine_unit ninexnine_unit_5852(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C10I)
);

ninexnine_unit ninexnine_unit_5853(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D10I)
);

ninexnine_unit ninexnine_unit_5854(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E10I)
);

ninexnine_unit ninexnine_unit_5855(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F10I)
);

assign C310I=c3010I+c3110I+c3210I+c3310I+c3410I+c3510I+c3610I+c3710I+c3810I+c3910I+c3A10I+c3B10I+c3C10I+c3D10I+c3E10I+c3F10I;
assign A310I=(C310I>=0)?1:0;

assign P410I=A310I;

ninexnine_unit ninexnine_unit_5856(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3011I)
);

ninexnine_unit ninexnine_unit_5857(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3111I)
);

ninexnine_unit ninexnine_unit_5858(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3211I)
);

ninexnine_unit ninexnine_unit_5859(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3311I)
);

ninexnine_unit ninexnine_unit_5860(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3411I)
);

ninexnine_unit ninexnine_unit_5861(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3511I)
);

ninexnine_unit ninexnine_unit_5862(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3611I)
);

ninexnine_unit ninexnine_unit_5863(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3711I)
);

ninexnine_unit ninexnine_unit_5864(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3811I)
);

ninexnine_unit ninexnine_unit_5865(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3911I)
);

ninexnine_unit ninexnine_unit_5866(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A11I)
);

ninexnine_unit ninexnine_unit_5867(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B11I)
);

ninexnine_unit ninexnine_unit_5868(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C11I)
);

ninexnine_unit ninexnine_unit_5869(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D11I)
);

ninexnine_unit ninexnine_unit_5870(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E11I)
);

ninexnine_unit ninexnine_unit_5871(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F11I)
);

assign C311I=c3011I+c3111I+c3211I+c3311I+c3411I+c3511I+c3611I+c3711I+c3811I+c3911I+c3A11I+c3B11I+c3C11I+c3D11I+c3E11I+c3F11I;
assign A311I=(C311I>=0)?1:0;

assign P411I=A311I;

ninexnine_unit ninexnine_unit_5872(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3012I)
);

ninexnine_unit ninexnine_unit_5873(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3112I)
);

ninexnine_unit ninexnine_unit_5874(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3212I)
);

ninexnine_unit ninexnine_unit_5875(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3312I)
);

ninexnine_unit ninexnine_unit_5876(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3412I)
);

ninexnine_unit ninexnine_unit_5877(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3512I)
);

ninexnine_unit ninexnine_unit_5878(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3612I)
);

ninexnine_unit ninexnine_unit_5879(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3712I)
);

ninexnine_unit ninexnine_unit_5880(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3812I)
);

ninexnine_unit ninexnine_unit_5881(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3912I)
);

ninexnine_unit ninexnine_unit_5882(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A12I)
);

ninexnine_unit ninexnine_unit_5883(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B12I)
);

ninexnine_unit ninexnine_unit_5884(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C12I)
);

ninexnine_unit ninexnine_unit_5885(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D12I)
);

ninexnine_unit ninexnine_unit_5886(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E12I)
);

ninexnine_unit ninexnine_unit_5887(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F12I)
);

assign C312I=c3012I+c3112I+c3212I+c3312I+c3412I+c3512I+c3612I+c3712I+c3812I+c3912I+c3A12I+c3B12I+c3C12I+c3D12I+c3E12I+c3F12I;
assign A312I=(C312I>=0)?1:0;

assign P412I=A312I;

ninexnine_unit ninexnine_unit_5888(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3020I)
);

ninexnine_unit ninexnine_unit_5889(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3120I)
);

ninexnine_unit ninexnine_unit_5890(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3220I)
);

ninexnine_unit ninexnine_unit_5891(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3320I)
);

ninexnine_unit ninexnine_unit_5892(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3420I)
);

ninexnine_unit ninexnine_unit_5893(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3520I)
);

ninexnine_unit ninexnine_unit_5894(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3620I)
);

ninexnine_unit ninexnine_unit_5895(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3720I)
);

ninexnine_unit ninexnine_unit_5896(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3820I)
);

ninexnine_unit ninexnine_unit_5897(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3920I)
);

ninexnine_unit ninexnine_unit_5898(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A20I)
);

ninexnine_unit ninexnine_unit_5899(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B20I)
);

ninexnine_unit ninexnine_unit_5900(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C20I)
);

ninexnine_unit ninexnine_unit_5901(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D20I)
);

ninexnine_unit ninexnine_unit_5902(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E20I)
);

ninexnine_unit ninexnine_unit_5903(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F20I)
);

assign C320I=c3020I+c3120I+c3220I+c3320I+c3420I+c3520I+c3620I+c3720I+c3820I+c3920I+c3A20I+c3B20I+c3C20I+c3D20I+c3E20I+c3F20I;
assign A320I=(C320I>=0)?1:0;

assign P420I=A320I;

ninexnine_unit ninexnine_unit_5904(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3021I)
);

ninexnine_unit ninexnine_unit_5905(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3121I)
);

ninexnine_unit ninexnine_unit_5906(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3221I)
);

ninexnine_unit ninexnine_unit_5907(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3321I)
);

ninexnine_unit ninexnine_unit_5908(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3421I)
);

ninexnine_unit ninexnine_unit_5909(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3521I)
);

ninexnine_unit ninexnine_unit_5910(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3621I)
);

ninexnine_unit ninexnine_unit_5911(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3721I)
);

ninexnine_unit ninexnine_unit_5912(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3821I)
);

ninexnine_unit ninexnine_unit_5913(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3921I)
);

ninexnine_unit ninexnine_unit_5914(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A21I)
);

ninexnine_unit ninexnine_unit_5915(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B21I)
);

ninexnine_unit ninexnine_unit_5916(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C21I)
);

ninexnine_unit ninexnine_unit_5917(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D21I)
);

ninexnine_unit ninexnine_unit_5918(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E21I)
);

ninexnine_unit ninexnine_unit_5919(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F21I)
);

assign C321I=c3021I+c3121I+c3221I+c3321I+c3421I+c3521I+c3621I+c3721I+c3821I+c3921I+c3A21I+c3B21I+c3C21I+c3D21I+c3E21I+c3F21I;
assign A321I=(C321I>=0)?1:0;

assign P421I=A321I;

ninexnine_unit ninexnine_unit_5920(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3I000),
				.b1(W3I010),
				.b2(W3I020),
				.b3(W3I100),
				.b4(W3I110),
				.b5(W3I120),
				.b6(W3I200),
				.b7(W3I210),
				.b8(W3I220),
				.c(c3022I)
);

ninexnine_unit ninexnine_unit_5921(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3I001),
				.b1(W3I011),
				.b2(W3I021),
				.b3(W3I101),
				.b4(W3I111),
				.b5(W3I121),
				.b6(W3I201),
				.b7(W3I211),
				.b8(W3I221),
				.c(c3122I)
);

ninexnine_unit ninexnine_unit_5922(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3I002),
				.b1(W3I012),
				.b2(W3I022),
				.b3(W3I102),
				.b4(W3I112),
				.b5(W3I122),
				.b6(W3I202),
				.b7(W3I212),
				.b8(W3I222),
				.c(c3222I)
);

ninexnine_unit ninexnine_unit_5923(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3I003),
				.b1(W3I013),
				.b2(W3I023),
				.b3(W3I103),
				.b4(W3I113),
				.b5(W3I123),
				.b6(W3I203),
				.b7(W3I213),
				.b8(W3I223),
				.c(c3322I)
);

ninexnine_unit ninexnine_unit_5924(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3I004),
				.b1(W3I014),
				.b2(W3I024),
				.b3(W3I104),
				.b4(W3I114),
				.b5(W3I124),
				.b6(W3I204),
				.b7(W3I214),
				.b8(W3I224),
				.c(c3422I)
);

ninexnine_unit ninexnine_unit_5925(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3I005),
				.b1(W3I015),
				.b2(W3I025),
				.b3(W3I105),
				.b4(W3I115),
				.b5(W3I125),
				.b6(W3I205),
				.b7(W3I215),
				.b8(W3I225),
				.c(c3522I)
);

ninexnine_unit ninexnine_unit_5926(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3I006),
				.b1(W3I016),
				.b2(W3I026),
				.b3(W3I106),
				.b4(W3I116),
				.b5(W3I126),
				.b6(W3I206),
				.b7(W3I216),
				.b8(W3I226),
				.c(c3622I)
);

ninexnine_unit ninexnine_unit_5927(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3I007),
				.b1(W3I017),
				.b2(W3I027),
				.b3(W3I107),
				.b4(W3I117),
				.b5(W3I127),
				.b6(W3I207),
				.b7(W3I217),
				.b8(W3I227),
				.c(c3722I)
);

ninexnine_unit ninexnine_unit_5928(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3I008),
				.b1(W3I018),
				.b2(W3I028),
				.b3(W3I108),
				.b4(W3I118),
				.b5(W3I128),
				.b6(W3I208),
				.b7(W3I218),
				.b8(W3I228),
				.c(c3822I)
);

ninexnine_unit ninexnine_unit_5929(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3I009),
				.b1(W3I019),
				.b2(W3I029),
				.b3(W3I109),
				.b4(W3I119),
				.b5(W3I129),
				.b6(W3I209),
				.b7(W3I219),
				.b8(W3I229),
				.c(c3922I)
);

ninexnine_unit ninexnine_unit_5930(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3I00A),
				.b1(W3I01A),
				.b2(W3I02A),
				.b3(W3I10A),
				.b4(W3I11A),
				.b5(W3I12A),
				.b6(W3I20A),
				.b7(W3I21A),
				.b8(W3I22A),
				.c(c3A22I)
);

ninexnine_unit ninexnine_unit_5931(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3I00B),
				.b1(W3I01B),
				.b2(W3I02B),
				.b3(W3I10B),
				.b4(W3I11B),
				.b5(W3I12B),
				.b6(W3I20B),
				.b7(W3I21B),
				.b8(W3I22B),
				.c(c3B22I)
);

ninexnine_unit ninexnine_unit_5932(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3I00C),
				.b1(W3I01C),
				.b2(W3I02C),
				.b3(W3I10C),
				.b4(W3I11C),
				.b5(W3I12C),
				.b6(W3I20C),
				.b7(W3I21C),
				.b8(W3I22C),
				.c(c3C22I)
);

ninexnine_unit ninexnine_unit_5933(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3I00D),
				.b1(W3I01D),
				.b2(W3I02D),
				.b3(W3I10D),
				.b4(W3I11D),
				.b5(W3I12D),
				.b6(W3I20D),
				.b7(W3I21D),
				.b8(W3I22D),
				.c(c3D22I)
);

ninexnine_unit ninexnine_unit_5934(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3I00E),
				.b1(W3I01E),
				.b2(W3I02E),
				.b3(W3I10E),
				.b4(W3I11E),
				.b5(W3I12E),
				.b6(W3I20E),
				.b7(W3I21E),
				.b8(W3I22E),
				.c(c3E22I)
);

ninexnine_unit ninexnine_unit_5935(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3I00F),
				.b1(W3I01F),
				.b2(W3I02F),
				.b3(W3I10F),
				.b4(W3I11F),
				.b5(W3I12F),
				.b6(W3I20F),
				.b7(W3I21F),
				.b8(W3I22F),
				.c(c3F22I)
);

assign C322I=c3022I+c3122I+c3222I+c3322I+c3422I+c3522I+c3622I+c3722I+c3822I+c3922I+c3A22I+c3B22I+c3C22I+c3D22I+c3E22I+c3F22I;
assign A322I=(C322I>=0)?1:0;

assign P422I=A322I;

ninexnine_unit ninexnine_unit_5936(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3000J)
);

ninexnine_unit ninexnine_unit_5937(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3100J)
);

ninexnine_unit ninexnine_unit_5938(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3200J)
);

ninexnine_unit ninexnine_unit_5939(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3300J)
);

ninexnine_unit ninexnine_unit_5940(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3400J)
);

ninexnine_unit ninexnine_unit_5941(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3500J)
);

ninexnine_unit ninexnine_unit_5942(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3600J)
);

ninexnine_unit ninexnine_unit_5943(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3700J)
);

ninexnine_unit ninexnine_unit_5944(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3800J)
);

ninexnine_unit ninexnine_unit_5945(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3900J)
);

ninexnine_unit ninexnine_unit_5946(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A00J)
);

ninexnine_unit ninexnine_unit_5947(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B00J)
);

ninexnine_unit ninexnine_unit_5948(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C00J)
);

ninexnine_unit ninexnine_unit_5949(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D00J)
);

ninexnine_unit ninexnine_unit_5950(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E00J)
);

ninexnine_unit ninexnine_unit_5951(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F00J)
);

assign C300J=c3000J+c3100J+c3200J+c3300J+c3400J+c3500J+c3600J+c3700J+c3800J+c3900J+c3A00J+c3B00J+c3C00J+c3D00J+c3E00J+c3F00J;
assign A300J=(C300J>=0)?1:0;

assign P400J=A300J;

ninexnine_unit ninexnine_unit_5952(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3001J)
);

ninexnine_unit ninexnine_unit_5953(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3101J)
);

ninexnine_unit ninexnine_unit_5954(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3201J)
);

ninexnine_unit ninexnine_unit_5955(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3301J)
);

ninexnine_unit ninexnine_unit_5956(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3401J)
);

ninexnine_unit ninexnine_unit_5957(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3501J)
);

ninexnine_unit ninexnine_unit_5958(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3601J)
);

ninexnine_unit ninexnine_unit_5959(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3701J)
);

ninexnine_unit ninexnine_unit_5960(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3801J)
);

ninexnine_unit ninexnine_unit_5961(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3901J)
);

ninexnine_unit ninexnine_unit_5962(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A01J)
);

ninexnine_unit ninexnine_unit_5963(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B01J)
);

ninexnine_unit ninexnine_unit_5964(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C01J)
);

ninexnine_unit ninexnine_unit_5965(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D01J)
);

ninexnine_unit ninexnine_unit_5966(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E01J)
);

ninexnine_unit ninexnine_unit_5967(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F01J)
);

assign C301J=c3001J+c3101J+c3201J+c3301J+c3401J+c3501J+c3601J+c3701J+c3801J+c3901J+c3A01J+c3B01J+c3C01J+c3D01J+c3E01J+c3F01J;
assign A301J=(C301J>=0)?1:0;

assign P401J=A301J;

ninexnine_unit ninexnine_unit_5968(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3002J)
);

ninexnine_unit ninexnine_unit_5969(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3102J)
);

ninexnine_unit ninexnine_unit_5970(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3202J)
);

ninexnine_unit ninexnine_unit_5971(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3302J)
);

ninexnine_unit ninexnine_unit_5972(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3402J)
);

ninexnine_unit ninexnine_unit_5973(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3502J)
);

ninexnine_unit ninexnine_unit_5974(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3602J)
);

ninexnine_unit ninexnine_unit_5975(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3702J)
);

ninexnine_unit ninexnine_unit_5976(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3802J)
);

ninexnine_unit ninexnine_unit_5977(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3902J)
);

ninexnine_unit ninexnine_unit_5978(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A02J)
);

ninexnine_unit ninexnine_unit_5979(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B02J)
);

ninexnine_unit ninexnine_unit_5980(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C02J)
);

ninexnine_unit ninexnine_unit_5981(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D02J)
);

ninexnine_unit ninexnine_unit_5982(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E02J)
);

ninexnine_unit ninexnine_unit_5983(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F02J)
);

assign C302J=c3002J+c3102J+c3202J+c3302J+c3402J+c3502J+c3602J+c3702J+c3802J+c3902J+c3A02J+c3B02J+c3C02J+c3D02J+c3E02J+c3F02J;
assign A302J=(C302J>=0)?1:0;

assign P402J=A302J;

ninexnine_unit ninexnine_unit_5984(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3010J)
);

ninexnine_unit ninexnine_unit_5985(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3110J)
);

ninexnine_unit ninexnine_unit_5986(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3210J)
);

ninexnine_unit ninexnine_unit_5987(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3310J)
);

ninexnine_unit ninexnine_unit_5988(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3410J)
);

ninexnine_unit ninexnine_unit_5989(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3510J)
);

ninexnine_unit ninexnine_unit_5990(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3610J)
);

ninexnine_unit ninexnine_unit_5991(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3710J)
);

ninexnine_unit ninexnine_unit_5992(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3810J)
);

ninexnine_unit ninexnine_unit_5993(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3910J)
);

ninexnine_unit ninexnine_unit_5994(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A10J)
);

ninexnine_unit ninexnine_unit_5995(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B10J)
);

ninexnine_unit ninexnine_unit_5996(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C10J)
);

ninexnine_unit ninexnine_unit_5997(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D10J)
);

ninexnine_unit ninexnine_unit_5998(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E10J)
);

ninexnine_unit ninexnine_unit_5999(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F10J)
);

assign C310J=c3010J+c3110J+c3210J+c3310J+c3410J+c3510J+c3610J+c3710J+c3810J+c3910J+c3A10J+c3B10J+c3C10J+c3D10J+c3E10J+c3F10J;
assign A310J=(C310J>=0)?1:0;

assign P410J=A310J;

ninexnine_unit ninexnine_unit_6000(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3011J)
);

ninexnine_unit ninexnine_unit_6001(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3111J)
);

ninexnine_unit ninexnine_unit_6002(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3211J)
);

ninexnine_unit ninexnine_unit_6003(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3311J)
);

ninexnine_unit ninexnine_unit_6004(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3411J)
);

ninexnine_unit ninexnine_unit_6005(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3511J)
);

ninexnine_unit ninexnine_unit_6006(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3611J)
);

ninexnine_unit ninexnine_unit_6007(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3711J)
);

ninexnine_unit ninexnine_unit_6008(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3811J)
);

ninexnine_unit ninexnine_unit_6009(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3911J)
);

ninexnine_unit ninexnine_unit_6010(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A11J)
);

ninexnine_unit ninexnine_unit_6011(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B11J)
);

ninexnine_unit ninexnine_unit_6012(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C11J)
);

ninexnine_unit ninexnine_unit_6013(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D11J)
);

ninexnine_unit ninexnine_unit_6014(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E11J)
);

ninexnine_unit ninexnine_unit_6015(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F11J)
);

assign C311J=c3011J+c3111J+c3211J+c3311J+c3411J+c3511J+c3611J+c3711J+c3811J+c3911J+c3A11J+c3B11J+c3C11J+c3D11J+c3E11J+c3F11J;
assign A311J=(C311J>=0)?1:0;

assign P411J=A311J;

ninexnine_unit ninexnine_unit_6016(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3012J)
);

ninexnine_unit ninexnine_unit_6017(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3112J)
);

ninexnine_unit ninexnine_unit_6018(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3212J)
);

ninexnine_unit ninexnine_unit_6019(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3312J)
);

ninexnine_unit ninexnine_unit_6020(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3412J)
);

ninexnine_unit ninexnine_unit_6021(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3512J)
);

ninexnine_unit ninexnine_unit_6022(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3612J)
);

ninexnine_unit ninexnine_unit_6023(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3712J)
);

ninexnine_unit ninexnine_unit_6024(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3812J)
);

ninexnine_unit ninexnine_unit_6025(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3912J)
);

ninexnine_unit ninexnine_unit_6026(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A12J)
);

ninexnine_unit ninexnine_unit_6027(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B12J)
);

ninexnine_unit ninexnine_unit_6028(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C12J)
);

ninexnine_unit ninexnine_unit_6029(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D12J)
);

ninexnine_unit ninexnine_unit_6030(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E12J)
);

ninexnine_unit ninexnine_unit_6031(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F12J)
);

assign C312J=c3012J+c3112J+c3212J+c3312J+c3412J+c3512J+c3612J+c3712J+c3812J+c3912J+c3A12J+c3B12J+c3C12J+c3D12J+c3E12J+c3F12J;
assign A312J=(C312J>=0)?1:0;

assign P412J=A312J;

ninexnine_unit ninexnine_unit_6032(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3020J)
);

ninexnine_unit ninexnine_unit_6033(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3120J)
);

ninexnine_unit ninexnine_unit_6034(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3220J)
);

ninexnine_unit ninexnine_unit_6035(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3320J)
);

ninexnine_unit ninexnine_unit_6036(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3420J)
);

ninexnine_unit ninexnine_unit_6037(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3520J)
);

ninexnine_unit ninexnine_unit_6038(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3620J)
);

ninexnine_unit ninexnine_unit_6039(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3720J)
);

ninexnine_unit ninexnine_unit_6040(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3820J)
);

ninexnine_unit ninexnine_unit_6041(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3920J)
);

ninexnine_unit ninexnine_unit_6042(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A20J)
);

ninexnine_unit ninexnine_unit_6043(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B20J)
);

ninexnine_unit ninexnine_unit_6044(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C20J)
);

ninexnine_unit ninexnine_unit_6045(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D20J)
);

ninexnine_unit ninexnine_unit_6046(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E20J)
);

ninexnine_unit ninexnine_unit_6047(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F20J)
);

assign C320J=c3020J+c3120J+c3220J+c3320J+c3420J+c3520J+c3620J+c3720J+c3820J+c3920J+c3A20J+c3B20J+c3C20J+c3D20J+c3E20J+c3F20J;
assign A320J=(C320J>=0)?1:0;

assign P420J=A320J;

ninexnine_unit ninexnine_unit_6048(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3021J)
);

ninexnine_unit ninexnine_unit_6049(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3121J)
);

ninexnine_unit ninexnine_unit_6050(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3221J)
);

ninexnine_unit ninexnine_unit_6051(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3321J)
);

ninexnine_unit ninexnine_unit_6052(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3421J)
);

ninexnine_unit ninexnine_unit_6053(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3521J)
);

ninexnine_unit ninexnine_unit_6054(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3621J)
);

ninexnine_unit ninexnine_unit_6055(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3721J)
);

ninexnine_unit ninexnine_unit_6056(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3821J)
);

ninexnine_unit ninexnine_unit_6057(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3921J)
);

ninexnine_unit ninexnine_unit_6058(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A21J)
);

ninexnine_unit ninexnine_unit_6059(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B21J)
);

ninexnine_unit ninexnine_unit_6060(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C21J)
);

ninexnine_unit ninexnine_unit_6061(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D21J)
);

ninexnine_unit ninexnine_unit_6062(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E21J)
);

ninexnine_unit ninexnine_unit_6063(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F21J)
);

assign C321J=c3021J+c3121J+c3221J+c3321J+c3421J+c3521J+c3621J+c3721J+c3821J+c3921J+c3A21J+c3B21J+c3C21J+c3D21J+c3E21J+c3F21J;
assign A321J=(C321J>=0)?1:0;

assign P421J=A321J;

ninexnine_unit ninexnine_unit_6064(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3J000),
				.b1(W3J010),
				.b2(W3J020),
				.b3(W3J100),
				.b4(W3J110),
				.b5(W3J120),
				.b6(W3J200),
				.b7(W3J210),
				.b8(W3J220),
				.c(c3022J)
);

ninexnine_unit ninexnine_unit_6065(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3J001),
				.b1(W3J011),
				.b2(W3J021),
				.b3(W3J101),
				.b4(W3J111),
				.b5(W3J121),
				.b6(W3J201),
				.b7(W3J211),
				.b8(W3J221),
				.c(c3122J)
);

ninexnine_unit ninexnine_unit_6066(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3J002),
				.b1(W3J012),
				.b2(W3J022),
				.b3(W3J102),
				.b4(W3J112),
				.b5(W3J122),
				.b6(W3J202),
				.b7(W3J212),
				.b8(W3J222),
				.c(c3222J)
);

ninexnine_unit ninexnine_unit_6067(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3J003),
				.b1(W3J013),
				.b2(W3J023),
				.b3(W3J103),
				.b4(W3J113),
				.b5(W3J123),
				.b6(W3J203),
				.b7(W3J213),
				.b8(W3J223),
				.c(c3322J)
);

ninexnine_unit ninexnine_unit_6068(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3J004),
				.b1(W3J014),
				.b2(W3J024),
				.b3(W3J104),
				.b4(W3J114),
				.b5(W3J124),
				.b6(W3J204),
				.b7(W3J214),
				.b8(W3J224),
				.c(c3422J)
);

ninexnine_unit ninexnine_unit_6069(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3J005),
				.b1(W3J015),
				.b2(W3J025),
				.b3(W3J105),
				.b4(W3J115),
				.b5(W3J125),
				.b6(W3J205),
				.b7(W3J215),
				.b8(W3J225),
				.c(c3522J)
);

ninexnine_unit ninexnine_unit_6070(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3J006),
				.b1(W3J016),
				.b2(W3J026),
				.b3(W3J106),
				.b4(W3J116),
				.b5(W3J126),
				.b6(W3J206),
				.b7(W3J216),
				.b8(W3J226),
				.c(c3622J)
);

ninexnine_unit ninexnine_unit_6071(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3J007),
				.b1(W3J017),
				.b2(W3J027),
				.b3(W3J107),
				.b4(W3J117),
				.b5(W3J127),
				.b6(W3J207),
				.b7(W3J217),
				.b8(W3J227),
				.c(c3722J)
);

ninexnine_unit ninexnine_unit_6072(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3J008),
				.b1(W3J018),
				.b2(W3J028),
				.b3(W3J108),
				.b4(W3J118),
				.b5(W3J128),
				.b6(W3J208),
				.b7(W3J218),
				.b8(W3J228),
				.c(c3822J)
);

ninexnine_unit ninexnine_unit_6073(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3J009),
				.b1(W3J019),
				.b2(W3J029),
				.b3(W3J109),
				.b4(W3J119),
				.b5(W3J129),
				.b6(W3J209),
				.b7(W3J219),
				.b8(W3J229),
				.c(c3922J)
);

ninexnine_unit ninexnine_unit_6074(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3J00A),
				.b1(W3J01A),
				.b2(W3J02A),
				.b3(W3J10A),
				.b4(W3J11A),
				.b5(W3J12A),
				.b6(W3J20A),
				.b7(W3J21A),
				.b8(W3J22A),
				.c(c3A22J)
);

ninexnine_unit ninexnine_unit_6075(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3J00B),
				.b1(W3J01B),
				.b2(W3J02B),
				.b3(W3J10B),
				.b4(W3J11B),
				.b5(W3J12B),
				.b6(W3J20B),
				.b7(W3J21B),
				.b8(W3J22B),
				.c(c3B22J)
);

ninexnine_unit ninexnine_unit_6076(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3J00C),
				.b1(W3J01C),
				.b2(W3J02C),
				.b3(W3J10C),
				.b4(W3J11C),
				.b5(W3J12C),
				.b6(W3J20C),
				.b7(W3J21C),
				.b8(W3J22C),
				.c(c3C22J)
);

ninexnine_unit ninexnine_unit_6077(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3J00D),
				.b1(W3J01D),
				.b2(W3J02D),
				.b3(W3J10D),
				.b4(W3J11D),
				.b5(W3J12D),
				.b6(W3J20D),
				.b7(W3J21D),
				.b8(W3J22D),
				.c(c3D22J)
);

ninexnine_unit ninexnine_unit_6078(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3J00E),
				.b1(W3J01E),
				.b2(W3J02E),
				.b3(W3J10E),
				.b4(W3J11E),
				.b5(W3J12E),
				.b6(W3J20E),
				.b7(W3J21E),
				.b8(W3J22E),
				.c(c3E22J)
);

ninexnine_unit ninexnine_unit_6079(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3J00F),
				.b1(W3J01F),
				.b2(W3J02F),
				.b3(W3J10F),
				.b4(W3J11F),
				.b5(W3J12F),
				.b6(W3J20F),
				.b7(W3J21F),
				.b8(W3J22F),
				.c(c3F22J)
);

assign C322J=c3022J+c3122J+c3222J+c3322J+c3422J+c3522J+c3622J+c3722J+c3822J+c3922J+c3A22J+c3B22J+c3C22J+c3D22J+c3E22J+c3F22J;
assign A322J=(C322J>=0)?1:0;

assign P422J=A322J;

ninexnine_unit ninexnine_unit_6080(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3000K)
);

ninexnine_unit ninexnine_unit_6081(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3100K)
);

ninexnine_unit ninexnine_unit_6082(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3200K)
);

ninexnine_unit ninexnine_unit_6083(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3300K)
);

ninexnine_unit ninexnine_unit_6084(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3400K)
);

ninexnine_unit ninexnine_unit_6085(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3500K)
);

ninexnine_unit ninexnine_unit_6086(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3600K)
);

ninexnine_unit ninexnine_unit_6087(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3700K)
);

ninexnine_unit ninexnine_unit_6088(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3800K)
);

ninexnine_unit ninexnine_unit_6089(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3900K)
);

ninexnine_unit ninexnine_unit_6090(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A00K)
);

ninexnine_unit ninexnine_unit_6091(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B00K)
);

ninexnine_unit ninexnine_unit_6092(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C00K)
);

ninexnine_unit ninexnine_unit_6093(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D00K)
);

ninexnine_unit ninexnine_unit_6094(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E00K)
);

ninexnine_unit ninexnine_unit_6095(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F00K)
);

assign C300K=c3000K+c3100K+c3200K+c3300K+c3400K+c3500K+c3600K+c3700K+c3800K+c3900K+c3A00K+c3B00K+c3C00K+c3D00K+c3E00K+c3F00K;
assign A300K=(C300K>=0)?1:0;

assign P400K=A300K;

ninexnine_unit ninexnine_unit_6096(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3001K)
);

ninexnine_unit ninexnine_unit_6097(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3101K)
);

ninexnine_unit ninexnine_unit_6098(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3201K)
);

ninexnine_unit ninexnine_unit_6099(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3301K)
);

ninexnine_unit ninexnine_unit_6100(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3401K)
);

ninexnine_unit ninexnine_unit_6101(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3501K)
);

ninexnine_unit ninexnine_unit_6102(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3601K)
);

ninexnine_unit ninexnine_unit_6103(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3701K)
);

ninexnine_unit ninexnine_unit_6104(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3801K)
);

ninexnine_unit ninexnine_unit_6105(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3901K)
);

ninexnine_unit ninexnine_unit_6106(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A01K)
);

ninexnine_unit ninexnine_unit_6107(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B01K)
);

ninexnine_unit ninexnine_unit_6108(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C01K)
);

ninexnine_unit ninexnine_unit_6109(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D01K)
);

ninexnine_unit ninexnine_unit_6110(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E01K)
);

ninexnine_unit ninexnine_unit_6111(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F01K)
);

assign C301K=c3001K+c3101K+c3201K+c3301K+c3401K+c3501K+c3601K+c3701K+c3801K+c3901K+c3A01K+c3B01K+c3C01K+c3D01K+c3E01K+c3F01K;
assign A301K=(C301K>=0)?1:0;

assign P401K=A301K;

ninexnine_unit ninexnine_unit_6112(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3002K)
);

ninexnine_unit ninexnine_unit_6113(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3102K)
);

ninexnine_unit ninexnine_unit_6114(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3202K)
);

ninexnine_unit ninexnine_unit_6115(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3302K)
);

ninexnine_unit ninexnine_unit_6116(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3402K)
);

ninexnine_unit ninexnine_unit_6117(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3502K)
);

ninexnine_unit ninexnine_unit_6118(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3602K)
);

ninexnine_unit ninexnine_unit_6119(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3702K)
);

ninexnine_unit ninexnine_unit_6120(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3802K)
);

ninexnine_unit ninexnine_unit_6121(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3902K)
);

ninexnine_unit ninexnine_unit_6122(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A02K)
);

ninexnine_unit ninexnine_unit_6123(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B02K)
);

ninexnine_unit ninexnine_unit_6124(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C02K)
);

ninexnine_unit ninexnine_unit_6125(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D02K)
);

ninexnine_unit ninexnine_unit_6126(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E02K)
);

ninexnine_unit ninexnine_unit_6127(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F02K)
);

assign C302K=c3002K+c3102K+c3202K+c3302K+c3402K+c3502K+c3602K+c3702K+c3802K+c3902K+c3A02K+c3B02K+c3C02K+c3D02K+c3E02K+c3F02K;
assign A302K=(C302K>=0)?1:0;

assign P402K=A302K;

ninexnine_unit ninexnine_unit_6128(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3010K)
);

ninexnine_unit ninexnine_unit_6129(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3110K)
);

ninexnine_unit ninexnine_unit_6130(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3210K)
);

ninexnine_unit ninexnine_unit_6131(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3310K)
);

ninexnine_unit ninexnine_unit_6132(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3410K)
);

ninexnine_unit ninexnine_unit_6133(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3510K)
);

ninexnine_unit ninexnine_unit_6134(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3610K)
);

ninexnine_unit ninexnine_unit_6135(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3710K)
);

ninexnine_unit ninexnine_unit_6136(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3810K)
);

ninexnine_unit ninexnine_unit_6137(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3910K)
);

ninexnine_unit ninexnine_unit_6138(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A10K)
);

ninexnine_unit ninexnine_unit_6139(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B10K)
);

ninexnine_unit ninexnine_unit_6140(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C10K)
);

ninexnine_unit ninexnine_unit_6141(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D10K)
);

ninexnine_unit ninexnine_unit_6142(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E10K)
);

ninexnine_unit ninexnine_unit_6143(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F10K)
);

assign C310K=c3010K+c3110K+c3210K+c3310K+c3410K+c3510K+c3610K+c3710K+c3810K+c3910K+c3A10K+c3B10K+c3C10K+c3D10K+c3E10K+c3F10K;
assign A310K=(C310K>=0)?1:0;

assign P410K=A310K;

ninexnine_unit ninexnine_unit_6144(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3011K)
);

ninexnine_unit ninexnine_unit_6145(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3111K)
);

ninexnine_unit ninexnine_unit_6146(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3211K)
);

ninexnine_unit ninexnine_unit_6147(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3311K)
);

ninexnine_unit ninexnine_unit_6148(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3411K)
);

ninexnine_unit ninexnine_unit_6149(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3511K)
);

ninexnine_unit ninexnine_unit_6150(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3611K)
);

ninexnine_unit ninexnine_unit_6151(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3711K)
);

ninexnine_unit ninexnine_unit_6152(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3811K)
);

ninexnine_unit ninexnine_unit_6153(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3911K)
);

ninexnine_unit ninexnine_unit_6154(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A11K)
);

ninexnine_unit ninexnine_unit_6155(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B11K)
);

ninexnine_unit ninexnine_unit_6156(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C11K)
);

ninexnine_unit ninexnine_unit_6157(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D11K)
);

ninexnine_unit ninexnine_unit_6158(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E11K)
);

ninexnine_unit ninexnine_unit_6159(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F11K)
);

assign C311K=c3011K+c3111K+c3211K+c3311K+c3411K+c3511K+c3611K+c3711K+c3811K+c3911K+c3A11K+c3B11K+c3C11K+c3D11K+c3E11K+c3F11K;
assign A311K=(C311K>=0)?1:0;

assign P411K=A311K;

ninexnine_unit ninexnine_unit_6160(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3012K)
);

ninexnine_unit ninexnine_unit_6161(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3112K)
);

ninexnine_unit ninexnine_unit_6162(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3212K)
);

ninexnine_unit ninexnine_unit_6163(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3312K)
);

ninexnine_unit ninexnine_unit_6164(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3412K)
);

ninexnine_unit ninexnine_unit_6165(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3512K)
);

ninexnine_unit ninexnine_unit_6166(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3612K)
);

ninexnine_unit ninexnine_unit_6167(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3712K)
);

ninexnine_unit ninexnine_unit_6168(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3812K)
);

ninexnine_unit ninexnine_unit_6169(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3912K)
);

ninexnine_unit ninexnine_unit_6170(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A12K)
);

ninexnine_unit ninexnine_unit_6171(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B12K)
);

ninexnine_unit ninexnine_unit_6172(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C12K)
);

ninexnine_unit ninexnine_unit_6173(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D12K)
);

ninexnine_unit ninexnine_unit_6174(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E12K)
);

ninexnine_unit ninexnine_unit_6175(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F12K)
);

assign C312K=c3012K+c3112K+c3212K+c3312K+c3412K+c3512K+c3612K+c3712K+c3812K+c3912K+c3A12K+c3B12K+c3C12K+c3D12K+c3E12K+c3F12K;
assign A312K=(C312K>=0)?1:0;

assign P412K=A312K;

ninexnine_unit ninexnine_unit_6176(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3020K)
);

ninexnine_unit ninexnine_unit_6177(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3120K)
);

ninexnine_unit ninexnine_unit_6178(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3220K)
);

ninexnine_unit ninexnine_unit_6179(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3320K)
);

ninexnine_unit ninexnine_unit_6180(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3420K)
);

ninexnine_unit ninexnine_unit_6181(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3520K)
);

ninexnine_unit ninexnine_unit_6182(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3620K)
);

ninexnine_unit ninexnine_unit_6183(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3720K)
);

ninexnine_unit ninexnine_unit_6184(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3820K)
);

ninexnine_unit ninexnine_unit_6185(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3920K)
);

ninexnine_unit ninexnine_unit_6186(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A20K)
);

ninexnine_unit ninexnine_unit_6187(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B20K)
);

ninexnine_unit ninexnine_unit_6188(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C20K)
);

ninexnine_unit ninexnine_unit_6189(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D20K)
);

ninexnine_unit ninexnine_unit_6190(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E20K)
);

ninexnine_unit ninexnine_unit_6191(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F20K)
);

assign C320K=c3020K+c3120K+c3220K+c3320K+c3420K+c3520K+c3620K+c3720K+c3820K+c3920K+c3A20K+c3B20K+c3C20K+c3D20K+c3E20K+c3F20K;
assign A320K=(C320K>=0)?1:0;

assign P420K=A320K;

ninexnine_unit ninexnine_unit_6192(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3021K)
);

ninexnine_unit ninexnine_unit_6193(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3121K)
);

ninexnine_unit ninexnine_unit_6194(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3221K)
);

ninexnine_unit ninexnine_unit_6195(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3321K)
);

ninexnine_unit ninexnine_unit_6196(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3421K)
);

ninexnine_unit ninexnine_unit_6197(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3521K)
);

ninexnine_unit ninexnine_unit_6198(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3621K)
);

ninexnine_unit ninexnine_unit_6199(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3721K)
);

ninexnine_unit ninexnine_unit_6200(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3821K)
);

ninexnine_unit ninexnine_unit_6201(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3921K)
);

ninexnine_unit ninexnine_unit_6202(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A21K)
);

ninexnine_unit ninexnine_unit_6203(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B21K)
);

ninexnine_unit ninexnine_unit_6204(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C21K)
);

ninexnine_unit ninexnine_unit_6205(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D21K)
);

ninexnine_unit ninexnine_unit_6206(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E21K)
);

ninexnine_unit ninexnine_unit_6207(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F21K)
);

assign C321K=c3021K+c3121K+c3221K+c3321K+c3421K+c3521K+c3621K+c3721K+c3821K+c3921K+c3A21K+c3B21K+c3C21K+c3D21K+c3E21K+c3F21K;
assign A321K=(C321K>=0)?1:0;

assign P421K=A321K;

ninexnine_unit ninexnine_unit_6208(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3K000),
				.b1(W3K010),
				.b2(W3K020),
				.b3(W3K100),
				.b4(W3K110),
				.b5(W3K120),
				.b6(W3K200),
				.b7(W3K210),
				.b8(W3K220),
				.c(c3022K)
);

ninexnine_unit ninexnine_unit_6209(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3K001),
				.b1(W3K011),
				.b2(W3K021),
				.b3(W3K101),
				.b4(W3K111),
				.b5(W3K121),
				.b6(W3K201),
				.b7(W3K211),
				.b8(W3K221),
				.c(c3122K)
);

ninexnine_unit ninexnine_unit_6210(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3K002),
				.b1(W3K012),
				.b2(W3K022),
				.b3(W3K102),
				.b4(W3K112),
				.b5(W3K122),
				.b6(W3K202),
				.b7(W3K212),
				.b8(W3K222),
				.c(c3222K)
);

ninexnine_unit ninexnine_unit_6211(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3K003),
				.b1(W3K013),
				.b2(W3K023),
				.b3(W3K103),
				.b4(W3K113),
				.b5(W3K123),
				.b6(W3K203),
				.b7(W3K213),
				.b8(W3K223),
				.c(c3322K)
);

ninexnine_unit ninexnine_unit_6212(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3K004),
				.b1(W3K014),
				.b2(W3K024),
				.b3(W3K104),
				.b4(W3K114),
				.b5(W3K124),
				.b6(W3K204),
				.b7(W3K214),
				.b8(W3K224),
				.c(c3422K)
);

ninexnine_unit ninexnine_unit_6213(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3K005),
				.b1(W3K015),
				.b2(W3K025),
				.b3(W3K105),
				.b4(W3K115),
				.b5(W3K125),
				.b6(W3K205),
				.b7(W3K215),
				.b8(W3K225),
				.c(c3522K)
);

ninexnine_unit ninexnine_unit_6214(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3K006),
				.b1(W3K016),
				.b2(W3K026),
				.b3(W3K106),
				.b4(W3K116),
				.b5(W3K126),
				.b6(W3K206),
				.b7(W3K216),
				.b8(W3K226),
				.c(c3622K)
);

ninexnine_unit ninexnine_unit_6215(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3K007),
				.b1(W3K017),
				.b2(W3K027),
				.b3(W3K107),
				.b4(W3K117),
				.b5(W3K127),
				.b6(W3K207),
				.b7(W3K217),
				.b8(W3K227),
				.c(c3722K)
);

ninexnine_unit ninexnine_unit_6216(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3K008),
				.b1(W3K018),
				.b2(W3K028),
				.b3(W3K108),
				.b4(W3K118),
				.b5(W3K128),
				.b6(W3K208),
				.b7(W3K218),
				.b8(W3K228),
				.c(c3822K)
);

ninexnine_unit ninexnine_unit_6217(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3K009),
				.b1(W3K019),
				.b2(W3K029),
				.b3(W3K109),
				.b4(W3K119),
				.b5(W3K129),
				.b6(W3K209),
				.b7(W3K219),
				.b8(W3K229),
				.c(c3922K)
);

ninexnine_unit ninexnine_unit_6218(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3K00A),
				.b1(W3K01A),
				.b2(W3K02A),
				.b3(W3K10A),
				.b4(W3K11A),
				.b5(W3K12A),
				.b6(W3K20A),
				.b7(W3K21A),
				.b8(W3K22A),
				.c(c3A22K)
);

ninexnine_unit ninexnine_unit_6219(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3K00B),
				.b1(W3K01B),
				.b2(W3K02B),
				.b3(W3K10B),
				.b4(W3K11B),
				.b5(W3K12B),
				.b6(W3K20B),
				.b7(W3K21B),
				.b8(W3K22B),
				.c(c3B22K)
);

ninexnine_unit ninexnine_unit_6220(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3K00C),
				.b1(W3K01C),
				.b2(W3K02C),
				.b3(W3K10C),
				.b4(W3K11C),
				.b5(W3K12C),
				.b6(W3K20C),
				.b7(W3K21C),
				.b8(W3K22C),
				.c(c3C22K)
);

ninexnine_unit ninexnine_unit_6221(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3K00D),
				.b1(W3K01D),
				.b2(W3K02D),
				.b3(W3K10D),
				.b4(W3K11D),
				.b5(W3K12D),
				.b6(W3K20D),
				.b7(W3K21D),
				.b8(W3K22D),
				.c(c3D22K)
);

ninexnine_unit ninexnine_unit_6222(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3K00E),
				.b1(W3K01E),
				.b2(W3K02E),
				.b3(W3K10E),
				.b4(W3K11E),
				.b5(W3K12E),
				.b6(W3K20E),
				.b7(W3K21E),
				.b8(W3K22E),
				.c(c3E22K)
);

ninexnine_unit ninexnine_unit_6223(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3K00F),
				.b1(W3K01F),
				.b2(W3K02F),
				.b3(W3K10F),
				.b4(W3K11F),
				.b5(W3K12F),
				.b6(W3K20F),
				.b7(W3K21F),
				.b8(W3K22F),
				.c(c3F22K)
);

assign C322K=c3022K+c3122K+c3222K+c3322K+c3422K+c3522K+c3622K+c3722K+c3822K+c3922K+c3A22K+c3B22K+c3C22K+c3D22K+c3E22K+c3F22K;
assign A322K=(C322K>=0)?1:0;

assign P422K=A322K;

ninexnine_unit ninexnine_unit_6224(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3000L)
);

ninexnine_unit ninexnine_unit_6225(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3100L)
);

ninexnine_unit ninexnine_unit_6226(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3200L)
);

ninexnine_unit ninexnine_unit_6227(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3300L)
);

ninexnine_unit ninexnine_unit_6228(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3400L)
);

ninexnine_unit ninexnine_unit_6229(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3500L)
);

ninexnine_unit ninexnine_unit_6230(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3600L)
);

ninexnine_unit ninexnine_unit_6231(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3700L)
);

ninexnine_unit ninexnine_unit_6232(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3800L)
);

ninexnine_unit ninexnine_unit_6233(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3900L)
);

ninexnine_unit ninexnine_unit_6234(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A00L)
);

ninexnine_unit ninexnine_unit_6235(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B00L)
);

ninexnine_unit ninexnine_unit_6236(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C00L)
);

ninexnine_unit ninexnine_unit_6237(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D00L)
);

ninexnine_unit ninexnine_unit_6238(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E00L)
);

ninexnine_unit ninexnine_unit_6239(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F00L)
);

assign C300L=c3000L+c3100L+c3200L+c3300L+c3400L+c3500L+c3600L+c3700L+c3800L+c3900L+c3A00L+c3B00L+c3C00L+c3D00L+c3E00L+c3F00L;
assign A300L=(C300L>=0)?1:0;

assign P400L=A300L;

ninexnine_unit ninexnine_unit_6240(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3001L)
);

ninexnine_unit ninexnine_unit_6241(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3101L)
);

ninexnine_unit ninexnine_unit_6242(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3201L)
);

ninexnine_unit ninexnine_unit_6243(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3301L)
);

ninexnine_unit ninexnine_unit_6244(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3401L)
);

ninexnine_unit ninexnine_unit_6245(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3501L)
);

ninexnine_unit ninexnine_unit_6246(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3601L)
);

ninexnine_unit ninexnine_unit_6247(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3701L)
);

ninexnine_unit ninexnine_unit_6248(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3801L)
);

ninexnine_unit ninexnine_unit_6249(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3901L)
);

ninexnine_unit ninexnine_unit_6250(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A01L)
);

ninexnine_unit ninexnine_unit_6251(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B01L)
);

ninexnine_unit ninexnine_unit_6252(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C01L)
);

ninexnine_unit ninexnine_unit_6253(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D01L)
);

ninexnine_unit ninexnine_unit_6254(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E01L)
);

ninexnine_unit ninexnine_unit_6255(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F01L)
);

assign C301L=c3001L+c3101L+c3201L+c3301L+c3401L+c3501L+c3601L+c3701L+c3801L+c3901L+c3A01L+c3B01L+c3C01L+c3D01L+c3E01L+c3F01L;
assign A301L=(C301L>=0)?1:0;

assign P401L=A301L;

ninexnine_unit ninexnine_unit_6256(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3002L)
);

ninexnine_unit ninexnine_unit_6257(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3102L)
);

ninexnine_unit ninexnine_unit_6258(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3202L)
);

ninexnine_unit ninexnine_unit_6259(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3302L)
);

ninexnine_unit ninexnine_unit_6260(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3402L)
);

ninexnine_unit ninexnine_unit_6261(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3502L)
);

ninexnine_unit ninexnine_unit_6262(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3602L)
);

ninexnine_unit ninexnine_unit_6263(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3702L)
);

ninexnine_unit ninexnine_unit_6264(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3802L)
);

ninexnine_unit ninexnine_unit_6265(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3902L)
);

ninexnine_unit ninexnine_unit_6266(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A02L)
);

ninexnine_unit ninexnine_unit_6267(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B02L)
);

ninexnine_unit ninexnine_unit_6268(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C02L)
);

ninexnine_unit ninexnine_unit_6269(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D02L)
);

ninexnine_unit ninexnine_unit_6270(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E02L)
);

ninexnine_unit ninexnine_unit_6271(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F02L)
);

assign C302L=c3002L+c3102L+c3202L+c3302L+c3402L+c3502L+c3602L+c3702L+c3802L+c3902L+c3A02L+c3B02L+c3C02L+c3D02L+c3E02L+c3F02L;
assign A302L=(C302L>=0)?1:0;

assign P402L=A302L;

ninexnine_unit ninexnine_unit_6272(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3010L)
);

ninexnine_unit ninexnine_unit_6273(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3110L)
);

ninexnine_unit ninexnine_unit_6274(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3210L)
);

ninexnine_unit ninexnine_unit_6275(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3310L)
);

ninexnine_unit ninexnine_unit_6276(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3410L)
);

ninexnine_unit ninexnine_unit_6277(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3510L)
);

ninexnine_unit ninexnine_unit_6278(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3610L)
);

ninexnine_unit ninexnine_unit_6279(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3710L)
);

ninexnine_unit ninexnine_unit_6280(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3810L)
);

ninexnine_unit ninexnine_unit_6281(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3910L)
);

ninexnine_unit ninexnine_unit_6282(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A10L)
);

ninexnine_unit ninexnine_unit_6283(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B10L)
);

ninexnine_unit ninexnine_unit_6284(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C10L)
);

ninexnine_unit ninexnine_unit_6285(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D10L)
);

ninexnine_unit ninexnine_unit_6286(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E10L)
);

ninexnine_unit ninexnine_unit_6287(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F10L)
);

assign C310L=c3010L+c3110L+c3210L+c3310L+c3410L+c3510L+c3610L+c3710L+c3810L+c3910L+c3A10L+c3B10L+c3C10L+c3D10L+c3E10L+c3F10L;
assign A310L=(C310L>=0)?1:0;

assign P410L=A310L;

ninexnine_unit ninexnine_unit_6288(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3011L)
);

ninexnine_unit ninexnine_unit_6289(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3111L)
);

ninexnine_unit ninexnine_unit_6290(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3211L)
);

ninexnine_unit ninexnine_unit_6291(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3311L)
);

ninexnine_unit ninexnine_unit_6292(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3411L)
);

ninexnine_unit ninexnine_unit_6293(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3511L)
);

ninexnine_unit ninexnine_unit_6294(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3611L)
);

ninexnine_unit ninexnine_unit_6295(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3711L)
);

ninexnine_unit ninexnine_unit_6296(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3811L)
);

ninexnine_unit ninexnine_unit_6297(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3911L)
);

ninexnine_unit ninexnine_unit_6298(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A11L)
);

ninexnine_unit ninexnine_unit_6299(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B11L)
);

ninexnine_unit ninexnine_unit_6300(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C11L)
);

ninexnine_unit ninexnine_unit_6301(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D11L)
);

ninexnine_unit ninexnine_unit_6302(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E11L)
);

ninexnine_unit ninexnine_unit_6303(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F11L)
);

assign C311L=c3011L+c3111L+c3211L+c3311L+c3411L+c3511L+c3611L+c3711L+c3811L+c3911L+c3A11L+c3B11L+c3C11L+c3D11L+c3E11L+c3F11L;
assign A311L=(C311L>=0)?1:0;

assign P411L=A311L;

ninexnine_unit ninexnine_unit_6304(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3012L)
);

ninexnine_unit ninexnine_unit_6305(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3112L)
);

ninexnine_unit ninexnine_unit_6306(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3212L)
);

ninexnine_unit ninexnine_unit_6307(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3312L)
);

ninexnine_unit ninexnine_unit_6308(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3412L)
);

ninexnine_unit ninexnine_unit_6309(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3512L)
);

ninexnine_unit ninexnine_unit_6310(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3612L)
);

ninexnine_unit ninexnine_unit_6311(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3712L)
);

ninexnine_unit ninexnine_unit_6312(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3812L)
);

ninexnine_unit ninexnine_unit_6313(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3912L)
);

ninexnine_unit ninexnine_unit_6314(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A12L)
);

ninexnine_unit ninexnine_unit_6315(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B12L)
);

ninexnine_unit ninexnine_unit_6316(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C12L)
);

ninexnine_unit ninexnine_unit_6317(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D12L)
);

ninexnine_unit ninexnine_unit_6318(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E12L)
);

ninexnine_unit ninexnine_unit_6319(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F12L)
);

assign C312L=c3012L+c3112L+c3212L+c3312L+c3412L+c3512L+c3612L+c3712L+c3812L+c3912L+c3A12L+c3B12L+c3C12L+c3D12L+c3E12L+c3F12L;
assign A312L=(C312L>=0)?1:0;

assign P412L=A312L;

ninexnine_unit ninexnine_unit_6320(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3020L)
);

ninexnine_unit ninexnine_unit_6321(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3120L)
);

ninexnine_unit ninexnine_unit_6322(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3220L)
);

ninexnine_unit ninexnine_unit_6323(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3320L)
);

ninexnine_unit ninexnine_unit_6324(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3420L)
);

ninexnine_unit ninexnine_unit_6325(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3520L)
);

ninexnine_unit ninexnine_unit_6326(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3620L)
);

ninexnine_unit ninexnine_unit_6327(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3720L)
);

ninexnine_unit ninexnine_unit_6328(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3820L)
);

ninexnine_unit ninexnine_unit_6329(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3920L)
);

ninexnine_unit ninexnine_unit_6330(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A20L)
);

ninexnine_unit ninexnine_unit_6331(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B20L)
);

ninexnine_unit ninexnine_unit_6332(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C20L)
);

ninexnine_unit ninexnine_unit_6333(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D20L)
);

ninexnine_unit ninexnine_unit_6334(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E20L)
);

ninexnine_unit ninexnine_unit_6335(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F20L)
);

assign C320L=c3020L+c3120L+c3220L+c3320L+c3420L+c3520L+c3620L+c3720L+c3820L+c3920L+c3A20L+c3B20L+c3C20L+c3D20L+c3E20L+c3F20L;
assign A320L=(C320L>=0)?1:0;

assign P420L=A320L;

ninexnine_unit ninexnine_unit_6336(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3021L)
);

ninexnine_unit ninexnine_unit_6337(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3121L)
);

ninexnine_unit ninexnine_unit_6338(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3221L)
);

ninexnine_unit ninexnine_unit_6339(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3321L)
);

ninexnine_unit ninexnine_unit_6340(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3421L)
);

ninexnine_unit ninexnine_unit_6341(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3521L)
);

ninexnine_unit ninexnine_unit_6342(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3621L)
);

ninexnine_unit ninexnine_unit_6343(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3721L)
);

ninexnine_unit ninexnine_unit_6344(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3821L)
);

ninexnine_unit ninexnine_unit_6345(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3921L)
);

ninexnine_unit ninexnine_unit_6346(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A21L)
);

ninexnine_unit ninexnine_unit_6347(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B21L)
);

ninexnine_unit ninexnine_unit_6348(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C21L)
);

ninexnine_unit ninexnine_unit_6349(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D21L)
);

ninexnine_unit ninexnine_unit_6350(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E21L)
);

ninexnine_unit ninexnine_unit_6351(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F21L)
);

assign C321L=c3021L+c3121L+c3221L+c3321L+c3421L+c3521L+c3621L+c3721L+c3821L+c3921L+c3A21L+c3B21L+c3C21L+c3D21L+c3E21L+c3F21L;
assign A321L=(C321L>=0)?1:0;

assign P421L=A321L;

ninexnine_unit ninexnine_unit_6352(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3L000),
				.b1(W3L010),
				.b2(W3L020),
				.b3(W3L100),
				.b4(W3L110),
				.b5(W3L120),
				.b6(W3L200),
				.b7(W3L210),
				.b8(W3L220),
				.c(c3022L)
);

ninexnine_unit ninexnine_unit_6353(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3L001),
				.b1(W3L011),
				.b2(W3L021),
				.b3(W3L101),
				.b4(W3L111),
				.b5(W3L121),
				.b6(W3L201),
				.b7(W3L211),
				.b8(W3L221),
				.c(c3122L)
);

ninexnine_unit ninexnine_unit_6354(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3L002),
				.b1(W3L012),
				.b2(W3L022),
				.b3(W3L102),
				.b4(W3L112),
				.b5(W3L122),
				.b6(W3L202),
				.b7(W3L212),
				.b8(W3L222),
				.c(c3222L)
);

ninexnine_unit ninexnine_unit_6355(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3L003),
				.b1(W3L013),
				.b2(W3L023),
				.b3(W3L103),
				.b4(W3L113),
				.b5(W3L123),
				.b6(W3L203),
				.b7(W3L213),
				.b8(W3L223),
				.c(c3322L)
);

ninexnine_unit ninexnine_unit_6356(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3L004),
				.b1(W3L014),
				.b2(W3L024),
				.b3(W3L104),
				.b4(W3L114),
				.b5(W3L124),
				.b6(W3L204),
				.b7(W3L214),
				.b8(W3L224),
				.c(c3422L)
);

ninexnine_unit ninexnine_unit_6357(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3L005),
				.b1(W3L015),
				.b2(W3L025),
				.b3(W3L105),
				.b4(W3L115),
				.b5(W3L125),
				.b6(W3L205),
				.b7(W3L215),
				.b8(W3L225),
				.c(c3522L)
);

ninexnine_unit ninexnine_unit_6358(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3L006),
				.b1(W3L016),
				.b2(W3L026),
				.b3(W3L106),
				.b4(W3L116),
				.b5(W3L126),
				.b6(W3L206),
				.b7(W3L216),
				.b8(W3L226),
				.c(c3622L)
);

ninexnine_unit ninexnine_unit_6359(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3L007),
				.b1(W3L017),
				.b2(W3L027),
				.b3(W3L107),
				.b4(W3L117),
				.b5(W3L127),
				.b6(W3L207),
				.b7(W3L217),
				.b8(W3L227),
				.c(c3722L)
);

ninexnine_unit ninexnine_unit_6360(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3L008),
				.b1(W3L018),
				.b2(W3L028),
				.b3(W3L108),
				.b4(W3L118),
				.b5(W3L128),
				.b6(W3L208),
				.b7(W3L218),
				.b8(W3L228),
				.c(c3822L)
);

ninexnine_unit ninexnine_unit_6361(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3L009),
				.b1(W3L019),
				.b2(W3L029),
				.b3(W3L109),
				.b4(W3L119),
				.b5(W3L129),
				.b6(W3L209),
				.b7(W3L219),
				.b8(W3L229),
				.c(c3922L)
);

ninexnine_unit ninexnine_unit_6362(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3L00A),
				.b1(W3L01A),
				.b2(W3L02A),
				.b3(W3L10A),
				.b4(W3L11A),
				.b5(W3L12A),
				.b6(W3L20A),
				.b7(W3L21A),
				.b8(W3L22A),
				.c(c3A22L)
);

ninexnine_unit ninexnine_unit_6363(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3L00B),
				.b1(W3L01B),
				.b2(W3L02B),
				.b3(W3L10B),
				.b4(W3L11B),
				.b5(W3L12B),
				.b6(W3L20B),
				.b7(W3L21B),
				.b8(W3L22B),
				.c(c3B22L)
);

ninexnine_unit ninexnine_unit_6364(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3L00C),
				.b1(W3L01C),
				.b2(W3L02C),
				.b3(W3L10C),
				.b4(W3L11C),
				.b5(W3L12C),
				.b6(W3L20C),
				.b7(W3L21C),
				.b8(W3L22C),
				.c(c3C22L)
);

ninexnine_unit ninexnine_unit_6365(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3L00D),
				.b1(W3L01D),
				.b2(W3L02D),
				.b3(W3L10D),
				.b4(W3L11D),
				.b5(W3L12D),
				.b6(W3L20D),
				.b7(W3L21D),
				.b8(W3L22D),
				.c(c3D22L)
);

ninexnine_unit ninexnine_unit_6366(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3L00E),
				.b1(W3L01E),
				.b2(W3L02E),
				.b3(W3L10E),
				.b4(W3L11E),
				.b5(W3L12E),
				.b6(W3L20E),
				.b7(W3L21E),
				.b8(W3L22E),
				.c(c3E22L)
);

ninexnine_unit ninexnine_unit_6367(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3L00F),
				.b1(W3L01F),
				.b2(W3L02F),
				.b3(W3L10F),
				.b4(W3L11F),
				.b5(W3L12F),
				.b6(W3L20F),
				.b7(W3L21F),
				.b8(W3L22F),
				.c(c3F22L)
);

assign C322L=c3022L+c3122L+c3222L+c3322L+c3422L+c3522L+c3622L+c3722L+c3822L+c3922L+c3A22L+c3B22L+c3C22L+c3D22L+c3E22L+c3F22L;
assign A322L=(C322L>=0)?1:0;

assign P422L=A322L;

ninexnine_unit ninexnine_unit_6368(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3000M)
);

ninexnine_unit ninexnine_unit_6369(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3100M)
);

ninexnine_unit ninexnine_unit_6370(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3200M)
);

ninexnine_unit ninexnine_unit_6371(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3300M)
);

ninexnine_unit ninexnine_unit_6372(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3400M)
);

ninexnine_unit ninexnine_unit_6373(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3500M)
);

ninexnine_unit ninexnine_unit_6374(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3600M)
);

ninexnine_unit ninexnine_unit_6375(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3700M)
);

ninexnine_unit ninexnine_unit_6376(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3800M)
);

ninexnine_unit ninexnine_unit_6377(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3900M)
);

ninexnine_unit ninexnine_unit_6378(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A00M)
);

ninexnine_unit ninexnine_unit_6379(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B00M)
);

ninexnine_unit ninexnine_unit_6380(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C00M)
);

ninexnine_unit ninexnine_unit_6381(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D00M)
);

ninexnine_unit ninexnine_unit_6382(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E00M)
);

ninexnine_unit ninexnine_unit_6383(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F00M)
);

assign C300M=c3000M+c3100M+c3200M+c3300M+c3400M+c3500M+c3600M+c3700M+c3800M+c3900M+c3A00M+c3B00M+c3C00M+c3D00M+c3E00M+c3F00M;
assign A300M=(C300M>=0)?1:0;

assign P400M=A300M;

ninexnine_unit ninexnine_unit_6384(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3001M)
);

ninexnine_unit ninexnine_unit_6385(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3101M)
);

ninexnine_unit ninexnine_unit_6386(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3201M)
);

ninexnine_unit ninexnine_unit_6387(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3301M)
);

ninexnine_unit ninexnine_unit_6388(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3401M)
);

ninexnine_unit ninexnine_unit_6389(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3501M)
);

ninexnine_unit ninexnine_unit_6390(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3601M)
);

ninexnine_unit ninexnine_unit_6391(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3701M)
);

ninexnine_unit ninexnine_unit_6392(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3801M)
);

ninexnine_unit ninexnine_unit_6393(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3901M)
);

ninexnine_unit ninexnine_unit_6394(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A01M)
);

ninexnine_unit ninexnine_unit_6395(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B01M)
);

ninexnine_unit ninexnine_unit_6396(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C01M)
);

ninexnine_unit ninexnine_unit_6397(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D01M)
);

ninexnine_unit ninexnine_unit_6398(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E01M)
);

ninexnine_unit ninexnine_unit_6399(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F01M)
);

assign C301M=c3001M+c3101M+c3201M+c3301M+c3401M+c3501M+c3601M+c3701M+c3801M+c3901M+c3A01M+c3B01M+c3C01M+c3D01M+c3E01M+c3F01M;
assign A301M=(C301M>=0)?1:0;

assign P401M=A301M;

ninexnine_unit ninexnine_unit_6400(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3002M)
);

ninexnine_unit ninexnine_unit_6401(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3102M)
);

ninexnine_unit ninexnine_unit_6402(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3202M)
);

ninexnine_unit ninexnine_unit_6403(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3302M)
);

ninexnine_unit ninexnine_unit_6404(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3402M)
);

ninexnine_unit ninexnine_unit_6405(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3502M)
);

ninexnine_unit ninexnine_unit_6406(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3602M)
);

ninexnine_unit ninexnine_unit_6407(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3702M)
);

ninexnine_unit ninexnine_unit_6408(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3802M)
);

ninexnine_unit ninexnine_unit_6409(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3902M)
);

ninexnine_unit ninexnine_unit_6410(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A02M)
);

ninexnine_unit ninexnine_unit_6411(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B02M)
);

ninexnine_unit ninexnine_unit_6412(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C02M)
);

ninexnine_unit ninexnine_unit_6413(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D02M)
);

ninexnine_unit ninexnine_unit_6414(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E02M)
);

ninexnine_unit ninexnine_unit_6415(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F02M)
);

assign C302M=c3002M+c3102M+c3202M+c3302M+c3402M+c3502M+c3602M+c3702M+c3802M+c3902M+c3A02M+c3B02M+c3C02M+c3D02M+c3E02M+c3F02M;
assign A302M=(C302M>=0)?1:0;

assign P402M=A302M;

ninexnine_unit ninexnine_unit_6416(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3010M)
);

ninexnine_unit ninexnine_unit_6417(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3110M)
);

ninexnine_unit ninexnine_unit_6418(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3210M)
);

ninexnine_unit ninexnine_unit_6419(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3310M)
);

ninexnine_unit ninexnine_unit_6420(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3410M)
);

ninexnine_unit ninexnine_unit_6421(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3510M)
);

ninexnine_unit ninexnine_unit_6422(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3610M)
);

ninexnine_unit ninexnine_unit_6423(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3710M)
);

ninexnine_unit ninexnine_unit_6424(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3810M)
);

ninexnine_unit ninexnine_unit_6425(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3910M)
);

ninexnine_unit ninexnine_unit_6426(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A10M)
);

ninexnine_unit ninexnine_unit_6427(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B10M)
);

ninexnine_unit ninexnine_unit_6428(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C10M)
);

ninexnine_unit ninexnine_unit_6429(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D10M)
);

ninexnine_unit ninexnine_unit_6430(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E10M)
);

ninexnine_unit ninexnine_unit_6431(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F10M)
);

assign C310M=c3010M+c3110M+c3210M+c3310M+c3410M+c3510M+c3610M+c3710M+c3810M+c3910M+c3A10M+c3B10M+c3C10M+c3D10M+c3E10M+c3F10M;
assign A310M=(C310M>=0)?1:0;

assign P410M=A310M;

ninexnine_unit ninexnine_unit_6432(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3011M)
);

ninexnine_unit ninexnine_unit_6433(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3111M)
);

ninexnine_unit ninexnine_unit_6434(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3211M)
);

ninexnine_unit ninexnine_unit_6435(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3311M)
);

ninexnine_unit ninexnine_unit_6436(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3411M)
);

ninexnine_unit ninexnine_unit_6437(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3511M)
);

ninexnine_unit ninexnine_unit_6438(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3611M)
);

ninexnine_unit ninexnine_unit_6439(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3711M)
);

ninexnine_unit ninexnine_unit_6440(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3811M)
);

ninexnine_unit ninexnine_unit_6441(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3911M)
);

ninexnine_unit ninexnine_unit_6442(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A11M)
);

ninexnine_unit ninexnine_unit_6443(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B11M)
);

ninexnine_unit ninexnine_unit_6444(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C11M)
);

ninexnine_unit ninexnine_unit_6445(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D11M)
);

ninexnine_unit ninexnine_unit_6446(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E11M)
);

ninexnine_unit ninexnine_unit_6447(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F11M)
);

assign C311M=c3011M+c3111M+c3211M+c3311M+c3411M+c3511M+c3611M+c3711M+c3811M+c3911M+c3A11M+c3B11M+c3C11M+c3D11M+c3E11M+c3F11M;
assign A311M=(C311M>=0)?1:0;

assign P411M=A311M;

ninexnine_unit ninexnine_unit_6448(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3012M)
);

ninexnine_unit ninexnine_unit_6449(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3112M)
);

ninexnine_unit ninexnine_unit_6450(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3212M)
);

ninexnine_unit ninexnine_unit_6451(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3312M)
);

ninexnine_unit ninexnine_unit_6452(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3412M)
);

ninexnine_unit ninexnine_unit_6453(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3512M)
);

ninexnine_unit ninexnine_unit_6454(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3612M)
);

ninexnine_unit ninexnine_unit_6455(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3712M)
);

ninexnine_unit ninexnine_unit_6456(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3812M)
);

ninexnine_unit ninexnine_unit_6457(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3912M)
);

ninexnine_unit ninexnine_unit_6458(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A12M)
);

ninexnine_unit ninexnine_unit_6459(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B12M)
);

ninexnine_unit ninexnine_unit_6460(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C12M)
);

ninexnine_unit ninexnine_unit_6461(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D12M)
);

ninexnine_unit ninexnine_unit_6462(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E12M)
);

ninexnine_unit ninexnine_unit_6463(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F12M)
);

assign C312M=c3012M+c3112M+c3212M+c3312M+c3412M+c3512M+c3612M+c3712M+c3812M+c3912M+c3A12M+c3B12M+c3C12M+c3D12M+c3E12M+c3F12M;
assign A312M=(C312M>=0)?1:0;

assign P412M=A312M;

ninexnine_unit ninexnine_unit_6464(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3020M)
);

ninexnine_unit ninexnine_unit_6465(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3120M)
);

ninexnine_unit ninexnine_unit_6466(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3220M)
);

ninexnine_unit ninexnine_unit_6467(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3320M)
);

ninexnine_unit ninexnine_unit_6468(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3420M)
);

ninexnine_unit ninexnine_unit_6469(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3520M)
);

ninexnine_unit ninexnine_unit_6470(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3620M)
);

ninexnine_unit ninexnine_unit_6471(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3720M)
);

ninexnine_unit ninexnine_unit_6472(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3820M)
);

ninexnine_unit ninexnine_unit_6473(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3920M)
);

ninexnine_unit ninexnine_unit_6474(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A20M)
);

ninexnine_unit ninexnine_unit_6475(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B20M)
);

ninexnine_unit ninexnine_unit_6476(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C20M)
);

ninexnine_unit ninexnine_unit_6477(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D20M)
);

ninexnine_unit ninexnine_unit_6478(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E20M)
);

ninexnine_unit ninexnine_unit_6479(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F20M)
);

assign C320M=c3020M+c3120M+c3220M+c3320M+c3420M+c3520M+c3620M+c3720M+c3820M+c3920M+c3A20M+c3B20M+c3C20M+c3D20M+c3E20M+c3F20M;
assign A320M=(C320M>=0)?1:0;

assign P420M=A320M;

ninexnine_unit ninexnine_unit_6480(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3021M)
);

ninexnine_unit ninexnine_unit_6481(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3121M)
);

ninexnine_unit ninexnine_unit_6482(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3221M)
);

ninexnine_unit ninexnine_unit_6483(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3321M)
);

ninexnine_unit ninexnine_unit_6484(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3421M)
);

ninexnine_unit ninexnine_unit_6485(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3521M)
);

ninexnine_unit ninexnine_unit_6486(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3621M)
);

ninexnine_unit ninexnine_unit_6487(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3721M)
);

ninexnine_unit ninexnine_unit_6488(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3821M)
);

ninexnine_unit ninexnine_unit_6489(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3921M)
);

ninexnine_unit ninexnine_unit_6490(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A21M)
);

ninexnine_unit ninexnine_unit_6491(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B21M)
);

ninexnine_unit ninexnine_unit_6492(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C21M)
);

ninexnine_unit ninexnine_unit_6493(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D21M)
);

ninexnine_unit ninexnine_unit_6494(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E21M)
);

ninexnine_unit ninexnine_unit_6495(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F21M)
);

assign C321M=c3021M+c3121M+c3221M+c3321M+c3421M+c3521M+c3621M+c3721M+c3821M+c3921M+c3A21M+c3B21M+c3C21M+c3D21M+c3E21M+c3F21M;
assign A321M=(C321M>=0)?1:0;

assign P421M=A321M;

ninexnine_unit ninexnine_unit_6496(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3M000),
				.b1(W3M010),
				.b2(W3M020),
				.b3(W3M100),
				.b4(W3M110),
				.b5(W3M120),
				.b6(W3M200),
				.b7(W3M210),
				.b8(W3M220),
				.c(c3022M)
);

ninexnine_unit ninexnine_unit_6497(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3M001),
				.b1(W3M011),
				.b2(W3M021),
				.b3(W3M101),
				.b4(W3M111),
				.b5(W3M121),
				.b6(W3M201),
				.b7(W3M211),
				.b8(W3M221),
				.c(c3122M)
);

ninexnine_unit ninexnine_unit_6498(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3M002),
				.b1(W3M012),
				.b2(W3M022),
				.b3(W3M102),
				.b4(W3M112),
				.b5(W3M122),
				.b6(W3M202),
				.b7(W3M212),
				.b8(W3M222),
				.c(c3222M)
);

ninexnine_unit ninexnine_unit_6499(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3M003),
				.b1(W3M013),
				.b2(W3M023),
				.b3(W3M103),
				.b4(W3M113),
				.b5(W3M123),
				.b6(W3M203),
				.b7(W3M213),
				.b8(W3M223),
				.c(c3322M)
);

ninexnine_unit ninexnine_unit_6500(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3M004),
				.b1(W3M014),
				.b2(W3M024),
				.b3(W3M104),
				.b4(W3M114),
				.b5(W3M124),
				.b6(W3M204),
				.b7(W3M214),
				.b8(W3M224),
				.c(c3422M)
);

ninexnine_unit ninexnine_unit_6501(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3M005),
				.b1(W3M015),
				.b2(W3M025),
				.b3(W3M105),
				.b4(W3M115),
				.b5(W3M125),
				.b6(W3M205),
				.b7(W3M215),
				.b8(W3M225),
				.c(c3522M)
);

ninexnine_unit ninexnine_unit_6502(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3M006),
				.b1(W3M016),
				.b2(W3M026),
				.b3(W3M106),
				.b4(W3M116),
				.b5(W3M126),
				.b6(W3M206),
				.b7(W3M216),
				.b8(W3M226),
				.c(c3622M)
);

ninexnine_unit ninexnine_unit_6503(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3M007),
				.b1(W3M017),
				.b2(W3M027),
				.b3(W3M107),
				.b4(W3M117),
				.b5(W3M127),
				.b6(W3M207),
				.b7(W3M217),
				.b8(W3M227),
				.c(c3722M)
);

ninexnine_unit ninexnine_unit_6504(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3M008),
				.b1(W3M018),
				.b2(W3M028),
				.b3(W3M108),
				.b4(W3M118),
				.b5(W3M128),
				.b6(W3M208),
				.b7(W3M218),
				.b8(W3M228),
				.c(c3822M)
);

ninexnine_unit ninexnine_unit_6505(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3M009),
				.b1(W3M019),
				.b2(W3M029),
				.b3(W3M109),
				.b4(W3M119),
				.b5(W3M129),
				.b6(W3M209),
				.b7(W3M219),
				.b8(W3M229),
				.c(c3922M)
);

ninexnine_unit ninexnine_unit_6506(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3M00A),
				.b1(W3M01A),
				.b2(W3M02A),
				.b3(W3M10A),
				.b4(W3M11A),
				.b5(W3M12A),
				.b6(W3M20A),
				.b7(W3M21A),
				.b8(W3M22A),
				.c(c3A22M)
);

ninexnine_unit ninexnine_unit_6507(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3M00B),
				.b1(W3M01B),
				.b2(W3M02B),
				.b3(W3M10B),
				.b4(W3M11B),
				.b5(W3M12B),
				.b6(W3M20B),
				.b7(W3M21B),
				.b8(W3M22B),
				.c(c3B22M)
);

ninexnine_unit ninexnine_unit_6508(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3M00C),
				.b1(W3M01C),
				.b2(W3M02C),
				.b3(W3M10C),
				.b4(W3M11C),
				.b5(W3M12C),
				.b6(W3M20C),
				.b7(W3M21C),
				.b8(W3M22C),
				.c(c3C22M)
);

ninexnine_unit ninexnine_unit_6509(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3M00D),
				.b1(W3M01D),
				.b2(W3M02D),
				.b3(W3M10D),
				.b4(W3M11D),
				.b5(W3M12D),
				.b6(W3M20D),
				.b7(W3M21D),
				.b8(W3M22D),
				.c(c3D22M)
);

ninexnine_unit ninexnine_unit_6510(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3M00E),
				.b1(W3M01E),
				.b2(W3M02E),
				.b3(W3M10E),
				.b4(W3M11E),
				.b5(W3M12E),
				.b6(W3M20E),
				.b7(W3M21E),
				.b8(W3M22E),
				.c(c3E22M)
);

ninexnine_unit ninexnine_unit_6511(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3M00F),
				.b1(W3M01F),
				.b2(W3M02F),
				.b3(W3M10F),
				.b4(W3M11F),
				.b5(W3M12F),
				.b6(W3M20F),
				.b7(W3M21F),
				.b8(W3M22F),
				.c(c3F22M)
);

assign C322M=c3022M+c3122M+c3222M+c3322M+c3422M+c3522M+c3622M+c3722M+c3822M+c3922M+c3A22M+c3B22M+c3C22M+c3D22M+c3E22M+c3F22M;
assign A322M=(C322M>=0)?1:0;

assign P422M=A322M;

ninexnine_unit ninexnine_unit_6512(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3000N)
);

ninexnine_unit ninexnine_unit_6513(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3100N)
);

ninexnine_unit ninexnine_unit_6514(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3200N)
);

ninexnine_unit ninexnine_unit_6515(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3300N)
);

ninexnine_unit ninexnine_unit_6516(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3400N)
);

ninexnine_unit ninexnine_unit_6517(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3500N)
);

ninexnine_unit ninexnine_unit_6518(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3600N)
);

ninexnine_unit ninexnine_unit_6519(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3700N)
);

ninexnine_unit ninexnine_unit_6520(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3800N)
);

ninexnine_unit ninexnine_unit_6521(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3900N)
);

ninexnine_unit ninexnine_unit_6522(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A00N)
);

ninexnine_unit ninexnine_unit_6523(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B00N)
);

ninexnine_unit ninexnine_unit_6524(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C00N)
);

ninexnine_unit ninexnine_unit_6525(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D00N)
);

ninexnine_unit ninexnine_unit_6526(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E00N)
);

ninexnine_unit ninexnine_unit_6527(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F00N)
);

assign C300N=c3000N+c3100N+c3200N+c3300N+c3400N+c3500N+c3600N+c3700N+c3800N+c3900N+c3A00N+c3B00N+c3C00N+c3D00N+c3E00N+c3F00N;
assign A300N=(C300N>=0)?1:0;

assign P400N=A300N;

ninexnine_unit ninexnine_unit_6528(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3001N)
);

ninexnine_unit ninexnine_unit_6529(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3101N)
);

ninexnine_unit ninexnine_unit_6530(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3201N)
);

ninexnine_unit ninexnine_unit_6531(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3301N)
);

ninexnine_unit ninexnine_unit_6532(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3401N)
);

ninexnine_unit ninexnine_unit_6533(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3501N)
);

ninexnine_unit ninexnine_unit_6534(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3601N)
);

ninexnine_unit ninexnine_unit_6535(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3701N)
);

ninexnine_unit ninexnine_unit_6536(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3801N)
);

ninexnine_unit ninexnine_unit_6537(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3901N)
);

ninexnine_unit ninexnine_unit_6538(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A01N)
);

ninexnine_unit ninexnine_unit_6539(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B01N)
);

ninexnine_unit ninexnine_unit_6540(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C01N)
);

ninexnine_unit ninexnine_unit_6541(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D01N)
);

ninexnine_unit ninexnine_unit_6542(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E01N)
);

ninexnine_unit ninexnine_unit_6543(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F01N)
);

assign C301N=c3001N+c3101N+c3201N+c3301N+c3401N+c3501N+c3601N+c3701N+c3801N+c3901N+c3A01N+c3B01N+c3C01N+c3D01N+c3E01N+c3F01N;
assign A301N=(C301N>=0)?1:0;

assign P401N=A301N;

ninexnine_unit ninexnine_unit_6544(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3002N)
);

ninexnine_unit ninexnine_unit_6545(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3102N)
);

ninexnine_unit ninexnine_unit_6546(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3202N)
);

ninexnine_unit ninexnine_unit_6547(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3302N)
);

ninexnine_unit ninexnine_unit_6548(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3402N)
);

ninexnine_unit ninexnine_unit_6549(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3502N)
);

ninexnine_unit ninexnine_unit_6550(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3602N)
);

ninexnine_unit ninexnine_unit_6551(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3702N)
);

ninexnine_unit ninexnine_unit_6552(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3802N)
);

ninexnine_unit ninexnine_unit_6553(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3902N)
);

ninexnine_unit ninexnine_unit_6554(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A02N)
);

ninexnine_unit ninexnine_unit_6555(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B02N)
);

ninexnine_unit ninexnine_unit_6556(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C02N)
);

ninexnine_unit ninexnine_unit_6557(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D02N)
);

ninexnine_unit ninexnine_unit_6558(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E02N)
);

ninexnine_unit ninexnine_unit_6559(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F02N)
);

assign C302N=c3002N+c3102N+c3202N+c3302N+c3402N+c3502N+c3602N+c3702N+c3802N+c3902N+c3A02N+c3B02N+c3C02N+c3D02N+c3E02N+c3F02N;
assign A302N=(C302N>=0)?1:0;

assign P402N=A302N;

ninexnine_unit ninexnine_unit_6560(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3010N)
);

ninexnine_unit ninexnine_unit_6561(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3110N)
);

ninexnine_unit ninexnine_unit_6562(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3210N)
);

ninexnine_unit ninexnine_unit_6563(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3310N)
);

ninexnine_unit ninexnine_unit_6564(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3410N)
);

ninexnine_unit ninexnine_unit_6565(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3510N)
);

ninexnine_unit ninexnine_unit_6566(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3610N)
);

ninexnine_unit ninexnine_unit_6567(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3710N)
);

ninexnine_unit ninexnine_unit_6568(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3810N)
);

ninexnine_unit ninexnine_unit_6569(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3910N)
);

ninexnine_unit ninexnine_unit_6570(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A10N)
);

ninexnine_unit ninexnine_unit_6571(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B10N)
);

ninexnine_unit ninexnine_unit_6572(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C10N)
);

ninexnine_unit ninexnine_unit_6573(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D10N)
);

ninexnine_unit ninexnine_unit_6574(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E10N)
);

ninexnine_unit ninexnine_unit_6575(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F10N)
);

assign C310N=c3010N+c3110N+c3210N+c3310N+c3410N+c3510N+c3610N+c3710N+c3810N+c3910N+c3A10N+c3B10N+c3C10N+c3D10N+c3E10N+c3F10N;
assign A310N=(C310N>=0)?1:0;

assign P410N=A310N;

ninexnine_unit ninexnine_unit_6576(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3011N)
);

ninexnine_unit ninexnine_unit_6577(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3111N)
);

ninexnine_unit ninexnine_unit_6578(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3211N)
);

ninexnine_unit ninexnine_unit_6579(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3311N)
);

ninexnine_unit ninexnine_unit_6580(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3411N)
);

ninexnine_unit ninexnine_unit_6581(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3511N)
);

ninexnine_unit ninexnine_unit_6582(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3611N)
);

ninexnine_unit ninexnine_unit_6583(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3711N)
);

ninexnine_unit ninexnine_unit_6584(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3811N)
);

ninexnine_unit ninexnine_unit_6585(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3911N)
);

ninexnine_unit ninexnine_unit_6586(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A11N)
);

ninexnine_unit ninexnine_unit_6587(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B11N)
);

ninexnine_unit ninexnine_unit_6588(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C11N)
);

ninexnine_unit ninexnine_unit_6589(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D11N)
);

ninexnine_unit ninexnine_unit_6590(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E11N)
);

ninexnine_unit ninexnine_unit_6591(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F11N)
);

assign C311N=c3011N+c3111N+c3211N+c3311N+c3411N+c3511N+c3611N+c3711N+c3811N+c3911N+c3A11N+c3B11N+c3C11N+c3D11N+c3E11N+c3F11N;
assign A311N=(C311N>=0)?1:0;

assign P411N=A311N;

ninexnine_unit ninexnine_unit_6592(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3012N)
);

ninexnine_unit ninexnine_unit_6593(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3112N)
);

ninexnine_unit ninexnine_unit_6594(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3212N)
);

ninexnine_unit ninexnine_unit_6595(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3312N)
);

ninexnine_unit ninexnine_unit_6596(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3412N)
);

ninexnine_unit ninexnine_unit_6597(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3512N)
);

ninexnine_unit ninexnine_unit_6598(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3612N)
);

ninexnine_unit ninexnine_unit_6599(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3712N)
);

ninexnine_unit ninexnine_unit_6600(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3812N)
);

ninexnine_unit ninexnine_unit_6601(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3912N)
);

ninexnine_unit ninexnine_unit_6602(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A12N)
);

ninexnine_unit ninexnine_unit_6603(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B12N)
);

ninexnine_unit ninexnine_unit_6604(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C12N)
);

ninexnine_unit ninexnine_unit_6605(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D12N)
);

ninexnine_unit ninexnine_unit_6606(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E12N)
);

ninexnine_unit ninexnine_unit_6607(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F12N)
);

assign C312N=c3012N+c3112N+c3212N+c3312N+c3412N+c3512N+c3612N+c3712N+c3812N+c3912N+c3A12N+c3B12N+c3C12N+c3D12N+c3E12N+c3F12N;
assign A312N=(C312N>=0)?1:0;

assign P412N=A312N;

ninexnine_unit ninexnine_unit_6608(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3020N)
);

ninexnine_unit ninexnine_unit_6609(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3120N)
);

ninexnine_unit ninexnine_unit_6610(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3220N)
);

ninexnine_unit ninexnine_unit_6611(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3320N)
);

ninexnine_unit ninexnine_unit_6612(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3420N)
);

ninexnine_unit ninexnine_unit_6613(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3520N)
);

ninexnine_unit ninexnine_unit_6614(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3620N)
);

ninexnine_unit ninexnine_unit_6615(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3720N)
);

ninexnine_unit ninexnine_unit_6616(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3820N)
);

ninexnine_unit ninexnine_unit_6617(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3920N)
);

ninexnine_unit ninexnine_unit_6618(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A20N)
);

ninexnine_unit ninexnine_unit_6619(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B20N)
);

ninexnine_unit ninexnine_unit_6620(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C20N)
);

ninexnine_unit ninexnine_unit_6621(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D20N)
);

ninexnine_unit ninexnine_unit_6622(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E20N)
);

ninexnine_unit ninexnine_unit_6623(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F20N)
);

assign C320N=c3020N+c3120N+c3220N+c3320N+c3420N+c3520N+c3620N+c3720N+c3820N+c3920N+c3A20N+c3B20N+c3C20N+c3D20N+c3E20N+c3F20N;
assign A320N=(C320N>=0)?1:0;

assign P420N=A320N;

ninexnine_unit ninexnine_unit_6624(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3021N)
);

ninexnine_unit ninexnine_unit_6625(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3121N)
);

ninexnine_unit ninexnine_unit_6626(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3221N)
);

ninexnine_unit ninexnine_unit_6627(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3321N)
);

ninexnine_unit ninexnine_unit_6628(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3421N)
);

ninexnine_unit ninexnine_unit_6629(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3521N)
);

ninexnine_unit ninexnine_unit_6630(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3621N)
);

ninexnine_unit ninexnine_unit_6631(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3721N)
);

ninexnine_unit ninexnine_unit_6632(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3821N)
);

ninexnine_unit ninexnine_unit_6633(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3921N)
);

ninexnine_unit ninexnine_unit_6634(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A21N)
);

ninexnine_unit ninexnine_unit_6635(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B21N)
);

ninexnine_unit ninexnine_unit_6636(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C21N)
);

ninexnine_unit ninexnine_unit_6637(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D21N)
);

ninexnine_unit ninexnine_unit_6638(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E21N)
);

ninexnine_unit ninexnine_unit_6639(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F21N)
);

assign C321N=c3021N+c3121N+c3221N+c3321N+c3421N+c3521N+c3621N+c3721N+c3821N+c3921N+c3A21N+c3B21N+c3C21N+c3D21N+c3E21N+c3F21N;
assign A321N=(C321N>=0)?1:0;

assign P421N=A321N;

ninexnine_unit ninexnine_unit_6640(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3N000),
				.b1(W3N010),
				.b2(W3N020),
				.b3(W3N100),
				.b4(W3N110),
				.b5(W3N120),
				.b6(W3N200),
				.b7(W3N210),
				.b8(W3N220),
				.c(c3022N)
);

ninexnine_unit ninexnine_unit_6641(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3N001),
				.b1(W3N011),
				.b2(W3N021),
				.b3(W3N101),
				.b4(W3N111),
				.b5(W3N121),
				.b6(W3N201),
				.b7(W3N211),
				.b8(W3N221),
				.c(c3122N)
);

ninexnine_unit ninexnine_unit_6642(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3N002),
				.b1(W3N012),
				.b2(W3N022),
				.b3(W3N102),
				.b4(W3N112),
				.b5(W3N122),
				.b6(W3N202),
				.b7(W3N212),
				.b8(W3N222),
				.c(c3222N)
);

ninexnine_unit ninexnine_unit_6643(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3N003),
				.b1(W3N013),
				.b2(W3N023),
				.b3(W3N103),
				.b4(W3N113),
				.b5(W3N123),
				.b6(W3N203),
				.b7(W3N213),
				.b8(W3N223),
				.c(c3322N)
);

ninexnine_unit ninexnine_unit_6644(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3N004),
				.b1(W3N014),
				.b2(W3N024),
				.b3(W3N104),
				.b4(W3N114),
				.b5(W3N124),
				.b6(W3N204),
				.b7(W3N214),
				.b8(W3N224),
				.c(c3422N)
);

ninexnine_unit ninexnine_unit_6645(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3N005),
				.b1(W3N015),
				.b2(W3N025),
				.b3(W3N105),
				.b4(W3N115),
				.b5(W3N125),
				.b6(W3N205),
				.b7(W3N215),
				.b8(W3N225),
				.c(c3522N)
);

ninexnine_unit ninexnine_unit_6646(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3N006),
				.b1(W3N016),
				.b2(W3N026),
				.b3(W3N106),
				.b4(W3N116),
				.b5(W3N126),
				.b6(W3N206),
				.b7(W3N216),
				.b8(W3N226),
				.c(c3622N)
);

ninexnine_unit ninexnine_unit_6647(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3N007),
				.b1(W3N017),
				.b2(W3N027),
				.b3(W3N107),
				.b4(W3N117),
				.b5(W3N127),
				.b6(W3N207),
				.b7(W3N217),
				.b8(W3N227),
				.c(c3722N)
);

ninexnine_unit ninexnine_unit_6648(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3N008),
				.b1(W3N018),
				.b2(W3N028),
				.b3(W3N108),
				.b4(W3N118),
				.b5(W3N128),
				.b6(W3N208),
				.b7(W3N218),
				.b8(W3N228),
				.c(c3822N)
);

ninexnine_unit ninexnine_unit_6649(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3N009),
				.b1(W3N019),
				.b2(W3N029),
				.b3(W3N109),
				.b4(W3N119),
				.b5(W3N129),
				.b6(W3N209),
				.b7(W3N219),
				.b8(W3N229),
				.c(c3922N)
);

ninexnine_unit ninexnine_unit_6650(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3N00A),
				.b1(W3N01A),
				.b2(W3N02A),
				.b3(W3N10A),
				.b4(W3N11A),
				.b5(W3N12A),
				.b6(W3N20A),
				.b7(W3N21A),
				.b8(W3N22A),
				.c(c3A22N)
);

ninexnine_unit ninexnine_unit_6651(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3N00B),
				.b1(W3N01B),
				.b2(W3N02B),
				.b3(W3N10B),
				.b4(W3N11B),
				.b5(W3N12B),
				.b6(W3N20B),
				.b7(W3N21B),
				.b8(W3N22B),
				.c(c3B22N)
);

ninexnine_unit ninexnine_unit_6652(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3N00C),
				.b1(W3N01C),
				.b2(W3N02C),
				.b3(W3N10C),
				.b4(W3N11C),
				.b5(W3N12C),
				.b6(W3N20C),
				.b7(W3N21C),
				.b8(W3N22C),
				.c(c3C22N)
);

ninexnine_unit ninexnine_unit_6653(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3N00D),
				.b1(W3N01D),
				.b2(W3N02D),
				.b3(W3N10D),
				.b4(W3N11D),
				.b5(W3N12D),
				.b6(W3N20D),
				.b7(W3N21D),
				.b8(W3N22D),
				.c(c3D22N)
);

ninexnine_unit ninexnine_unit_6654(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3N00E),
				.b1(W3N01E),
				.b2(W3N02E),
				.b3(W3N10E),
				.b4(W3N11E),
				.b5(W3N12E),
				.b6(W3N20E),
				.b7(W3N21E),
				.b8(W3N22E),
				.c(c3E22N)
);

ninexnine_unit ninexnine_unit_6655(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3N00F),
				.b1(W3N01F),
				.b2(W3N02F),
				.b3(W3N10F),
				.b4(W3N11F),
				.b5(W3N12F),
				.b6(W3N20F),
				.b7(W3N21F),
				.b8(W3N22F),
				.c(c3F22N)
);

assign C322N=c3022N+c3122N+c3222N+c3322N+c3422N+c3522N+c3622N+c3722N+c3822N+c3922N+c3A22N+c3B22N+c3C22N+c3D22N+c3E22N+c3F22N;
assign A322N=(C322N>=0)?1:0;

assign P422N=A322N;

ninexnine_unit ninexnine_unit_6656(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3000O)
);

ninexnine_unit ninexnine_unit_6657(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3100O)
);

ninexnine_unit ninexnine_unit_6658(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3200O)
);

ninexnine_unit ninexnine_unit_6659(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3300O)
);

ninexnine_unit ninexnine_unit_6660(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3400O)
);

ninexnine_unit ninexnine_unit_6661(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3500O)
);

ninexnine_unit ninexnine_unit_6662(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3600O)
);

ninexnine_unit ninexnine_unit_6663(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3700O)
);

ninexnine_unit ninexnine_unit_6664(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3800O)
);

ninexnine_unit ninexnine_unit_6665(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3900O)
);

ninexnine_unit ninexnine_unit_6666(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A00O)
);

ninexnine_unit ninexnine_unit_6667(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B00O)
);

ninexnine_unit ninexnine_unit_6668(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C00O)
);

ninexnine_unit ninexnine_unit_6669(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D00O)
);

ninexnine_unit ninexnine_unit_6670(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E00O)
);

ninexnine_unit ninexnine_unit_6671(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F00O)
);

assign C300O=c3000O+c3100O+c3200O+c3300O+c3400O+c3500O+c3600O+c3700O+c3800O+c3900O+c3A00O+c3B00O+c3C00O+c3D00O+c3E00O+c3F00O;
assign A300O=(C300O>=0)?1:0;

assign P400O=A300O;

ninexnine_unit ninexnine_unit_6672(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3001O)
);

ninexnine_unit ninexnine_unit_6673(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3101O)
);

ninexnine_unit ninexnine_unit_6674(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3201O)
);

ninexnine_unit ninexnine_unit_6675(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3301O)
);

ninexnine_unit ninexnine_unit_6676(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3401O)
);

ninexnine_unit ninexnine_unit_6677(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3501O)
);

ninexnine_unit ninexnine_unit_6678(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3601O)
);

ninexnine_unit ninexnine_unit_6679(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3701O)
);

ninexnine_unit ninexnine_unit_6680(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3801O)
);

ninexnine_unit ninexnine_unit_6681(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3901O)
);

ninexnine_unit ninexnine_unit_6682(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A01O)
);

ninexnine_unit ninexnine_unit_6683(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B01O)
);

ninexnine_unit ninexnine_unit_6684(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C01O)
);

ninexnine_unit ninexnine_unit_6685(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D01O)
);

ninexnine_unit ninexnine_unit_6686(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E01O)
);

ninexnine_unit ninexnine_unit_6687(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F01O)
);

assign C301O=c3001O+c3101O+c3201O+c3301O+c3401O+c3501O+c3601O+c3701O+c3801O+c3901O+c3A01O+c3B01O+c3C01O+c3D01O+c3E01O+c3F01O;
assign A301O=(C301O>=0)?1:0;

assign P401O=A301O;

ninexnine_unit ninexnine_unit_6688(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3002O)
);

ninexnine_unit ninexnine_unit_6689(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3102O)
);

ninexnine_unit ninexnine_unit_6690(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3202O)
);

ninexnine_unit ninexnine_unit_6691(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3302O)
);

ninexnine_unit ninexnine_unit_6692(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3402O)
);

ninexnine_unit ninexnine_unit_6693(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3502O)
);

ninexnine_unit ninexnine_unit_6694(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3602O)
);

ninexnine_unit ninexnine_unit_6695(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3702O)
);

ninexnine_unit ninexnine_unit_6696(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3802O)
);

ninexnine_unit ninexnine_unit_6697(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3902O)
);

ninexnine_unit ninexnine_unit_6698(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A02O)
);

ninexnine_unit ninexnine_unit_6699(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B02O)
);

ninexnine_unit ninexnine_unit_6700(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C02O)
);

ninexnine_unit ninexnine_unit_6701(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D02O)
);

ninexnine_unit ninexnine_unit_6702(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E02O)
);

ninexnine_unit ninexnine_unit_6703(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F02O)
);

assign C302O=c3002O+c3102O+c3202O+c3302O+c3402O+c3502O+c3602O+c3702O+c3802O+c3902O+c3A02O+c3B02O+c3C02O+c3D02O+c3E02O+c3F02O;
assign A302O=(C302O>=0)?1:0;

assign P402O=A302O;

ninexnine_unit ninexnine_unit_6704(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3010O)
);

ninexnine_unit ninexnine_unit_6705(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3110O)
);

ninexnine_unit ninexnine_unit_6706(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3210O)
);

ninexnine_unit ninexnine_unit_6707(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3310O)
);

ninexnine_unit ninexnine_unit_6708(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3410O)
);

ninexnine_unit ninexnine_unit_6709(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3510O)
);

ninexnine_unit ninexnine_unit_6710(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3610O)
);

ninexnine_unit ninexnine_unit_6711(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3710O)
);

ninexnine_unit ninexnine_unit_6712(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3810O)
);

ninexnine_unit ninexnine_unit_6713(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3910O)
);

ninexnine_unit ninexnine_unit_6714(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A10O)
);

ninexnine_unit ninexnine_unit_6715(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B10O)
);

ninexnine_unit ninexnine_unit_6716(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C10O)
);

ninexnine_unit ninexnine_unit_6717(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D10O)
);

ninexnine_unit ninexnine_unit_6718(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E10O)
);

ninexnine_unit ninexnine_unit_6719(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F10O)
);

assign C310O=c3010O+c3110O+c3210O+c3310O+c3410O+c3510O+c3610O+c3710O+c3810O+c3910O+c3A10O+c3B10O+c3C10O+c3D10O+c3E10O+c3F10O;
assign A310O=(C310O>=0)?1:0;

assign P410O=A310O;

ninexnine_unit ninexnine_unit_6720(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3011O)
);

ninexnine_unit ninexnine_unit_6721(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3111O)
);

ninexnine_unit ninexnine_unit_6722(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3211O)
);

ninexnine_unit ninexnine_unit_6723(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3311O)
);

ninexnine_unit ninexnine_unit_6724(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3411O)
);

ninexnine_unit ninexnine_unit_6725(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3511O)
);

ninexnine_unit ninexnine_unit_6726(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3611O)
);

ninexnine_unit ninexnine_unit_6727(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3711O)
);

ninexnine_unit ninexnine_unit_6728(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3811O)
);

ninexnine_unit ninexnine_unit_6729(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3911O)
);

ninexnine_unit ninexnine_unit_6730(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A11O)
);

ninexnine_unit ninexnine_unit_6731(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B11O)
);

ninexnine_unit ninexnine_unit_6732(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C11O)
);

ninexnine_unit ninexnine_unit_6733(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D11O)
);

ninexnine_unit ninexnine_unit_6734(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E11O)
);

ninexnine_unit ninexnine_unit_6735(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F11O)
);

assign C311O=c3011O+c3111O+c3211O+c3311O+c3411O+c3511O+c3611O+c3711O+c3811O+c3911O+c3A11O+c3B11O+c3C11O+c3D11O+c3E11O+c3F11O;
assign A311O=(C311O>=0)?1:0;

assign P411O=A311O;

ninexnine_unit ninexnine_unit_6736(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3012O)
);

ninexnine_unit ninexnine_unit_6737(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3112O)
);

ninexnine_unit ninexnine_unit_6738(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3212O)
);

ninexnine_unit ninexnine_unit_6739(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3312O)
);

ninexnine_unit ninexnine_unit_6740(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3412O)
);

ninexnine_unit ninexnine_unit_6741(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3512O)
);

ninexnine_unit ninexnine_unit_6742(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3612O)
);

ninexnine_unit ninexnine_unit_6743(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3712O)
);

ninexnine_unit ninexnine_unit_6744(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3812O)
);

ninexnine_unit ninexnine_unit_6745(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3912O)
);

ninexnine_unit ninexnine_unit_6746(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A12O)
);

ninexnine_unit ninexnine_unit_6747(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B12O)
);

ninexnine_unit ninexnine_unit_6748(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C12O)
);

ninexnine_unit ninexnine_unit_6749(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D12O)
);

ninexnine_unit ninexnine_unit_6750(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E12O)
);

ninexnine_unit ninexnine_unit_6751(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F12O)
);

assign C312O=c3012O+c3112O+c3212O+c3312O+c3412O+c3512O+c3612O+c3712O+c3812O+c3912O+c3A12O+c3B12O+c3C12O+c3D12O+c3E12O+c3F12O;
assign A312O=(C312O>=0)?1:0;

assign P412O=A312O;

ninexnine_unit ninexnine_unit_6752(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3020O)
);

ninexnine_unit ninexnine_unit_6753(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3120O)
);

ninexnine_unit ninexnine_unit_6754(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3220O)
);

ninexnine_unit ninexnine_unit_6755(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3320O)
);

ninexnine_unit ninexnine_unit_6756(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3420O)
);

ninexnine_unit ninexnine_unit_6757(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3520O)
);

ninexnine_unit ninexnine_unit_6758(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3620O)
);

ninexnine_unit ninexnine_unit_6759(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3720O)
);

ninexnine_unit ninexnine_unit_6760(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3820O)
);

ninexnine_unit ninexnine_unit_6761(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3920O)
);

ninexnine_unit ninexnine_unit_6762(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A20O)
);

ninexnine_unit ninexnine_unit_6763(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B20O)
);

ninexnine_unit ninexnine_unit_6764(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C20O)
);

ninexnine_unit ninexnine_unit_6765(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D20O)
);

ninexnine_unit ninexnine_unit_6766(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E20O)
);

ninexnine_unit ninexnine_unit_6767(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F20O)
);

assign C320O=c3020O+c3120O+c3220O+c3320O+c3420O+c3520O+c3620O+c3720O+c3820O+c3920O+c3A20O+c3B20O+c3C20O+c3D20O+c3E20O+c3F20O;
assign A320O=(C320O>=0)?1:0;

assign P420O=A320O;

ninexnine_unit ninexnine_unit_6768(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3021O)
);

ninexnine_unit ninexnine_unit_6769(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3121O)
);

ninexnine_unit ninexnine_unit_6770(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3221O)
);

ninexnine_unit ninexnine_unit_6771(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3321O)
);

ninexnine_unit ninexnine_unit_6772(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3421O)
);

ninexnine_unit ninexnine_unit_6773(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3521O)
);

ninexnine_unit ninexnine_unit_6774(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3621O)
);

ninexnine_unit ninexnine_unit_6775(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3721O)
);

ninexnine_unit ninexnine_unit_6776(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3821O)
);

ninexnine_unit ninexnine_unit_6777(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3921O)
);

ninexnine_unit ninexnine_unit_6778(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A21O)
);

ninexnine_unit ninexnine_unit_6779(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B21O)
);

ninexnine_unit ninexnine_unit_6780(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C21O)
);

ninexnine_unit ninexnine_unit_6781(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D21O)
);

ninexnine_unit ninexnine_unit_6782(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E21O)
);

ninexnine_unit ninexnine_unit_6783(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F21O)
);

assign C321O=c3021O+c3121O+c3221O+c3321O+c3421O+c3521O+c3621O+c3721O+c3821O+c3921O+c3A21O+c3B21O+c3C21O+c3D21O+c3E21O+c3F21O;
assign A321O=(C321O>=0)?1:0;

assign P421O=A321O;

ninexnine_unit ninexnine_unit_6784(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3O000),
				.b1(W3O010),
				.b2(W3O020),
				.b3(W3O100),
				.b4(W3O110),
				.b5(W3O120),
				.b6(W3O200),
				.b7(W3O210),
				.b8(W3O220),
				.c(c3022O)
);

ninexnine_unit ninexnine_unit_6785(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3O001),
				.b1(W3O011),
				.b2(W3O021),
				.b3(W3O101),
				.b4(W3O111),
				.b5(W3O121),
				.b6(W3O201),
				.b7(W3O211),
				.b8(W3O221),
				.c(c3122O)
);

ninexnine_unit ninexnine_unit_6786(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3O002),
				.b1(W3O012),
				.b2(W3O022),
				.b3(W3O102),
				.b4(W3O112),
				.b5(W3O122),
				.b6(W3O202),
				.b7(W3O212),
				.b8(W3O222),
				.c(c3222O)
);

ninexnine_unit ninexnine_unit_6787(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3O003),
				.b1(W3O013),
				.b2(W3O023),
				.b3(W3O103),
				.b4(W3O113),
				.b5(W3O123),
				.b6(W3O203),
				.b7(W3O213),
				.b8(W3O223),
				.c(c3322O)
);

ninexnine_unit ninexnine_unit_6788(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3O004),
				.b1(W3O014),
				.b2(W3O024),
				.b3(W3O104),
				.b4(W3O114),
				.b5(W3O124),
				.b6(W3O204),
				.b7(W3O214),
				.b8(W3O224),
				.c(c3422O)
);

ninexnine_unit ninexnine_unit_6789(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3O005),
				.b1(W3O015),
				.b2(W3O025),
				.b3(W3O105),
				.b4(W3O115),
				.b5(W3O125),
				.b6(W3O205),
				.b7(W3O215),
				.b8(W3O225),
				.c(c3522O)
);

ninexnine_unit ninexnine_unit_6790(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3O006),
				.b1(W3O016),
				.b2(W3O026),
				.b3(W3O106),
				.b4(W3O116),
				.b5(W3O126),
				.b6(W3O206),
				.b7(W3O216),
				.b8(W3O226),
				.c(c3622O)
);

ninexnine_unit ninexnine_unit_6791(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3O007),
				.b1(W3O017),
				.b2(W3O027),
				.b3(W3O107),
				.b4(W3O117),
				.b5(W3O127),
				.b6(W3O207),
				.b7(W3O217),
				.b8(W3O227),
				.c(c3722O)
);

ninexnine_unit ninexnine_unit_6792(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3O008),
				.b1(W3O018),
				.b2(W3O028),
				.b3(W3O108),
				.b4(W3O118),
				.b5(W3O128),
				.b6(W3O208),
				.b7(W3O218),
				.b8(W3O228),
				.c(c3822O)
);

ninexnine_unit ninexnine_unit_6793(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3O009),
				.b1(W3O019),
				.b2(W3O029),
				.b3(W3O109),
				.b4(W3O119),
				.b5(W3O129),
				.b6(W3O209),
				.b7(W3O219),
				.b8(W3O229),
				.c(c3922O)
);

ninexnine_unit ninexnine_unit_6794(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3O00A),
				.b1(W3O01A),
				.b2(W3O02A),
				.b3(W3O10A),
				.b4(W3O11A),
				.b5(W3O12A),
				.b6(W3O20A),
				.b7(W3O21A),
				.b8(W3O22A),
				.c(c3A22O)
);

ninexnine_unit ninexnine_unit_6795(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3O00B),
				.b1(W3O01B),
				.b2(W3O02B),
				.b3(W3O10B),
				.b4(W3O11B),
				.b5(W3O12B),
				.b6(W3O20B),
				.b7(W3O21B),
				.b8(W3O22B),
				.c(c3B22O)
);

ninexnine_unit ninexnine_unit_6796(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3O00C),
				.b1(W3O01C),
				.b2(W3O02C),
				.b3(W3O10C),
				.b4(W3O11C),
				.b5(W3O12C),
				.b6(W3O20C),
				.b7(W3O21C),
				.b8(W3O22C),
				.c(c3C22O)
);

ninexnine_unit ninexnine_unit_6797(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3O00D),
				.b1(W3O01D),
				.b2(W3O02D),
				.b3(W3O10D),
				.b4(W3O11D),
				.b5(W3O12D),
				.b6(W3O20D),
				.b7(W3O21D),
				.b8(W3O22D),
				.c(c3D22O)
);

ninexnine_unit ninexnine_unit_6798(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3O00E),
				.b1(W3O01E),
				.b2(W3O02E),
				.b3(W3O10E),
				.b4(W3O11E),
				.b5(W3O12E),
				.b6(W3O20E),
				.b7(W3O21E),
				.b8(W3O22E),
				.c(c3E22O)
);

ninexnine_unit ninexnine_unit_6799(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3O00F),
				.b1(W3O01F),
				.b2(W3O02F),
				.b3(W3O10F),
				.b4(W3O11F),
				.b5(W3O12F),
				.b6(W3O20F),
				.b7(W3O21F),
				.b8(W3O22F),
				.c(c3F22O)
);

assign C322O=c3022O+c3122O+c3222O+c3322O+c3422O+c3522O+c3622O+c3722O+c3822O+c3922O+c3A22O+c3B22O+c3C22O+c3D22O+c3E22O+c3F22O;
assign A322O=(C322O>=0)?1:0;

assign P422O=A322O;

ninexnine_unit ninexnine_unit_6800(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3000P)
);

ninexnine_unit ninexnine_unit_6801(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3100P)
);

ninexnine_unit ninexnine_unit_6802(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3200P)
);

ninexnine_unit ninexnine_unit_6803(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3300P)
);

ninexnine_unit ninexnine_unit_6804(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3400P)
);

ninexnine_unit ninexnine_unit_6805(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3500P)
);

ninexnine_unit ninexnine_unit_6806(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3600P)
);

ninexnine_unit ninexnine_unit_6807(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3700P)
);

ninexnine_unit ninexnine_unit_6808(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3800P)
);

ninexnine_unit ninexnine_unit_6809(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3900P)
);

ninexnine_unit ninexnine_unit_6810(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A00P)
);

ninexnine_unit ninexnine_unit_6811(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B00P)
);

ninexnine_unit ninexnine_unit_6812(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C00P)
);

ninexnine_unit ninexnine_unit_6813(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D00P)
);

ninexnine_unit ninexnine_unit_6814(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E00P)
);

ninexnine_unit ninexnine_unit_6815(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F00P)
);

assign C300P=c3000P+c3100P+c3200P+c3300P+c3400P+c3500P+c3600P+c3700P+c3800P+c3900P+c3A00P+c3B00P+c3C00P+c3D00P+c3E00P+c3F00P;
assign A300P=(C300P>=0)?1:0;

assign P400P=A300P;

ninexnine_unit ninexnine_unit_6816(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3001P)
);

ninexnine_unit ninexnine_unit_6817(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3101P)
);

ninexnine_unit ninexnine_unit_6818(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3201P)
);

ninexnine_unit ninexnine_unit_6819(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3301P)
);

ninexnine_unit ninexnine_unit_6820(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3401P)
);

ninexnine_unit ninexnine_unit_6821(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3501P)
);

ninexnine_unit ninexnine_unit_6822(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3601P)
);

ninexnine_unit ninexnine_unit_6823(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3701P)
);

ninexnine_unit ninexnine_unit_6824(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3801P)
);

ninexnine_unit ninexnine_unit_6825(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3901P)
);

ninexnine_unit ninexnine_unit_6826(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A01P)
);

ninexnine_unit ninexnine_unit_6827(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B01P)
);

ninexnine_unit ninexnine_unit_6828(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C01P)
);

ninexnine_unit ninexnine_unit_6829(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D01P)
);

ninexnine_unit ninexnine_unit_6830(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E01P)
);

ninexnine_unit ninexnine_unit_6831(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F01P)
);

assign C301P=c3001P+c3101P+c3201P+c3301P+c3401P+c3501P+c3601P+c3701P+c3801P+c3901P+c3A01P+c3B01P+c3C01P+c3D01P+c3E01P+c3F01P;
assign A301P=(C301P>=0)?1:0;

assign P401P=A301P;

ninexnine_unit ninexnine_unit_6832(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3002P)
);

ninexnine_unit ninexnine_unit_6833(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3102P)
);

ninexnine_unit ninexnine_unit_6834(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3202P)
);

ninexnine_unit ninexnine_unit_6835(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3302P)
);

ninexnine_unit ninexnine_unit_6836(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3402P)
);

ninexnine_unit ninexnine_unit_6837(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3502P)
);

ninexnine_unit ninexnine_unit_6838(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3602P)
);

ninexnine_unit ninexnine_unit_6839(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3702P)
);

ninexnine_unit ninexnine_unit_6840(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3802P)
);

ninexnine_unit ninexnine_unit_6841(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3902P)
);

ninexnine_unit ninexnine_unit_6842(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A02P)
);

ninexnine_unit ninexnine_unit_6843(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B02P)
);

ninexnine_unit ninexnine_unit_6844(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C02P)
);

ninexnine_unit ninexnine_unit_6845(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D02P)
);

ninexnine_unit ninexnine_unit_6846(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E02P)
);

ninexnine_unit ninexnine_unit_6847(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F02P)
);

assign C302P=c3002P+c3102P+c3202P+c3302P+c3402P+c3502P+c3602P+c3702P+c3802P+c3902P+c3A02P+c3B02P+c3C02P+c3D02P+c3E02P+c3F02P;
assign A302P=(C302P>=0)?1:0;

assign P402P=A302P;

ninexnine_unit ninexnine_unit_6848(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3010P)
);

ninexnine_unit ninexnine_unit_6849(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3110P)
);

ninexnine_unit ninexnine_unit_6850(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3210P)
);

ninexnine_unit ninexnine_unit_6851(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3310P)
);

ninexnine_unit ninexnine_unit_6852(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3410P)
);

ninexnine_unit ninexnine_unit_6853(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3510P)
);

ninexnine_unit ninexnine_unit_6854(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3610P)
);

ninexnine_unit ninexnine_unit_6855(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3710P)
);

ninexnine_unit ninexnine_unit_6856(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3810P)
);

ninexnine_unit ninexnine_unit_6857(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3910P)
);

ninexnine_unit ninexnine_unit_6858(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A10P)
);

ninexnine_unit ninexnine_unit_6859(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B10P)
);

ninexnine_unit ninexnine_unit_6860(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C10P)
);

ninexnine_unit ninexnine_unit_6861(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D10P)
);

ninexnine_unit ninexnine_unit_6862(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E10P)
);

ninexnine_unit ninexnine_unit_6863(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F10P)
);

assign C310P=c3010P+c3110P+c3210P+c3310P+c3410P+c3510P+c3610P+c3710P+c3810P+c3910P+c3A10P+c3B10P+c3C10P+c3D10P+c3E10P+c3F10P;
assign A310P=(C310P>=0)?1:0;

assign P410P=A310P;

ninexnine_unit ninexnine_unit_6864(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3011P)
);

ninexnine_unit ninexnine_unit_6865(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3111P)
);

ninexnine_unit ninexnine_unit_6866(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3211P)
);

ninexnine_unit ninexnine_unit_6867(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3311P)
);

ninexnine_unit ninexnine_unit_6868(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3411P)
);

ninexnine_unit ninexnine_unit_6869(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3511P)
);

ninexnine_unit ninexnine_unit_6870(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3611P)
);

ninexnine_unit ninexnine_unit_6871(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3711P)
);

ninexnine_unit ninexnine_unit_6872(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3811P)
);

ninexnine_unit ninexnine_unit_6873(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3911P)
);

ninexnine_unit ninexnine_unit_6874(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A11P)
);

ninexnine_unit ninexnine_unit_6875(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B11P)
);

ninexnine_unit ninexnine_unit_6876(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C11P)
);

ninexnine_unit ninexnine_unit_6877(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D11P)
);

ninexnine_unit ninexnine_unit_6878(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E11P)
);

ninexnine_unit ninexnine_unit_6879(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F11P)
);

assign C311P=c3011P+c3111P+c3211P+c3311P+c3411P+c3511P+c3611P+c3711P+c3811P+c3911P+c3A11P+c3B11P+c3C11P+c3D11P+c3E11P+c3F11P;
assign A311P=(C311P>=0)?1:0;

assign P411P=A311P;

ninexnine_unit ninexnine_unit_6880(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3012P)
);

ninexnine_unit ninexnine_unit_6881(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3112P)
);

ninexnine_unit ninexnine_unit_6882(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3212P)
);

ninexnine_unit ninexnine_unit_6883(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3312P)
);

ninexnine_unit ninexnine_unit_6884(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3412P)
);

ninexnine_unit ninexnine_unit_6885(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3512P)
);

ninexnine_unit ninexnine_unit_6886(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3612P)
);

ninexnine_unit ninexnine_unit_6887(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3712P)
);

ninexnine_unit ninexnine_unit_6888(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3812P)
);

ninexnine_unit ninexnine_unit_6889(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3912P)
);

ninexnine_unit ninexnine_unit_6890(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A12P)
);

ninexnine_unit ninexnine_unit_6891(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B12P)
);

ninexnine_unit ninexnine_unit_6892(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C12P)
);

ninexnine_unit ninexnine_unit_6893(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D12P)
);

ninexnine_unit ninexnine_unit_6894(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E12P)
);

ninexnine_unit ninexnine_unit_6895(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F12P)
);

assign C312P=c3012P+c3112P+c3212P+c3312P+c3412P+c3512P+c3612P+c3712P+c3812P+c3912P+c3A12P+c3B12P+c3C12P+c3D12P+c3E12P+c3F12P;
assign A312P=(C312P>=0)?1:0;

assign P412P=A312P;

ninexnine_unit ninexnine_unit_6896(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3020P)
);

ninexnine_unit ninexnine_unit_6897(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3120P)
);

ninexnine_unit ninexnine_unit_6898(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3220P)
);

ninexnine_unit ninexnine_unit_6899(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3320P)
);

ninexnine_unit ninexnine_unit_6900(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3420P)
);

ninexnine_unit ninexnine_unit_6901(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3520P)
);

ninexnine_unit ninexnine_unit_6902(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3620P)
);

ninexnine_unit ninexnine_unit_6903(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3720P)
);

ninexnine_unit ninexnine_unit_6904(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3820P)
);

ninexnine_unit ninexnine_unit_6905(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3920P)
);

ninexnine_unit ninexnine_unit_6906(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A20P)
);

ninexnine_unit ninexnine_unit_6907(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B20P)
);

ninexnine_unit ninexnine_unit_6908(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C20P)
);

ninexnine_unit ninexnine_unit_6909(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D20P)
);

ninexnine_unit ninexnine_unit_6910(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E20P)
);

ninexnine_unit ninexnine_unit_6911(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F20P)
);

assign C320P=c3020P+c3120P+c3220P+c3320P+c3420P+c3520P+c3620P+c3720P+c3820P+c3920P+c3A20P+c3B20P+c3C20P+c3D20P+c3E20P+c3F20P;
assign A320P=(C320P>=0)?1:0;

assign P420P=A320P;

ninexnine_unit ninexnine_unit_6912(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3021P)
);

ninexnine_unit ninexnine_unit_6913(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3121P)
);

ninexnine_unit ninexnine_unit_6914(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3221P)
);

ninexnine_unit ninexnine_unit_6915(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3321P)
);

ninexnine_unit ninexnine_unit_6916(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3421P)
);

ninexnine_unit ninexnine_unit_6917(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3521P)
);

ninexnine_unit ninexnine_unit_6918(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3621P)
);

ninexnine_unit ninexnine_unit_6919(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3721P)
);

ninexnine_unit ninexnine_unit_6920(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3821P)
);

ninexnine_unit ninexnine_unit_6921(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3921P)
);

ninexnine_unit ninexnine_unit_6922(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A21P)
);

ninexnine_unit ninexnine_unit_6923(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B21P)
);

ninexnine_unit ninexnine_unit_6924(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C21P)
);

ninexnine_unit ninexnine_unit_6925(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D21P)
);

ninexnine_unit ninexnine_unit_6926(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E21P)
);

ninexnine_unit ninexnine_unit_6927(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F21P)
);

assign C321P=c3021P+c3121P+c3221P+c3321P+c3421P+c3521P+c3621P+c3721P+c3821P+c3921P+c3A21P+c3B21P+c3C21P+c3D21P+c3E21P+c3F21P;
assign A321P=(C321P>=0)?1:0;

assign P421P=A321P;

ninexnine_unit ninexnine_unit_6928(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3P000),
				.b1(W3P010),
				.b2(W3P020),
				.b3(W3P100),
				.b4(W3P110),
				.b5(W3P120),
				.b6(W3P200),
				.b7(W3P210),
				.b8(W3P220),
				.c(c3022P)
);

ninexnine_unit ninexnine_unit_6929(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3P001),
				.b1(W3P011),
				.b2(W3P021),
				.b3(W3P101),
				.b4(W3P111),
				.b5(W3P121),
				.b6(W3P201),
				.b7(W3P211),
				.b8(W3P221),
				.c(c3122P)
);

ninexnine_unit ninexnine_unit_6930(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3P002),
				.b1(W3P012),
				.b2(W3P022),
				.b3(W3P102),
				.b4(W3P112),
				.b5(W3P122),
				.b6(W3P202),
				.b7(W3P212),
				.b8(W3P222),
				.c(c3222P)
);

ninexnine_unit ninexnine_unit_6931(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3P003),
				.b1(W3P013),
				.b2(W3P023),
				.b3(W3P103),
				.b4(W3P113),
				.b5(W3P123),
				.b6(W3P203),
				.b7(W3P213),
				.b8(W3P223),
				.c(c3322P)
);

ninexnine_unit ninexnine_unit_6932(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3P004),
				.b1(W3P014),
				.b2(W3P024),
				.b3(W3P104),
				.b4(W3P114),
				.b5(W3P124),
				.b6(W3P204),
				.b7(W3P214),
				.b8(W3P224),
				.c(c3422P)
);

ninexnine_unit ninexnine_unit_6933(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3P005),
				.b1(W3P015),
				.b2(W3P025),
				.b3(W3P105),
				.b4(W3P115),
				.b5(W3P125),
				.b6(W3P205),
				.b7(W3P215),
				.b8(W3P225),
				.c(c3522P)
);

ninexnine_unit ninexnine_unit_6934(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3P006),
				.b1(W3P016),
				.b2(W3P026),
				.b3(W3P106),
				.b4(W3P116),
				.b5(W3P126),
				.b6(W3P206),
				.b7(W3P216),
				.b8(W3P226),
				.c(c3622P)
);

ninexnine_unit ninexnine_unit_6935(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3P007),
				.b1(W3P017),
				.b2(W3P027),
				.b3(W3P107),
				.b4(W3P117),
				.b5(W3P127),
				.b6(W3P207),
				.b7(W3P217),
				.b8(W3P227),
				.c(c3722P)
);

ninexnine_unit ninexnine_unit_6936(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3P008),
				.b1(W3P018),
				.b2(W3P028),
				.b3(W3P108),
				.b4(W3P118),
				.b5(W3P128),
				.b6(W3P208),
				.b7(W3P218),
				.b8(W3P228),
				.c(c3822P)
);

ninexnine_unit ninexnine_unit_6937(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3P009),
				.b1(W3P019),
				.b2(W3P029),
				.b3(W3P109),
				.b4(W3P119),
				.b5(W3P129),
				.b6(W3P209),
				.b7(W3P219),
				.b8(W3P229),
				.c(c3922P)
);

ninexnine_unit ninexnine_unit_6938(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3P00A),
				.b1(W3P01A),
				.b2(W3P02A),
				.b3(W3P10A),
				.b4(W3P11A),
				.b5(W3P12A),
				.b6(W3P20A),
				.b7(W3P21A),
				.b8(W3P22A),
				.c(c3A22P)
);

ninexnine_unit ninexnine_unit_6939(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3P00B),
				.b1(W3P01B),
				.b2(W3P02B),
				.b3(W3P10B),
				.b4(W3P11B),
				.b5(W3P12B),
				.b6(W3P20B),
				.b7(W3P21B),
				.b8(W3P22B),
				.c(c3B22P)
);

ninexnine_unit ninexnine_unit_6940(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3P00C),
				.b1(W3P01C),
				.b2(W3P02C),
				.b3(W3P10C),
				.b4(W3P11C),
				.b5(W3P12C),
				.b6(W3P20C),
				.b7(W3P21C),
				.b8(W3P22C),
				.c(c3C22P)
);

ninexnine_unit ninexnine_unit_6941(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3P00D),
				.b1(W3P01D),
				.b2(W3P02D),
				.b3(W3P10D),
				.b4(W3P11D),
				.b5(W3P12D),
				.b6(W3P20D),
				.b7(W3P21D),
				.b8(W3P22D),
				.c(c3D22P)
);

ninexnine_unit ninexnine_unit_6942(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3P00E),
				.b1(W3P01E),
				.b2(W3P02E),
				.b3(W3P10E),
				.b4(W3P11E),
				.b5(W3P12E),
				.b6(W3P20E),
				.b7(W3P21E),
				.b8(W3P22E),
				.c(c3E22P)
);

ninexnine_unit ninexnine_unit_6943(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3P00F),
				.b1(W3P01F),
				.b2(W3P02F),
				.b3(W3P10F),
				.b4(W3P11F),
				.b5(W3P12F),
				.b6(W3P20F),
				.b7(W3P21F),
				.b8(W3P22F),
				.c(c3F22P)
);

assign C322P=c3022P+c3122P+c3222P+c3322P+c3422P+c3522P+c3622P+c3722P+c3822P+c3922P+c3A22P+c3B22P+c3C22P+c3D22P+c3E22P+c3F22P;
assign A322P=(C322P>=0)?1:0;

assign P422P=A322P;

ninexnine_unit ninexnine_unit_6944(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3000Q)
);

ninexnine_unit ninexnine_unit_6945(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3100Q)
);

ninexnine_unit ninexnine_unit_6946(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3200Q)
);

ninexnine_unit ninexnine_unit_6947(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3300Q)
);

ninexnine_unit ninexnine_unit_6948(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3400Q)
);

ninexnine_unit ninexnine_unit_6949(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3500Q)
);

ninexnine_unit ninexnine_unit_6950(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3600Q)
);

ninexnine_unit ninexnine_unit_6951(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3700Q)
);

ninexnine_unit ninexnine_unit_6952(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3800Q)
);

ninexnine_unit ninexnine_unit_6953(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3900Q)
);

ninexnine_unit ninexnine_unit_6954(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A00Q)
);

ninexnine_unit ninexnine_unit_6955(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B00Q)
);

ninexnine_unit ninexnine_unit_6956(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C00Q)
);

ninexnine_unit ninexnine_unit_6957(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D00Q)
);

ninexnine_unit ninexnine_unit_6958(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E00Q)
);

ninexnine_unit ninexnine_unit_6959(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F00Q)
);

assign C300Q=c3000Q+c3100Q+c3200Q+c3300Q+c3400Q+c3500Q+c3600Q+c3700Q+c3800Q+c3900Q+c3A00Q+c3B00Q+c3C00Q+c3D00Q+c3E00Q+c3F00Q;
assign A300Q=(C300Q>=0)?1:0;

assign P400Q=A300Q;

ninexnine_unit ninexnine_unit_6960(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3001Q)
);

ninexnine_unit ninexnine_unit_6961(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3101Q)
);

ninexnine_unit ninexnine_unit_6962(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3201Q)
);

ninexnine_unit ninexnine_unit_6963(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3301Q)
);

ninexnine_unit ninexnine_unit_6964(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3401Q)
);

ninexnine_unit ninexnine_unit_6965(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3501Q)
);

ninexnine_unit ninexnine_unit_6966(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3601Q)
);

ninexnine_unit ninexnine_unit_6967(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3701Q)
);

ninexnine_unit ninexnine_unit_6968(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3801Q)
);

ninexnine_unit ninexnine_unit_6969(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3901Q)
);

ninexnine_unit ninexnine_unit_6970(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A01Q)
);

ninexnine_unit ninexnine_unit_6971(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B01Q)
);

ninexnine_unit ninexnine_unit_6972(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C01Q)
);

ninexnine_unit ninexnine_unit_6973(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D01Q)
);

ninexnine_unit ninexnine_unit_6974(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E01Q)
);

ninexnine_unit ninexnine_unit_6975(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F01Q)
);

assign C301Q=c3001Q+c3101Q+c3201Q+c3301Q+c3401Q+c3501Q+c3601Q+c3701Q+c3801Q+c3901Q+c3A01Q+c3B01Q+c3C01Q+c3D01Q+c3E01Q+c3F01Q;
assign A301Q=(C301Q>=0)?1:0;

assign P401Q=A301Q;

ninexnine_unit ninexnine_unit_6976(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3002Q)
);

ninexnine_unit ninexnine_unit_6977(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3102Q)
);

ninexnine_unit ninexnine_unit_6978(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3202Q)
);

ninexnine_unit ninexnine_unit_6979(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3302Q)
);

ninexnine_unit ninexnine_unit_6980(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3402Q)
);

ninexnine_unit ninexnine_unit_6981(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3502Q)
);

ninexnine_unit ninexnine_unit_6982(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3602Q)
);

ninexnine_unit ninexnine_unit_6983(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3702Q)
);

ninexnine_unit ninexnine_unit_6984(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3802Q)
);

ninexnine_unit ninexnine_unit_6985(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3902Q)
);

ninexnine_unit ninexnine_unit_6986(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A02Q)
);

ninexnine_unit ninexnine_unit_6987(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B02Q)
);

ninexnine_unit ninexnine_unit_6988(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C02Q)
);

ninexnine_unit ninexnine_unit_6989(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D02Q)
);

ninexnine_unit ninexnine_unit_6990(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E02Q)
);

ninexnine_unit ninexnine_unit_6991(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F02Q)
);

assign C302Q=c3002Q+c3102Q+c3202Q+c3302Q+c3402Q+c3502Q+c3602Q+c3702Q+c3802Q+c3902Q+c3A02Q+c3B02Q+c3C02Q+c3D02Q+c3E02Q+c3F02Q;
assign A302Q=(C302Q>=0)?1:0;

assign P402Q=A302Q;

ninexnine_unit ninexnine_unit_6992(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3010Q)
);

ninexnine_unit ninexnine_unit_6993(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3110Q)
);

ninexnine_unit ninexnine_unit_6994(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3210Q)
);

ninexnine_unit ninexnine_unit_6995(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3310Q)
);

ninexnine_unit ninexnine_unit_6996(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3410Q)
);

ninexnine_unit ninexnine_unit_6997(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3510Q)
);

ninexnine_unit ninexnine_unit_6998(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3610Q)
);

ninexnine_unit ninexnine_unit_6999(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3710Q)
);

ninexnine_unit ninexnine_unit_7000(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3810Q)
);

ninexnine_unit ninexnine_unit_7001(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3910Q)
);

ninexnine_unit ninexnine_unit_7002(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A10Q)
);

ninexnine_unit ninexnine_unit_7003(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B10Q)
);

ninexnine_unit ninexnine_unit_7004(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C10Q)
);

ninexnine_unit ninexnine_unit_7005(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D10Q)
);

ninexnine_unit ninexnine_unit_7006(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E10Q)
);

ninexnine_unit ninexnine_unit_7007(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F10Q)
);

assign C310Q=c3010Q+c3110Q+c3210Q+c3310Q+c3410Q+c3510Q+c3610Q+c3710Q+c3810Q+c3910Q+c3A10Q+c3B10Q+c3C10Q+c3D10Q+c3E10Q+c3F10Q;
assign A310Q=(C310Q>=0)?1:0;

assign P410Q=A310Q;

ninexnine_unit ninexnine_unit_7008(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3011Q)
);

ninexnine_unit ninexnine_unit_7009(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3111Q)
);

ninexnine_unit ninexnine_unit_7010(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3211Q)
);

ninexnine_unit ninexnine_unit_7011(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3311Q)
);

ninexnine_unit ninexnine_unit_7012(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3411Q)
);

ninexnine_unit ninexnine_unit_7013(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3511Q)
);

ninexnine_unit ninexnine_unit_7014(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3611Q)
);

ninexnine_unit ninexnine_unit_7015(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3711Q)
);

ninexnine_unit ninexnine_unit_7016(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3811Q)
);

ninexnine_unit ninexnine_unit_7017(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3911Q)
);

ninexnine_unit ninexnine_unit_7018(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A11Q)
);

ninexnine_unit ninexnine_unit_7019(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B11Q)
);

ninexnine_unit ninexnine_unit_7020(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C11Q)
);

ninexnine_unit ninexnine_unit_7021(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D11Q)
);

ninexnine_unit ninexnine_unit_7022(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E11Q)
);

ninexnine_unit ninexnine_unit_7023(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F11Q)
);

assign C311Q=c3011Q+c3111Q+c3211Q+c3311Q+c3411Q+c3511Q+c3611Q+c3711Q+c3811Q+c3911Q+c3A11Q+c3B11Q+c3C11Q+c3D11Q+c3E11Q+c3F11Q;
assign A311Q=(C311Q>=0)?1:0;

assign P411Q=A311Q;

ninexnine_unit ninexnine_unit_7024(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3012Q)
);

ninexnine_unit ninexnine_unit_7025(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3112Q)
);

ninexnine_unit ninexnine_unit_7026(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3212Q)
);

ninexnine_unit ninexnine_unit_7027(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3312Q)
);

ninexnine_unit ninexnine_unit_7028(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3412Q)
);

ninexnine_unit ninexnine_unit_7029(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3512Q)
);

ninexnine_unit ninexnine_unit_7030(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3612Q)
);

ninexnine_unit ninexnine_unit_7031(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3712Q)
);

ninexnine_unit ninexnine_unit_7032(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3812Q)
);

ninexnine_unit ninexnine_unit_7033(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3912Q)
);

ninexnine_unit ninexnine_unit_7034(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A12Q)
);

ninexnine_unit ninexnine_unit_7035(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B12Q)
);

ninexnine_unit ninexnine_unit_7036(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C12Q)
);

ninexnine_unit ninexnine_unit_7037(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D12Q)
);

ninexnine_unit ninexnine_unit_7038(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E12Q)
);

ninexnine_unit ninexnine_unit_7039(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F12Q)
);

assign C312Q=c3012Q+c3112Q+c3212Q+c3312Q+c3412Q+c3512Q+c3612Q+c3712Q+c3812Q+c3912Q+c3A12Q+c3B12Q+c3C12Q+c3D12Q+c3E12Q+c3F12Q;
assign A312Q=(C312Q>=0)?1:0;

assign P412Q=A312Q;

ninexnine_unit ninexnine_unit_7040(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3020Q)
);

ninexnine_unit ninexnine_unit_7041(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3120Q)
);

ninexnine_unit ninexnine_unit_7042(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3220Q)
);

ninexnine_unit ninexnine_unit_7043(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3320Q)
);

ninexnine_unit ninexnine_unit_7044(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3420Q)
);

ninexnine_unit ninexnine_unit_7045(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3520Q)
);

ninexnine_unit ninexnine_unit_7046(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3620Q)
);

ninexnine_unit ninexnine_unit_7047(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3720Q)
);

ninexnine_unit ninexnine_unit_7048(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3820Q)
);

ninexnine_unit ninexnine_unit_7049(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3920Q)
);

ninexnine_unit ninexnine_unit_7050(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A20Q)
);

ninexnine_unit ninexnine_unit_7051(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B20Q)
);

ninexnine_unit ninexnine_unit_7052(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C20Q)
);

ninexnine_unit ninexnine_unit_7053(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D20Q)
);

ninexnine_unit ninexnine_unit_7054(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E20Q)
);

ninexnine_unit ninexnine_unit_7055(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F20Q)
);

assign C320Q=c3020Q+c3120Q+c3220Q+c3320Q+c3420Q+c3520Q+c3620Q+c3720Q+c3820Q+c3920Q+c3A20Q+c3B20Q+c3C20Q+c3D20Q+c3E20Q+c3F20Q;
assign A320Q=(C320Q>=0)?1:0;

assign P420Q=A320Q;

ninexnine_unit ninexnine_unit_7056(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3021Q)
);

ninexnine_unit ninexnine_unit_7057(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3121Q)
);

ninexnine_unit ninexnine_unit_7058(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3221Q)
);

ninexnine_unit ninexnine_unit_7059(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3321Q)
);

ninexnine_unit ninexnine_unit_7060(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3421Q)
);

ninexnine_unit ninexnine_unit_7061(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3521Q)
);

ninexnine_unit ninexnine_unit_7062(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3621Q)
);

ninexnine_unit ninexnine_unit_7063(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3721Q)
);

ninexnine_unit ninexnine_unit_7064(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3821Q)
);

ninexnine_unit ninexnine_unit_7065(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3921Q)
);

ninexnine_unit ninexnine_unit_7066(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A21Q)
);

ninexnine_unit ninexnine_unit_7067(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B21Q)
);

ninexnine_unit ninexnine_unit_7068(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C21Q)
);

ninexnine_unit ninexnine_unit_7069(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D21Q)
);

ninexnine_unit ninexnine_unit_7070(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E21Q)
);

ninexnine_unit ninexnine_unit_7071(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F21Q)
);

assign C321Q=c3021Q+c3121Q+c3221Q+c3321Q+c3421Q+c3521Q+c3621Q+c3721Q+c3821Q+c3921Q+c3A21Q+c3B21Q+c3C21Q+c3D21Q+c3E21Q+c3F21Q;
assign A321Q=(C321Q>=0)?1:0;

assign P421Q=A321Q;

ninexnine_unit ninexnine_unit_7072(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3Q000),
				.b1(W3Q010),
				.b2(W3Q020),
				.b3(W3Q100),
				.b4(W3Q110),
				.b5(W3Q120),
				.b6(W3Q200),
				.b7(W3Q210),
				.b8(W3Q220),
				.c(c3022Q)
);

ninexnine_unit ninexnine_unit_7073(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3Q001),
				.b1(W3Q011),
				.b2(W3Q021),
				.b3(W3Q101),
				.b4(W3Q111),
				.b5(W3Q121),
				.b6(W3Q201),
				.b7(W3Q211),
				.b8(W3Q221),
				.c(c3122Q)
);

ninexnine_unit ninexnine_unit_7074(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3Q002),
				.b1(W3Q012),
				.b2(W3Q022),
				.b3(W3Q102),
				.b4(W3Q112),
				.b5(W3Q122),
				.b6(W3Q202),
				.b7(W3Q212),
				.b8(W3Q222),
				.c(c3222Q)
);

ninexnine_unit ninexnine_unit_7075(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3Q003),
				.b1(W3Q013),
				.b2(W3Q023),
				.b3(W3Q103),
				.b4(W3Q113),
				.b5(W3Q123),
				.b6(W3Q203),
				.b7(W3Q213),
				.b8(W3Q223),
				.c(c3322Q)
);

ninexnine_unit ninexnine_unit_7076(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3Q004),
				.b1(W3Q014),
				.b2(W3Q024),
				.b3(W3Q104),
				.b4(W3Q114),
				.b5(W3Q124),
				.b6(W3Q204),
				.b7(W3Q214),
				.b8(W3Q224),
				.c(c3422Q)
);

ninexnine_unit ninexnine_unit_7077(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3Q005),
				.b1(W3Q015),
				.b2(W3Q025),
				.b3(W3Q105),
				.b4(W3Q115),
				.b5(W3Q125),
				.b6(W3Q205),
				.b7(W3Q215),
				.b8(W3Q225),
				.c(c3522Q)
);

ninexnine_unit ninexnine_unit_7078(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3Q006),
				.b1(W3Q016),
				.b2(W3Q026),
				.b3(W3Q106),
				.b4(W3Q116),
				.b5(W3Q126),
				.b6(W3Q206),
				.b7(W3Q216),
				.b8(W3Q226),
				.c(c3622Q)
);

ninexnine_unit ninexnine_unit_7079(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3Q007),
				.b1(W3Q017),
				.b2(W3Q027),
				.b3(W3Q107),
				.b4(W3Q117),
				.b5(W3Q127),
				.b6(W3Q207),
				.b7(W3Q217),
				.b8(W3Q227),
				.c(c3722Q)
);

ninexnine_unit ninexnine_unit_7080(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3Q008),
				.b1(W3Q018),
				.b2(W3Q028),
				.b3(W3Q108),
				.b4(W3Q118),
				.b5(W3Q128),
				.b6(W3Q208),
				.b7(W3Q218),
				.b8(W3Q228),
				.c(c3822Q)
);

ninexnine_unit ninexnine_unit_7081(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3Q009),
				.b1(W3Q019),
				.b2(W3Q029),
				.b3(W3Q109),
				.b4(W3Q119),
				.b5(W3Q129),
				.b6(W3Q209),
				.b7(W3Q219),
				.b8(W3Q229),
				.c(c3922Q)
);

ninexnine_unit ninexnine_unit_7082(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3Q00A),
				.b1(W3Q01A),
				.b2(W3Q02A),
				.b3(W3Q10A),
				.b4(W3Q11A),
				.b5(W3Q12A),
				.b6(W3Q20A),
				.b7(W3Q21A),
				.b8(W3Q22A),
				.c(c3A22Q)
);

ninexnine_unit ninexnine_unit_7083(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3Q00B),
				.b1(W3Q01B),
				.b2(W3Q02B),
				.b3(W3Q10B),
				.b4(W3Q11B),
				.b5(W3Q12B),
				.b6(W3Q20B),
				.b7(W3Q21B),
				.b8(W3Q22B),
				.c(c3B22Q)
);

ninexnine_unit ninexnine_unit_7084(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3Q00C),
				.b1(W3Q01C),
				.b2(W3Q02C),
				.b3(W3Q10C),
				.b4(W3Q11C),
				.b5(W3Q12C),
				.b6(W3Q20C),
				.b7(W3Q21C),
				.b8(W3Q22C),
				.c(c3C22Q)
);

ninexnine_unit ninexnine_unit_7085(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3Q00D),
				.b1(W3Q01D),
				.b2(W3Q02D),
				.b3(W3Q10D),
				.b4(W3Q11D),
				.b5(W3Q12D),
				.b6(W3Q20D),
				.b7(W3Q21D),
				.b8(W3Q22D),
				.c(c3D22Q)
);

ninexnine_unit ninexnine_unit_7086(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3Q00E),
				.b1(W3Q01E),
				.b2(W3Q02E),
				.b3(W3Q10E),
				.b4(W3Q11E),
				.b5(W3Q12E),
				.b6(W3Q20E),
				.b7(W3Q21E),
				.b8(W3Q22E),
				.c(c3E22Q)
);

ninexnine_unit ninexnine_unit_7087(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3Q00F),
				.b1(W3Q01F),
				.b2(W3Q02F),
				.b3(W3Q10F),
				.b4(W3Q11F),
				.b5(W3Q12F),
				.b6(W3Q20F),
				.b7(W3Q21F),
				.b8(W3Q22F),
				.c(c3F22Q)
);

assign C322Q=c3022Q+c3122Q+c3222Q+c3322Q+c3422Q+c3522Q+c3622Q+c3722Q+c3822Q+c3922Q+c3A22Q+c3B22Q+c3C22Q+c3D22Q+c3E22Q+c3F22Q;
assign A322Q=(C322Q>=0)?1:0;

assign P422Q=A322Q;

ninexnine_unit ninexnine_unit_7088(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3000R)
);

ninexnine_unit ninexnine_unit_7089(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3100R)
);

ninexnine_unit ninexnine_unit_7090(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3200R)
);

ninexnine_unit ninexnine_unit_7091(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3300R)
);

ninexnine_unit ninexnine_unit_7092(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3400R)
);

ninexnine_unit ninexnine_unit_7093(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3500R)
);

ninexnine_unit ninexnine_unit_7094(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3600R)
);

ninexnine_unit ninexnine_unit_7095(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3700R)
);

ninexnine_unit ninexnine_unit_7096(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3800R)
);

ninexnine_unit ninexnine_unit_7097(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3900R)
);

ninexnine_unit ninexnine_unit_7098(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A00R)
);

ninexnine_unit ninexnine_unit_7099(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B00R)
);

ninexnine_unit ninexnine_unit_7100(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C00R)
);

ninexnine_unit ninexnine_unit_7101(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D00R)
);

ninexnine_unit ninexnine_unit_7102(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E00R)
);

ninexnine_unit ninexnine_unit_7103(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F00R)
);

assign C300R=c3000R+c3100R+c3200R+c3300R+c3400R+c3500R+c3600R+c3700R+c3800R+c3900R+c3A00R+c3B00R+c3C00R+c3D00R+c3E00R+c3F00R;
assign A300R=(C300R>=0)?1:0;

assign P400R=A300R;

ninexnine_unit ninexnine_unit_7104(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3001R)
);

ninexnine_unit ninexnine_unit_7105(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3101R)
);

ninexnine_unit ninexnine_unit_7106(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3201R)
);

ninexnine_unit ninexnine_unit_7107(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3301R)
);

ninexnine_unit ninexnine_unit_7108(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3401R)
);

ninexnine_unit ninexnine_unit_7109(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3501R)
);

ninexnine_unit ninexnine_unit_7110(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3601R)
);

ninexnine_unit ninexnine_unit_7111(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3701R)
);

ninexnine_unit ninexnine_unit_7112(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3801R)
);

ninexnine_unit ninexnine_unit_7113(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3901R)
);

ninexnine_unit ninexnine_unit_7114(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A01R)
);

ninexnine_unit ninexnine_unit_7115(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B01R)
);

ninexnine_unit ninexnine_unit_7116(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C01R)
);

ninexnine_unit ninexnine_unit_7117(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D01R)
);

ninexnine_unit ninexnine_unit_7118(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E01R)
);

ninexnine_unit ninexnine_unit_7119(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F01R)
);

assign C301R=c3001R+c3101R+c3201R+c3301R+c3401R+c3501R+c3601R+c3701R+c3801R+c3901R+c3A01R+c3B01R+c3C01R+c3D01R+c3E01R+c3F01R;
assign A301R=(C301R>=0)?1:0;

assign P401R=A301R;

ninexnine_unit ninexnine_unit_7120(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3002R)
);

ninexnine_unit ninexnine_unit_7121(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3102R)
);

ninexnine_unit ninexnine_unit_7122(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3202R)
);

ninexnine_unit ninexnine_unit_7123(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3302R)
);

ninexnine_unit ninexnine_unit_7124(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3402R)
);

ninexnine_unit ninexnine_unit_7125(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3502R)
);

ninexnine_unit ninexnine_unit_7126(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3602R)
);

ninexnine_unit ninexnine_unit_7127(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3702R)
);

ninexnine_unit ninexnine_unit_7128(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3802R)
);

ninexnine_unit ninexnine_unit_7129(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3902R)
);

ninexnine_unit ninexnine_unit_7130(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A02R)
);

ninexnine_unit ninexnine_unit_7131(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B02R)
);

ninexnine_unit ninexnine_unit_7132(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C02R)
);

ninexnine_unit ninexnine_unit_7133(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D02R)
);

ninexnine_unit ninexnine_unit_7134(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E02R)
);

ninexnine_unit ninexnine_unit_7135(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F02R)
);

assign C302R=c3002R+c3102R+c3202R+c3302R+c3402R+c3502R+c3602R+c3702R+c3802R+c3902R+c3A02R+c3B02R+c3C02R+c3D02R+c3E02R+c3F02R;
assign A302R=(C302R>=0)?1:0;

assign P402R=A302R;

ninexnine_unit ninexnine_unit_7136(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3010R)
);

ninexnine_unit ninexnine_unit_7137(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3110R)
);

ninexnine_unit ninexnine_unit_7138(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3210R)
);

ninexnine_unit ninexnine_unit_7139(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3310R)
);

ninexnine_unit ninexnine_unit_7140(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3410R)
);

ninexnine_unit ninexnine_unit_7141(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3510R)
);

ninexnine_unit ninexnine_unit_7142(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3610R)
);

ninexnine_unit ninexnine_unit_7143(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3710R)
);

ninexnine_unit ninexnine_unit_7144(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3810R)
);

ninexnine_unit ninexnine_unit_7145(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3910R)
);

ninexnine_unit ninexnine_unit_7146(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A10R)
);

ninexnine_unit ninexnine_unit_7147(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B10R)
);

ninexnine_unit ninexnine_unit_7148(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C10R)
);

ninexnine_unit ninexnine_unit_7149(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D10R)
);

ninexnine_unit ninexnine_unit_7150(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E10R)
);

ninexnine_unit ninexnine_unit_7151(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F10R)
);

assign C310R=c3010R+c3110R+c3210R+c3310R+c3410R+c3510R+c3610R+c3710R+c3810R+c3910R+c3A10R+c3B10R+c3C10R+c3D10R+c3E10R+c3F10R;
assign A310R=(C310R>=0)?1:0;

assign P410R=A310R;

ninexnine_unit ninexnine_unit_7152(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3011R)
);

ninexnine_unit ninexnine_unit_7153(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3111R)
);

ninexnine_unit ninexnine_unit_7154(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3211R)
);

ninexnine_unit ninexnine_unit_7155(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3311R)
);

ninexnine_unit ninexnine_unit_7156(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3411R)
);

ninexnine_unit ninexnine_unit_7157(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3511R)
);

ninexnine_unit ninexnine_unit_7158(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3611R)
);

ninexnine_unit ninexnine_unit_7159(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3711R)
);

ninexnine_unit ninexnine_unit_7160(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3811R)
);

ninexnine_unit ninexnine_unit_7161(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3911R)
);

ninexnine_unit ninexnine_unit_7162(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A11R)
);

ninexnine_unit ninexnine_unit_7163(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B11R)
);

ninexnine_unit ninexnine_unit_7164(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C11R)
);

ninexnine_unit ninexnine_unit_7165(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D11R)
);

ninexnine_unit ninexnine_unit_7166(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E11R)
);

ninexnine_unit ninexnine_unit_7167(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F11R)
);

assign C311R=c3011R+c3111R+c3211R+c3311R+c3411R+c3511R+c3611R+c3711R+c3811R+c3911R+c3A11R+c3B11R+c3C11R+c3D11R+c3E11R+c3F11R;
assign A311R=(C311R>=0)?1:0;

assign P411R=A311R;

ninexnine_unit ninexnine_unit_7168(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3012R)
);

ninexnine_unit ninexnine_unit_7169(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3112R)
);

ninexnine_unit ninexnine_unit_7170(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3212R)
);

ninexnine_unit ninexnine_unit_7171(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3312R)
);

ninexnine_unit ninexnine_unit_7172(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3412R)
);

ninexnine_unit ninexnine_unit_7173(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3512R)
);

ninexnine_unit ninexnine_unit_7174(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3612R)
);

ninexnine_unit ninexnine_unit_7175(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3712R)
);

ninexnine_unit ninexnine_unit_7176(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3812R)
);

ninexnine_unit ninexnine_unit_7177(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3912R)
);

ninexnine_unit ninexnine_unit_7178(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A12R)
);

ninexnine_unit ninexnine_unit_7179(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B12R)
);

ninexnine_unit ninexnine_unit_7180(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C12R)
);

ninexnine_unit ninexnine_unit_7181(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D12R)
);

ninexnine_unit ninexnine_unit_7182(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E12R)
);

ninexnine_unit ninexnine_unit_7183(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F12R)
);

assign C312R=c3012R+c3112R+c3212R+c3312R+c3412R+c3512R+c3612R+c3712R+c3812R+c3912R+c3A12R+c3B12R+c3C12R+c3D12R+c3E12R+c3F12R;
assign A312R=(C312R>=0)?1:0;

assign P412R=A312R;

ninexnine_unit ninexnine_unit_7184(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3020R)
);

ninexnine_unit ninexnine_unit_7185(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3120R)
);

ninexnine_unit ninexnine_unit_7186(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3220R)
);

ninexnine_unit ninexnine_unit_7187(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3320R)
);

ninexnine_unit ninexnine_unit_7188(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3420R)
);

ninexnine_unit ninexnine_unit_7189(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3520R)
);

ninexnine_unit ninexnine_unit_7190(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3620R)
);

ninexnine_unit ninexnine_unit_7191(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3720R)
);

ninexnine_unit ninexnine_unit_7192(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3820R)
);

ninexnine_unit ninexnine_unit_7193(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3920R)
);

ninexnine_unit ninexnine_unit_7194(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A20R)
);

ninexnine_unit ninexnine_unit_7195(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B20R)
);

ninexnine_unit ninexnine_unit_7196(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C20R)
);

ninexnine_unit ninexnine_unit_7197(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D20R)
);

ninexnine_unit ninexnine_unit_7198(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E20R)
);

ninexnine_unit ninexnine_unit_7199(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F20R)
);

assign C320R=c3020R+c3120R+c3220R+c3320R+c3420R+c3520R+c3620R+c3720R+c3820R+c3920R+c3A20R+c3B20R+c3C20R+c3D20R+c3E20R+c3F20R;
assign A320R=(C320R>=0)?1:0;

assign P420R=A320R;

ninexnine_unit ninexnine_unit_7200(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3021R)
);

ninexnine_unit ninexnine_unit_7201(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3121R)
);

ninexnine_unit ninexnine_unit_7202(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3221R)
);

ninexnine_unit ninexnine_unit_7203(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3321R)
);

ninexnine_unit ninexnine_unit_7204(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3421R)
);

ninexnine_unit ninexnine_unit_7205(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3521R)
);

ninexnine_unit ninexnine_unit_7206(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3621R)
);

ninexnine_unit ninexnine_unit_7207(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3721R)
);

ninexnine_unit ninexnine_unit_7208(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3821R)
);

ninexnine_unit ninexnine_unit_7209(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3921R)
);

ninexnine_unit ninexnine_unit_7210(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A21R)
);

ninexnine_unit ninexnine_unit_7211(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B21R)
);

ninexnine_unit ninexnine_unit_7212(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C21R)
);

ninexnine_unit ninexnine_unit_7213(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D21R)
);

ninexnine_unit ninexnine_unit_7214(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E21R)
);

ninexnine_unit ninexnine_unit_7215(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F21R)
);

assign C321R=c3021R+c3121R+c3221R+c3321R+c3421R+c3521R+c3621R+c3721R+c3821R+c3921R+c3A21R+c3B21R+c3C21R+c3D21R+c3E21R+c3F21R;
assign A321R=(C321R>=0)?1:0;

assign P421R=A321R;

ninexnine_unit ninexnine_unit_7216(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3R000),
				.b1(W3R010),
				.b2(W3R020),
				.b3(W3R100),
				.b4(W3R110),
				.b5(W3R120),
				.b6(W3R200),
				.b7(W3R210),
				.b8(W3R220),
				.c(c3022R)
);

ninexnine_unit ninexnine_unit_7217(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3R001),
				.b1(W3R011),
				.b2(W3R021),
				.b3(W3R101),
				.b4(W3R111),
				.b5(W3R121),
				.b6(W3R201),
				.b7(W3R211),
				.b8(W3R221),
				.c(c3122R)
);

ninexnine_unit ninexnine_unit_7218(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3R002),
				.b1(W3R012),
				.b2(W3R022),
				.b3(W3R102),
				.b4(W3R112),
				.b5(W3R122),
				.b6(W3R202),
				.b7(W3R212),
				.b8(W3R222),
				.c(c3222R)
);

ninexnine_unit ninexnine_unit_7219(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3R003),
				.b1(W3R013),
				.b2(W3R023),
				.b3(W3R103),
				.b4(W3R113),
				.b5(W3R123),
				.b6(W3R203),
				.b7(W3R213),
				.b8(W3R223),
				.c(c3322R)
);

ninexnine_unit ninexnine_unit_7220(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3R004),
				.b1(W3R014),
				.b2(W3R024),
				.b3(W3R104),
				.b4(W3R114),
				.b5(W3R124),
				.b6(W3R204),
				.b7(W3R214),
				.b8(W3R224),
				.c(c3422R)
);

ninexnine_unit ninexnine_unit_7221(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3R005),
				.b1(W3R015),
				.b2(W3R025),
				.b3(W3R105),
				.b4(W3R115),
				.b5(W3R125),
				.b6(W3R205),
				.b7(W3R215),
				.b8(W3R225),
				.c(c3522R)
);

ninexnine_unit ninexnine_unit_7222(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3R006),
				.b1(W3R016),
				.b2(W3R026),
				.b3(W3R106),
				.b4(W3R116),
				.b5(W3R126),
				.b6(W3R206),
				.b7(W3R216),
				.b8(W3R226),
				.c(c3622R)
);

ninexnine_unit ninexnine_unit_7223(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3R007),
				.b1(W3R017),
				.b2(W3R027),
				.b3(W3R107),
				.b4(W3R117),
				.b5(W3R127),
				.b6(W3R207),
				.b7(W3R217),
				.b8(W3R227),
				.c(c3722R)
);

ninexnine_unit ninexnine_unit_7224(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3R008),
				.b1(W3R018),
				.b2(W3R028),
				.b3(W3R108),
				.b4(W3R118),
				.b5(W3R128),
				.b6(W3R208),
				.b7(W3R218),
				.b8(W3R228),
				.c(c3822R)
);

ninexnine_unit ninexnine_unit_7225(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3R009),
				.b1(W3R019),
				.b2(W3R029),
				.b3(W3R109),
				.b4(W3R119),
				.b5(W3R129),
				.b6(W3R209),
				.b7(W3R219),
				.b8(W3R229),
				.c(c3922R)
);

ninexnine_unit ninexnine_unit_7226(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3R00A),
				.b1(W3R01A),
				.b2(W3R02A),
				.b3(W3R10A),
				.b4(W3R11A),
				.b5(W3R12A),
				.b6(W3R20A),
				.b7(W3R21A),
				.b8(W3R22A),
				.c(c3A22R)
);

ninexnine_unit ninexnine_unit_7227(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3R00B),
				.b1(W3R01B),
				.b2(W3R02B),
				.b3(W3R10B),
				.b4(W3R11B),
				.b5(W3R12B),
				.b6(W3R20B),
				.b7(W3R21B),
				.b8(W3R22B),
				.c(c3B22R)
);

ninexnine_unit ninexnine_unit_7228(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3R00C),
				.b1(W3R01C),
				.b2(W3R02C),
				.b3(W3R10C),
				.b4(W3R11C),
				.b5(W3R12C),
				.b6(W3R20C),
				.b7(W3R21C),
				.b8(W3R22C),
				.c(c3C22R)
);

ninexnine_unit ninexnine_unit_7229(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3R00D),
				.b1(W3R01D),
				.b2(W3R02D),
				.b3(W3R10D),
				.b4(W3R11D),
				.b5(W3R12D),
				.b6(W3R20D),
				.b7(W3R21D),
				.b8(W3R22D),
				.c(c3D22R)
);

ninexnine_unit ninexnine_unit_7230(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3R00E),
				.b1(W3R01E),
				.b2(W3R02E),
				.b3(W3R10E),
				.b4(W3R11E),
				.b5(W3R12E),
				.b6(W3R20E),
				.b7(W3R21E),
				.b8(W3R22E),
				.c(c3E22R)
);

ninexnine_unit ninexnine_unit_7231(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3R00F),
				.b1(W3R01F),
				.b2(W3R02F),
				.b3(W3R10F),
				.b4(W3R11F),
				.b5(W3R12F),
				.b6(W3R20F),
				.b7(W3R21F),
				.b8(W3R22F),
				.c(c3F22R)
);

assign C322R=c3022R+c3122R+c3222R+c3322R+c3422R+c3522R+c3622R+c3722R+c3822R+c3922R+c3A22R+c3B22R+c3C22R+c3D22R+c3E22R+c3F22R;
assign A322R=(C322R>=0)?1:0;

assign P422R=A322R;

ninexnine_unit ninexnine_unit_7232(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3000S)
);

ninexnine_unit ninexnine_unit_7233(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3100S)
);

ninexnine_unit ninexnine_unit_7234(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3200S)
);

ninexnine_unit ninexnine_unit_7235(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3300S)
);

ninexnine_unit ninexnine_unit_7236(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3400S)
);

ninexnine_unit ninexnine_unit_7237(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3500S)
);

ninexnine_unit ninexnine_unit_7238(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3600S)
);

ninexnine_unit ninexnine_unit_7239(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3700S)
);

ninexnine_unit ninexnine_unit_7240(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3800S)
);

ninexnine_unit ninexnine_unit_7241(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3900S)
);

ninexnine_unit ninexnine_unit_7242(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A00S)
);

ninexnine_unit ninexnine_unit_7243(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B00S)
);

ninexnine_unit ninexnine_unit_7244(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C00S)
);

ninexnine_unit ninexnine_unit_7245(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D00S)
);

ninexnine_unit ninexnine_unit_7246(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E00S)
);

ninexnine_unit ninexnine_unit_7247(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F00S)
);

assign C300S=c3000S+c3100S+c3200S+c3300S+c3400S+c3500S+c3600S+c3700S+c3800S+c3900S+c3A00S+c3B00S+c3C00S+c3D00S+c3E00S+c3F00S;
assign A300S=(C300S>=0)?1:0;

assign P400S=A300S;

ninexnine_unit ninexnine_unit_7248(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3001S)
);

ninexnine_unit ninexnine_unit_7249(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3101S)
);

ninexnine_unit ninexnine_unit_7250(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3201S)
);

ninexnine_unit ninexnine_unit_7251(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3301S)
);

ninexnine_unit ninexnine_unit_7252(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3401S)
);

ninexnine_unit ninexnine_unit_7253(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3501S)
);

ninexnine_unit ninexnine_unit_7254(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3601S)
);

ninexnine_unit ninexnine_unit_7255(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3701S)
);

ninexnine_unit ninexnine_unit_7256(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3801S)
);

ninexnine_unit ninexnine_unit_7257(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3901S)
);

ninexnine_unit ninexnine_unit_7258(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A01S)
);

ninexnine_unit ninexnine_unit_7259(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B01S)
);

ninexnine_unit ninexnine_unit_7260(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C01S)
);

ninexnine_unit ninexnine_unit_7261(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D01S)
);

ninexnine_unit ninexnine_unit_7262(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E01S)
);

ninexnine_unit ninexnine_unit_7263(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F01S)
);

assign C301S=c3001S+c3101S+c3201S+c3301S+c3401S+c3501S+c3601S+c3701S+c3801S+c3901S+c3A01S+c3B01S+c3C01S+c3D01S+c3E01S+c3F01S;
assign A301S=(C301S>=0)?1:0;

assign P401S=A301S;

ninexnine_unit ninexnine_unit_7264(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3002S)
);

ninexnine_unit ninexnine_unit_7265(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3102S)
);

ninexnine_unit ninexnine_unit_7266(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3202S)
);

ninexnine_unit ninexnine_unit_7267(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3302S)
);

ninexnine_unit ninexnine_unit_7268(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3402S)
);

ninexnine_unit ninexnine_unit_7269(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3502S)
);

ninexnine_unit ninexnine_unit_7270(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3602S)
);

ninexnine_unit ninexnine_unit_7271(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3702S)
);

ninexnine_unit ninexnine_unit_7272(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3802S)
);

ninexnine_unit ninexnine_unit_7273(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3902S)
);

ninexnine_unit ninexnine_unit_7274(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A02S)
);

ninexnine_unit ninexnine_unit_7275(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B02S)
);

ninexnine_unit ninexnine_unit_7276(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C02S)
);

ninexnine_unit ninexnine_unit_7277(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D02S)
);

ninexnine_unit ninexnine_unit_7278(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E02S)
);

ninexnine_unit ninexnine_unit_7279(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F02S)
);

assign C302S=c3002S+c3102S+c3202S+c3302S+c3402S+c3502S+c3602S+c3702S+c3802S+c3902S+c3A02S+c3B02S+c3C02S+c3D02S+c3E02S+c3F02S;
assign A302S=(C302S>=0)?1:0;

assign P402S=A302S;

ninexnine_unit ninexnine_unit_7280(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3010S)
);

ninexnine_unit ninexnine_unit_7281(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3110S)
);

ninexnine_unit ninexnine_unit_7282(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3210S)
);

ninexnine_unit ninexnine_unit_7283(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3310S)
);

ninexnine_unit ninexnine_unit_7284(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3410S)
);

ninexnine_unit ninexnine_unit_7285(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3510S)
);

ninexnine_unit ninexnine_unit_7286(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3610S)
);

ninexnine_unit ninexnine_unit_7287(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3710S)
);

ninexnine_unit ninexnine_unit_7288(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3810S)
);

ninexnine_unit ninexnine_unit_7289(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3910S)
);

ninexnine_unit ninexnine_unit_7290(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A10S)
);

ninexnine_unit ninexnine_unit_7291(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B10S)
);

ninexnine_unit ninexnine_unit_7292(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C10S)
);

ninexnine_unit ninexnine_unit_7293(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D10S)
);

ninexnine_unit ninexnine_unit_7294(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E10S)
);

ninexnine_unit ninexnine_unit_7295(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F10S)
);

assign C310S=c3010S+c3110S+c3210S+c3310S+c3410S+c3510S+c3610S+c3710S+c3810S+c3910S+c3A10S+c3B10S+c3C10S+c3D10S+c3E10S+c3F10S;
assign A310S=(C310S>=0)?1:0;

assign P410S=A310S;

ninexnine_unit ninexnine_unit_7296(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3011S)
);

ninexnine_unit ninexnine_unit_7297(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3111S)
);

ninexnine_unit ninexnine_unit_7298(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3211S)
);

ninexnine_unit ninexnine_unit_7299(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3311S)
);

ninexnine_unit ninexnine_unit_7300(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3411S)
);

ninexnine_unit ninexnine_unit_7301(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3511S)
);

ninexnine_unit ninexnine_unit_7302(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3611S)
);

ninexnine_unit ninexnine_unit_7303(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3711S)
);

ninexnine_unit ninexnine_unit_7304(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3811S)
);

ninexnine_unit ninexnine_unit_7305(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3911S)
);

ninexnine_unit ninexnine_unit_7306(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A11S)
);

ninexnine_unit ninexnine_unit_7307(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B11S)
);

ninexnine_unit ninexnine_unit_7308(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C11S)
);

ninexnine_unit ninexnine_unit_7309(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D11S)
);

ninexnine_unit ninexnine_unit_7310(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E11S)
);

ninexnine_unit ninexnine_unit_7311(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F11S)
);

assign C311S=c3011S+c3111S+c3211S+c3311S+c3411S+c3511S+c3611S+c3711S+c3811S+c3911S+c3A11S+c3B11S+c3C11S+c3D11S+c3E11S+c3F11S;
assign A311S=(C311S>=0)?1:0;

assign P411S=A311S;

ninexnine_unit ninexnine_unit_7312(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3012S)
);

ninexnine_unit ninexnine_unit_7313(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3112S)
);

ninexnine_unit ninexnine_unit_7314(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3212S)
);

ninexnine_unit ninexnine_unit_7315(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3312S)
);

ninexnine_unit ninexnine_unit_7316(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3412S)
);

ninexnine_unit ninexnine_unit_7317(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3512S)
);

ninexnine_unit ninexnine_unit_7318(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3612S)
);

ninexnine_unit ninexnine_unit_7319(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3712S)
);

ninexnine_unit ninexnine_unit_7320(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3812S)
);

ninexnine_unit ninexnine_unit_7321(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3912S)
);

ninexnine_unit ninexnine_unit_7322(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A12S)
);

ninexnine_unit ninexnine_unit_7323(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B12S)
);

ninexnine_unit ninexnine_unit_7324(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C12S)
);

ninexnine_unit ninexnine_unit_7325(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D12S)
);

ninexnine_unit ninexnine_unit_7326(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E12S)
);

ninexnine_unit ninexnine_unit_7327(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F12S)
);

assign C312S=c3012S+c3112S+c3212S+c3312S+c3412S+c3512S+c3612S+c3712S+c3812S+c3912S+c3A12S+c3B12S+c3C12S+c3D12S+c3E12S+c3F12S;
assign A312S=(C312S>=0)?1:0;

assign P412S=A312S;

ninexnine_unit ninexnine_unit_7328(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3020S)
);

ninexnine_unit ninexnine_unit_7329(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3120S)
);

ninexnine_unit ninexnine_unit_7330(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3220S)
);

ninexnine_unit ninexnine_unit_7331(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3320S)
);

ninexnine_unit ninexnine_unit_7332(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3420S)
);

ninexnine_unit ninexnine_unit_7333(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3520S)
);

ninexnine_unit ninexnine_unit_7334(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3620S)
);

ninexnine_unit ninexnine_unit_7335(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3720S)
);

ninexnine_unit ninexnine_unit_7336(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3820S)
);

ninexnine_unit ninexnine_unit_7337(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3920S)
);

ninexnine_unit ninexnine_unit_7338(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A20S)
);

ninexnine_unit ninexnine_unit_7339(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B20S)
);

ninexnine_unit ninexnine_unit_7340(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C20S)
);

ninexnine_unit ninexnine_unit_7341(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D20S)
);

ninexnine_unit ninexnine_unit_7342(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E20S)
);

ninexnine_unit ninexnine_unit_7343(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F20S)
);

assign C320S=c3020S+c3120S+c3220S+c3320S+c3420S+c3520S+c3620S+c3720S+c3820S+c3920S+c3A20S+c3B20S+c3C20S+c3D20S+c3E20S+c3F20S;
assign A320S=(C320S>=0)?1:0;

assign P420S=A320S;

ninexnine_unit ninexnine_unit_7344(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3021S)
);

ninexnine_unit ninexnine_unit_7345(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3121S)
);

ninexnine_unit ninexnine_unit_7346(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3221S)
);

ninexnine_unit ninexnine_unit_7347(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3321S)
);

ninexnine_unit ninexnine_unit_7348(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3421S)
);

ninexnine_unit ninexnine_unit_7349(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3521S)
);

ninexnine_unit ninexnine_unit_7350(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3621S)
);

ninexnine_unit ninexnine_unit_7351(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3721S)
);

ninexnine_unit ninexnine_unit_7352(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3821S)
);

ninexnine_unit ninexnine_unit_7353(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3921S)
);

ninexnine_unit ninexnine_unit_7354(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A21S)
);

ninexnine_unit ninexnine_unit_7355(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B21S)
);

ninexnine_unit ninexnine_unit_7356(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C21S)
);

ninexnine_unit ninexnine_unit_7357(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D21S)
);

ninexnine_unit ninexnine_unit_7358(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E21S)
);

ninexnine_unit ninexnine_unit_7359(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F21S)
);

assign C321S=c3021S+c3121S+c3221S+c3321S+c3421S+c3521S+c3621S+c3721S+c3821S+c3921S+c3A21S+c3B21S+c3C21S+c3D21S+c3E21S+c3F21S;
assign A321S=(C321S>=0)?1:0;

assign P421S=A321S;

ninexnine_unit ninexnine_unit_7360(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3S000),
				.b1(W3S010),
				.b2(W3S020),
				.b3(W3S100),
				.b4(W3S110),
				.b5(W3S120),
				.b6(W3S200),
				.b7(W3S210),
				.b8(W3S220),
				.c(c3022S)
);

ninexnine_unit ninexnine_unit_7361(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3S001),
				.b1(W3S011),
				.b2(W3S021),
				.b3(W3S101),
				.b4(W3S111),
				.b5(W3S121),
				.b6(W3S201),
				.b7(W3S211),
				.b8(W3S221),
				.c(c3122S)
);

ninexnine_unit ninexnine_unit_7362(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3S002),
				.b1(W3S012),
				.b2(W3S022),
				.b3(W3S102),
				.b4(W3S112),
				.b5(W3S122),
				.b6(W3S202),
				.b7(W3S212),
				.b8(W3S222),
				.c(c3222S)
);

ninexnine_unit ninexnine_unit_7363(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3S003),
				.b1(W3S013),
				.b2(W3S023),
				.b3(W3S103),
				.b4(W3S113),
				.b5(W3S123),
				.b6(W3S203),
				.b7(W3S213),
				.b8(W3S223),
				.c(c3322S)
);

ninexnine_unit ninexnine_unit_7364(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3S004),
				.b1(W3S014),
				.b2(W3S024),
				.b3(W3S104),
				.b4(W3S114),
				.b5(W3S124),
				.b6(W3S204),
				.b7(W3S214),
				.b8(W3S224),
				.c(c3422S)
);

ninexnine_unit ninexnine_unit_7365(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3S005),
				.b1(W3S015),
				.b2(W3S025),
				.b3(W3S105),
				.b4(W3S115),
				.b5(W3S125),
				.b6(W3S205),
				.b7(W3S215),
				.b8(W3S225),
				.c(c3522S)
);

ninexnine_unit ninexnine_unit_7366(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3S006),
				.b1(W3S016),
				.b2(W3S026),
				.b3(W3S106),
				.b4(W3S116),
				.b5(W3S126),
				.b6(W3S206),
				.b7(W3S216),
				.b8(W3S226),
				.c(c3622S)
);

ninexnine_unit ninexnine_unit_7367(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3S007),
				.b1(W3S017),
				.b2(W3S027),
				.b3(W3S107),
				.b4(W3S117),
				.b5(W3S127),
				.b6(W3S207),
				.b7(W3S217),
				.b8(W3S227),
				.c(c3722S)
);

ninexnine_unit ninexnine_unit_7368(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3S008),
				.b1(W3S018),
				.b2(W3S028),
				.b3(W3S108),
				.b4(W3S118),
				.b5(W3S128),
				.b6(W3S208),
				.b7(W3S218),
				.b8(W3S228),
				.c(c3822S)
);

ninexnine_unit ninexnine_unit_7369(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3S009),
				.b1(W3S019),
				.b2(W3S029),
				.b3(W3S109),
				.b4(W3S119),
				.b5(W3S129),
				.b6(W3S209),
				.b7(W3S219),
				.b8(W3S229),
				.c(c3922S)
);

ninexnine_unit ninexnine_unit_7370(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3S00A),
				.b1(W3S01A),
				.b2(W3S02A),
				.b3(W3S10A),
				.b4(W3S11A),
				.b5(W3S12A),
				.b6(W3S20A),
				.b7(W3S21A),
				.b8(W3S22A),
				.c(c3A22S)
);

ninexnine_unit ninexnine_unit_7371(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3S00B),
				.b1(W3S01B),
				.b2(W3S02B),
				.b3(W3S10B),
				.b4(W3S11B),
				.b5(W3S12B),
				.b6(W3S20B),
				.b7(W3S21B),
				.b8(W3S22B),
				.c(c3B22S)
);

ninexnine_unit ninexnine_unit_7372(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3S00C),
				.b1(W3S01C),
				.b2(W3S02C),
				.b3(W3S10C),
				.b4(W3S11C),
				.b5(W3S12C),
				.b6(W3S20C),
				.b7(W3S21C),
				.b8(W3S22C),
				.c(c3C22S)
);

ninexnine_unit ninexnine_unit_7373(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3S00D),
				.b1(W3S01D),
				.b2(W3S02D),
				.b3(W3S10D),
				.b4(W3S11D),
				.b5(W3S12D),
				.b6(W3S20D),
				.b7(W3S21D),
				.b8(W3S22D),
				.c(c3D22S)
);

ninexnine_unit ninexnine_unit_7374(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3S00E),
				.b1(W3S01E),
				.b2(W3S02E),
				.b3(W3S10E),
				.b4(W3S11E),
				.b5(W3S12E),
				.b6(W3S20E),
				.b7(W3S21E),
				.b8(W3S22E),
				.c(c3E22S)
);

ninexnine_unit ninexnine_unit_7375(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3S00F),
				.b1(W3S01F),
				.b2(W3S02F),
				.b3(W3S10F),
				.b4(W3S11F),
				.b5(W3S12F),
				.b6(W3S20F),
				.b7(W3S21F),
				.b8(W3S22F),
				.c(c3F22S)
);

assign C322S=c3022S+c3122S+c3222S+c3322S+c3422S+c3522S+c3622S+c3722S+c3822S+c3922S+c3A22S+c3B22S+c3C22S+c3D22S+c3E22S+c3F22S;
assign A322S=(C322S>=0)?1:0;

assign P422S=A322S;

ninexnine_unit ninexnine_unit_7376(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3000T)
);

ninexnine_unit ninexnine_unit_7377(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3100T)
);

ninexnine_unit ninexnine_unit_7378(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3200T)
);

ninexnine_unit ninexnine_unit_7379(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3300T)
);

ninexnine_unit ninexnine_unit_7380(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3400T)
);

ninexnine_unit ninexnine_unit_7381(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3500T)
);

ninexnine_unit ninexnine_unit_7382(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3600T)
);

ninexnine_unit ninexnine_unit_7383(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3700T)
);

ninexnine_unit ninexnine_unit_7384(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3800T)
);

ninexnine_unit ninexnine_unit_7385(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3900T)
);

ninexnine_unit ninexnine_unit_7386(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A00T)
);

ninexnine_unit ninexnine_unit_7387(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B00T)
);

ninexnine_unit ninexnine_unit_7388(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C00T)
);

ninexnine_unit ninexnine_unit_7389(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D00T)
);

ninexnine_unit ninexnine_unit_7390(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E00T)
);

ninexnine_unit ninexnine_unit_7391(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F00T)
);

assign C300T=c3000T+c3100T+c3200T+c3300T+c3400T+c3500T+c3600T+c3700T+c3800T+c3900T+c3A00T+c3B00T+c3C00T+c3D00T+c3E00T+c3F00T;
assign A300T=(C300T>=0)?1:0;

assign P400T=A300T;

ninexnine_unit ninexnine_unit_7392(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3001T)
);

ninexnine_unit ninexnine_unit_7393(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3101T)
);

ninexnine_unit ninexnine_unit_7394(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3201T)
);

ninexnine_unit ninexnine_unit_7395(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3301T)
);

ninexnine_unit ninexnine_unit_7396(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3401T)
);

ninexnine_unit ninexnine_unit_7397(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3501T)
);

ninexnine_unit ninexnine_unit_7398(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3601T)
);

ninexnine_unit ninexnine_unit_7399(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3701T)
);

ninexnine_unit ninexnine_unit_7400(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3801T)
);

ninexnine_unit ninexnine_unit_7401(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3901T)
);

ninexnine_unit ninexnine_unit_7402(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A01T)
);

ninexnine_unit ninexnine_unit_7403(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B01T)
);

ninexnine_unit ninexnine_unit_7404(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C01T)
);

ninexnine_unit ninexnine_unit_7405(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D01T)
);

ninexnine_unit ninexnine_unit_7406(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E01T)
);

ninexnine_unit ninexnine_unit_7407(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F01T)
);

assign C301T=c3001T+c3101T+c3201T+c3301T+c3401T+c3501T+c3601T+c3701T+c3801T+c3901T+c3A01T+c3B01T+c3C01T+c3D01T+c3E01T+c3F01T;
assign A301T=(C301T>=0)?1:0;

assign P401T=A301T;

ninexnine_unit ninexnine_unit_7408(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3002T)
);

ninexnine_unit ninexnine_unit_7409(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3102T)
);

ninexnine_unit ninexnine_unit_7410(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3202T)
);

ninexnine_unit ninexnine_unit_7411(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3302T)
);

ninexnine_unit ninexnine_unit_7412(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3402T)
);

ninexnine_unit ninexnine_unit_7413(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3502T)
);

ninexnine_unit ninexnine_unit_7414(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3602T)
);

ninexnine_unit ninexnine_unit_7415(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3702T)
);

ninexnine_unit ninexnine_unit_7416(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3802T)
);

ninexnine_unit ninexnine_unit_7417(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3902T)
);

ninexnine_unit ninexnine_unit_7418(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A02T)
);

ninexnine_unit ninexnine_unit_7419(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B02T)
);

ninexnine_unit ninexnine_unit_7420(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C02T)
);

ninexnine_unit ninexnine_unit_7421(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D02T)
);

ninexnine_unit ninexnine_unit_7422(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E02T)
);

ninexnine_unit ninexnine_unit_7423(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F02T)
);

assign C302T=c3002T+c3102T+c3202T+c3302T+c3402T+c3502T+c3602T+c3702T+c3802T+c3902T+c3A02T+c3B02T+c3C02T+c3D02T+c3E02T+c3F02T;
assign A302T=(C302T>=0)?1:0;

assign P402T=A302T;

ninexnine_unit ninexnine_unit_7424(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3010T)
);

ninexnine_unit ninexnine_unit_7425(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3110T)
);

ninexnine_unit ninexnine_unit_7426(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3210T)
);

ninexnine_unit ninexnine_unit_7427(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3310T)
);

ninexnine_unit ninexnine_unit_7428(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3410T)
);

ninexnine_unit ninexnine_unit_7429(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3510T)
);

ninexnine_unit ninexnine_unit_7430(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3610T)
);

ninexnine_unit ninexnine_unit_7431(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3710T)
);

ninexnine_unit ninexnine_unit_7432(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3810T)
);

ninexnine_unit ninexnine_unit_7433(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3910T)
);

ninexnine_unit ninexnine_unit_7434(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A10T)
);

ninexnine_unit ninexnine_unit_7435(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B10T)
);

ninexnine_unit ninexnine_unit_7436(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C10T)
);

ninexnine_unit ninexnine_unit_7437(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D10T)
);

ninexnine_unit ninexnine_unit_7438(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E10T)
);

ninexnine_unit ninexnine_unit_7439(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F10T)
);

assign C310T=c3010T+c3110T+c3210T+c3310T+c3410T+c3510T+c3610T+c3710T+c3810T+c3910T+c3A10T+c3B10T+c3C10T+c3D10T+c3E10T+c3F10T;
assign A310T=(C310T>=0)?1:0;

assign P410T=A310T;

ninexnine_unit ninexnine_unit_7440(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3011T)
);

ninexnine_unit ninexnine_unit_7441(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3111T)
);

ninexnine_unit ninexnine_unit_7442(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3211T)
);

ninexnine_unit ninexnine_unit_7443(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3311T)
);

ninexnine_unit ninexnine_unit_7444(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3411T)
);

ninexnine_unit ninexnine_unit_7445(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3511T)
);

ninexnine_unit ninexnine_unit_7446(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3611T)
);

ninexnine_unit ninexnine_unit_7447(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3711T)
);

ninexnine_unit ninexnine_unit_7448(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3811T)
);

ninexnine_unit ninexnine_unit_7449(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3911T)
);

ninexnine_unit ninexnine_unit_7450(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A11T)
);

ninexnine_unit ninexnine_unit_7451(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B11T)
);

ninexnine_unit ninexnine_unit_7452(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C11T)
);

ninexnine_unit ninexnine_unit_7453(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D11T)
);

ninexnine_unit ninexnine_unit_7454(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E11T)
);

ninexnine_unit ninexnine_unit_7455(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F11T)
);

assign C311T=c3011T+c3111T+c3211T+c3311T+c3411T+c3511T+c3611T+c3711T+c3811T+c3911T+c3A11T+c3B11T+c3C11T+c3D11T+c3E11T+c3F11T;
assign A311T=(C311T>=0)?1:0;

assign P411T=A311T;

ninexnine_unit ninexnine_unit_7456(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3012T)
);

ninexnine_unit ninexnine_unit_7457(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3112T)
);

ninexnine_unit ninexnine_unit_7458(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3212T)
);

ninexnine_unit ninexnine_unit_7459(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3312T)
);

ninexnine_unit ninexnine_unit_7460(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3412T)
);

ninexnine_unit ninexnine_unit_7461(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3512T)
);

ninexnine_unit ninexnine_unit_7462(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3612T)
);

ninexnine_unit ninexnine_unit_7463(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3712T)
);

ninexnine_unit ninexnine_unit_7464(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3812T)
);

ninexnine_unit ninexnine_unit_7465(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3912T)
);

ninexnine_unit ninexnine_unit_7466(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A12T)
);

ninexnine_unit ninexnine_unit_7467(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B12T)
);

ninexnine_unit ninexnine_unit_7468(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C12T)
);

ninexnine_unit ninexnine_unit_7469(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D12T)
);

ninexnine_unit ninexnine_unit_7470(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E12T)
);

ninexnine_unit ninexnine_unit_7471(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F12T)
);

assign C312T=c3012T+c3112T+c3212T+c3312T+c3412T+c3512T+c3612T+c3712T+c3812T+c3912T+c3A12T+c3B12T+c3C12T+c3D12T+c3E12T+c3F12T;
assign A312T=(C312T>=0)?1:0;

assign P412T=A312T;

ninexnine_unit ninexnine_unit_7472(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3020T)
);

ninexnine_unit ninexnine_unit_7473(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3120T)
);

ninexnine_unit ninexnine_unit_7474(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3220T)
);

ninexnine_unit ninexnine_unit_7475(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3320T)
);

ninexnine_unit ninexnine_unit_7476(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3420T)
);

ninexnine_unit ninexnine_unit_7477(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3520T)
);

ninexnine_unit ninexnine_unit_7478(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3620T)
);

ninexnine_unit ninexnine_unit_7479(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3720T)
);

ninexnine_unit ninexnine_unit_7480(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3820T)
);

ninexnine_unit ninexnine_unit_7481(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3920T)
);

ninexnine_unit ninexnine_unit_7482(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A20T)
);

ninexnine_unit ninexnine_unit_7483(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B20T)
);

ninexnine_unit ninexnine_unit_7484(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C20T)
);

ninexnine_unit ninexnine_unit_7485(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D20T)
);

ninexnine_unit ninexnine_unit_7486(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E20T)
);

ninexnine_unit ninexnine_unit_7487(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F20T)
);

assign C320T=c3020T+c3120T+c3220T+c3320T+c3420T+c3520T+c3620T+c3720T+c3820T+c3920T+c3A20T+c3B20T+c3C20T+c3D20T+c3E20T+c3F20T;
assign A320T=(C320T>=0)?1:0;

assign P420T=A320T;

ninexnine_unit ninexnine_unit_7488(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3021T)
);

ninexnine_unit ninexnine_unit_7489(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3121T)
);

ninexnine_unit ninexnine_unit_7490(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3221T)
);

ninexnine_unit ninexnine_unit_7491(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3321T)
);

ninexnine_unit ninexnine_unit_7492(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3421T)
);

ninexnine_unit ninexnine_unit_7493(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3521T)
);

ninexnine_unit ninexnine_unit_7494(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3621T)
);

ninexnine_unit ninexnine_unit_7495(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3721T)
);

ninexnine_unit ninexnine_unit_7496(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3821T)
);

ninexnine_unit ninexnine_unit_7497(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3921T)
);

ninexnine_unit ninexnine_unit_7498(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A21T)
);

ninexnine_unit ninexnine_unit_7499(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B21T)
);

ninexnine_unit ninexnine_unit_7500(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C21T)
);

ninexnine_unit ninexnine_unit_7501(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D21T)
);

ninexnine_unit ninexnine_unit_7502(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E21T)
);

ninexnine_unit ninexnine_unit_7503(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F21T)
);

assign C321T=c3021T+c3121T+c3221T+c3321T+c3421T+c3521T+c3621T+c3721T+c3821T+c3921T+c3A21T+c3B21T+c3C21T+c3D21T+c3E21T+c3F21T;
assign A321T=(C321T>=0)?1:0;

assign P421T=A321T;

ninexnine_unit ninexnine_unit_7504(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3T000),
				.b1(W3T010),
				.b2(W3T020),
				.b3(W3T100),
				.b4(W3T110),
				.b5(W3T120),
				.b6(W3T200),
				.b7(W3T210),
				.b8(W3T220),
				.c(c3022T)
);

ninexnine_unit ninexnine_unit_7505(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3T001),
				.b1(W3T011),
				.b2(W3T021),
				.b3(W3T101),
				.b4(W3T111),
				.b5(W3T121),
				.b6(W3T201),
				.b7(W3T211),
				.b8(W3T221),
				.c(c3122T)
);

ninexnine_unit ninexnine_unit_7506(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3T002),
				.b1(W3T012),
				.b2(W3T022),
				.b3(W3T102),
				.b4(W3T112),
				.b5(W3T122),
				.b6(W3T202),
				.b7(W3T212),
				.b8(W3T222),
				.c(c3222T)
);

ninexnine_unit ninexnine_unit_7507(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3T003),
				.b1(W3T013),
				.b2(W3T023),
				.b3(W3T103),
				.b4(W3T113),
				.b5(W3T123),
				.b6(W3T203),
				.b7(W3T213),
				.b8(W3T223),
				.c(c3322T)
);

ninexnine_unit ninexnine_unit_7508(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3T004),
				.b1(W3T014),
				.b2(W3T024),
				.b3(W3T104),
				.b4(W3T114),
				.b5(W3T124),
				.b6(W3T204),
				.b7(W3T214),
				.b8(W3T224),
				.c(c3422T)
);

ninexnine_unit ninexnine_unit_7509(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3T005),
				.b1(W3T015),
				.b2(W3T025),
				.b3(W3T105),
				.b4(W3T115),
				.b5(W3T125),
				.b6(W3T205),
				.b7(W3T215),
				.b8(W3T225),
				.c(c3522T)
);

ninexnine_unit ninexnine_unit_7510(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3T006),
				.b1(W3T016),
				.b2(W3T026),
				.b3(W3T106),
				.b4(W3T116),
				.b5(W3T126),
				.b6(W3T206),
				.b7(W3T216),
				.b8(W3T226),
				.c(c3622T)
);

ninexnine_unit ninexnine_unit_7511(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3T007),
				.b1(W3T017),
				.b2(W3T027),
				.b3(W3T107),
				.b4(W3T117),
				.b5(W3T127),
				.b6(W3T207),
				.b7(W3T217),
				.b8(W3T227),
				.c(c3722T)
);

ninexnine_unit ninexnine_unit_7512(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3T008),
				.b1(W3T018),
				.b2(W3T028),
				.b3(W3T108),
				.b4(W3T118),
				.b5(W3T128),
				.b6(W3T208),
				.b7(W3T218),
				.b8(W3T228),
				.c(c3822T)
);

ninexnine_unit ninexnine_unit_7513(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3T009),
				.b1(W3T019),
				.b2(W3T029),
				.b3(W3T109),
				.b4(W3T119),
				.b5(W3T129),
				.b6(W3T209),
				.b7(W3T219),
				.b8(W3T229),
				.c(c3922T)
);

ninexnine_unit ninexnine_unit_7514(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3T00A),
				.b1(W3T01A),
				.b2(W3T02A),
				.b3(W3T10A),
				.b4(W3T11A),
				.b5(W3T12A),
				.b6(W3T20A),
				.b7(W3T21A),
				.b8(W3T22A),
				.c(c3A22T)
);

ninexnine_unit ninexnine_unit_7515(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3T00B),
				.b1(W3T01B),
				.b2(W3T02B),
				.b3(W3T10B),
				.b4(W3T11B),
				.b5(W3T12B),
				.b6(W3T20B),
				.b7(W3T21B),
				.b8(W3T22B),
				.c(c3B22T)
);

ninexnine_unit ninexnine_unit_7516(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3T00C),
				.b1(W3T01C),
				.b2(W3T02C),
				.b3(W3T10C),
				.b4(W3T11C),
				.b5(W3T12C),
				.b6(W3T20C),
				.b7(W3T21C),
				.b8(W3T22C),
				.c(c3C22T)
);

ninexnine_unit ninexnine_unit_7517(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3T00D),
				.b1(W3T01D),
				.b2(W3T02D),
				.b3(W3T10D),
				.b4(W3T11D),
				.b5(W3T12D),
				.b6(W3T20D),
				.b7(W3T21D),
				.b8(W3T22D),
				.c(c3D22T)
);

ninexnine_unit ninexnine_unit_7518(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3T00E),
				.b1(W3T01E),
				.b2(W3T02E),
				.b3(W3T10E),
				.b4(W3T11E),
				.b5(W3T12E),
				.b6(W3T20E),
				.b7(W3T21E),
				.b8(W3T22E),
				.c(c3E22T)
);

ninexnine_unit ninexnine_unit_7519(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3T00F),
				.b1(W3T01F),
				.b2(W3T02F),
				.b3(W3T10F),
				.b4(W3T11F),
				.b5(W3T12F),
				.b6(W3T20F),
				.b7(W3T21F),
				.b8(W3T22F),
				.c(c3F22T)
);

assign C322T=c3022T+c3122T+c3222T+c3322T+c3422T+c3522T+c3622T+c3722T+c3822T+c3922T+c3A22T+c3B22T+c3C22T+c3D22T+c3E22T+c3F22T;
assign A322T=(C322T>=0)?1:0;

assign P422T=A322T;

ninexnine_unit ninexnine_unit_7520(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3000U)
);

ninexnine_unit ninexnine_unit_7521(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3100U)
);

ninexnine_unit ninexnine_unit_7522(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3200U)
);

ninexnine_unit ninexnine_unit_7523(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3300U)
);

ninexnine_unit ninexnine_unit_7524(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3400U)
);

ninexnine_unit ninexnine_unit_7525(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3500U)
);

ninexnine_unit ninexnine_unit_7526(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3600U)
);

ninexnine_unit ninexnine_unit_7527(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3700U)
);

ninexnine_unit ninexnine_unit_7528(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3800U)
);

ninexnine_unit ninexnine_unit_7529(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3900U)
);

ninexnine_unit ninexnine_unit_7530(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A00U)
);

ninexnine_unit ninexnine_unit_7531(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B00U)
);

ninexnine_unit ninexnine_unit_7532(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C00U)
);

ninexnine_unit ninexnine_unit_7533(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D00U)
);

ninexnine_unit ninexnine_unit_7534(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E00U)
);

ninexnine_unit ninexnine_unit_7535(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F00U)
);

assign C300U=c3000U+c3100U+c3200U+c3300U+c3400U+c3500U+c3600U+c3700U+c3800U+c3900U+c3A00U+c3B00U+c3C00U+c3D00U+c3E00U+c3F00U;
assign A300U=(C300U>=0)?1:0;

assign P400U=A300U;

ninexnine_unit ninexnine_unit_7536(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3001U)
);

ninexnine_unit ninexnine_unit_7537(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3101U)
);

ninexnine_unit ninexnine_unit_7538(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3201U)
);

ninexnine_unit ninexnine_unit_7539(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3301U)
);

ninexnine_unit ninexnine_unit_7540(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3401U)
);

ninexnine_unit ninexnine_unit_7541(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3501U)
);

ninexnine_unit ninexnine_unit_7542(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3601U)
);

ninexnine_unit ninexnine_unit_7543(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3701U)
);

ninexnine_unit ninexnine_unit_7544(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3801U)
);

ninexnine_unit ninexnine_unit_7545(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3901U)
);

ninexnine_unit ninexnine_unit_7546(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A01U)
);

ninexnine_unit ninexnine_unit_7547(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B01U)
);

ninexnine_unit ninexnine_unit_7548(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C01U)
);

ninexnine_unit ninexnine_unit_7549(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D01U)
);

ninexnine_unit ninexnine_unit_7550(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E01U)
);

ninexnine_unit ninexnine_unit_7551(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F01U)
);

assign C301U=c3001U+c3101U+c3201U+c3301U+c3401U+c3501U+c3601U+c3701U+c3801U+c3901U+c3A01U+c3B01U+c3C01U+c3D01U+c3E01U+c3F01U;
assign A301U=(C301U>=0)?1:0;

assign P401U=A301U;

ninexnine_unit ninexnine_unit_7552(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3002U)
);

ninexnine_unit ninexnine_unit_7553(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3102U)
);

ninexnine_unit ninexnine_unit_7554(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3202U)
);

ninexnine_unit ninexnine_unit_7555(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3302U)
);

ninexnine_unit ninexnine_unit_7556(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3402U)
);

ninexnine_unit ninexnine_unit_7557(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3502U)
);

ninexnine_unit ninexnine_unit_7558(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3602U)
);

ninexnine_unit ninexnine_unit_7559(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3702U)
);

ninexnine_unit ninexnine_unit_7560(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3802U)
);

ninexnine_unit ninexnine_unit_7561(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3902U)
);

ninexnine_unit ninexnine_unit_7562(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A02U)
);

ninexnine_unit ninexnine_unit_7563(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B02U)
);

ninexnine_unit ninexnine_unit_7564(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C02U)
);

ninexnine_unit ninexnine_unit_7565(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D02U)
);

ninexnine_unit ninexnine_unit_7566(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E02U)
);

ninexnine_unit ninexnine_unit_7567(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F02U)
);

assign C302U=c3002U+c3102U+c3202U+c3302U+c3402U+c3502U+c3602U+c3702U+c3802U+c3902U+c3A02U+c3B02U+c3C02U+c3D02U+c3E02U+c3F02U;
assign A302U=(C302U>=0)?1:0;

assign P402U=A302U;

ninexnine_unit ninexnine_unit_7568(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3010U)
);

ninexnine_unit ninexnine_unit_7569(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3110U)
);

ninexnine_unit ninexnine_unit_7570(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3210U)
);

ninexnine_unit ninexnine_unit_7571(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3310U)
);

ninexnine_unit ninexnine_unit_7572(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3410U)
);

ninexnine_unit ninexnine_unit_7573(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3510U)
);

ninexnine_unit ninexnine_unit_7574(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3610U)
);

ninexnine_unit ninexnine_unit_7575(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3710U)
);

ninexnine_unit ninexnine_unit_7576(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3810U)
);

ninexnine_unit ninexnine_unit_7577(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3910U)
);

ninexnine_unit ninexnine_unit_7578(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A10U)
);

ninexnine_unit ninexnine_unit_7579(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B10U)
);

ninexnine_unit ninexnine_unit_7580(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C10U)
);

ninexnine_unit ninexnine_unit_7581(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D10U)
);

ninexnine_unit ninexnine_unit_7582(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E10U)
);

ninexnine_unit ninexnine_unit_7583(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F10U)
);

assign C310U=c3010U+c3110U+c3210U+c3310U+c3410U+c3510U+c3610U+c3710U+c3810U+c3910U+c3A10U+c3B10U+c3C10U+c3D10U+c3E10U+c3F10U;
assign A310U=(C310U>=0)?1:0;

assign P410U=A310U;

ninexnine_unit ninexnine_unit_7584(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3011U)
);

ninexnine_unit ninexnine_unit_7585(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3111U)
);

ninexnine_unit ninexnine_unit_7586(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3211U)
);

ninexnine_unit ninexnine_unit_7587(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3311U)
);

ninexnine_unit ninexnine_unit_7588(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3411U)
);

ninexnine_unit ninexnine_unit_7589(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3511U)
);

ninexnine_unit ninexnine_unit_7590(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3611U)
);

ninexnine_unit ninexnine_unit_7591(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3711U)
);

ninexnine_unit ninexnine_unit_7592(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3811U)
);

ninexnine_unit ninexnine_unit_7593(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3911U)
);

ninexnine_unit ninexnine_unit_7594(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A11U)
);

ninexnine_unit ninexnine_unit_7595(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B11U)
);

ninexnine_unit ninexnine_unit_7596(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C11U)
);

ninexnine_unit ninexnine_unit_7597(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D11U)
);

ninexnine_unit ninexnine_unit_7598(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E11U)
);

ninexnine_unit ninexnine_unit_7599(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F11U)
);

assign C311U=c3011U+c3111U+c3211U+c3311U+c3411U+c3511U+c3611U+c3711U+c3811U+c3911U+c3A11U+c3B11U+c3C11U+c3D11U+c3E11U+c3F11U;
assign A311U=(C311U>=0)?1:0;

assign P411U=A311U;

ninexnine_unit ninexnine_unit_7600(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3012U)
);

ninexnine_unit ninexnine_unit_7601(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3112U)
);

ninexnine_unit ninexnine_unit_7602(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3212U)
);

ninexnine_unit ninexnine_unit_7603(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3312U)
);

ninexnine_unit ninexnine_unit_7604(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3412U)
);

ninexnine_unit ninexnine_unit_7605(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3512U)
);

ninexnine_unit ninexnine_unit_7606(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3612U)
);

ninexnine_unit ninexnine_unit_7607(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3712U)
);

ninexnine_unit ninexnine_unit_7608(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3812U)
);

ninexnine_unit ninexnine_unit_7609(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3912U)
);

ninexnine_unit ninexnine_unit_7610(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A12U)
);

ninexnine_unit ninexnine_unit_7611(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B12U)
);

ninexnine_unit ninexnine_unit_7612(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C12U)
);

ninexnine_unit ninexnine_unit_7613(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D12U)
);

ninexnine_unit ninexnine_unit_7614(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E12U)
);

ninexnine_unit ninexnine_unit_7615(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F12U)
);

assign C312U=c3012U+c3112U+c3212U+c3312U+c3412U+c3512U+c3612U+c3712U+c3812U+c3912U+c3A12U+c3B12U+c3C12U+c3D12U+c3E12U+c3F12U;
assign A312U=(C312U>=0)?1:0;

assign P412U=A312U;

ninexnine_unit ninexnine_unit_7616(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3020U)
);

ninexnine_unit ninexnine_unit_7617(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3120U)
);

ninexnine_unit ninexnine_unit_7618(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3220U)
);

ninexnine_unit ninexnine_unit_7619(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3320U)
);

ninexnine_unit ninexnine_unit_7620(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3420U)
);

ninexnine_unit ninexnine_unit_7621(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3520U)
);

ninexnine_unit ninexnine_unit_7622(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3620U)
);

ninexnine_unit ninexnine_unit_7623(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3720U)
);

ninexnine_unit ninexnine_unit_7624(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3820U)
);

ninexnine_unit ninexnine_unit_7625(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3920U)
);

ninexnine_unit ninexnine_unit_7626(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A20U)
);

ninexnine_unit ninexnine_unit_7627(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B20U)
);

ninexnine_unit ninexnine_unit_7628(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C20U)
);

ninexnine_unit ninexnine_unit_7629(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D20U)
);

ninexnine_unit ninexnine_unit_7630(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E20U)
);

ninexnine_unit ninexnine_unit_7631(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F20U)
);

assign C320U=c3020U+c3120U+c3220U+c3320U+c3420U+c3520U+c3620U+c3720U+c3820U+c3920U+c3A20U+c3B20U+c3C20U+c3D20U+c3E20U+c3F20U;
assign A320U=(C320U>=0)?1:0;

assign P420U=A320U;

ninexnine_unit ninexnine_unit_7632(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3021U)
);

ninexnine_unit ninexnine_unit_7633(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3121U)
);

ninexnine_unit ninexnine_unit_7634(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3221U)
);

ninexnine_unit ninexnine_unit_7635(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3321U)
);

ninexnine_unit ninexnine_unit_7636(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3421U)
);

ninexnine_unit ninexnine_unit_7637(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3521U)
);

ninexnine_unit ninexnine_unit_7638(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3621U)
);

ninexnine_unit ninexnine_unit_7639(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3721U)
);

ninexnine_unit ninexnine_unit_7640(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3821U)
);

ninexnine_unit ninexnine_unit_7641(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3921U)
);

ninexnine_unit ninexnine_unit_7642(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A21U)
);

ninexnine_unit ninexnine_unit_7643(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B21U)
);

ninexnine_unit ninexnine_unit_7644(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C21U)
);

ninexnine_unit ninexnine_unit_7645(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D21U)
);

ninexnine_unit ninexnine_unit_7646(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E21U)
);

ninexnine_unit ninexnine_unit_7647(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F21U)
);

assign C321U=c3021U+c3121U+c3221U+c3321U+c3421U+c3521U+c3621U+c3721U+c3821U+c3921U+c3A21U+c3B21U+c3C21U+c3D21U+c3E21U+c3F21U;
assign A321U=(C321U>=0)?1:0;

assign P421U=A321U;

ninexnine_unit ninexnine_unit_7648(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3U000),
				.b1(W3U010),
				.b2(W3U020),
				.b3(W3U100),
				.b4(W3U110),
				.b5(W3U120),
				.b6(W3U200),
				.b7(W3U210),
				.b8(W3U220),
				.c(c3022U)
);

ninexnine_unit ninexnine_unit_7649(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3U001),
				.b1(W3U011),
				.b2(W3U021),
				.b3(W3U101),
				.b4(W3U111),
				.b5(W3U121),
				.b6(W3U201),
				.b7(W3U211),
				.b8(W3U221),
				.c(c3122U)
);

ninexnine_unit ninexnine_unit_7650(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3U002),
				.b1(W3U012),
				.b2(W3U022),
				.b3(W3U102),
				.b4(W3U112),
				.b5(W3U122),
				.b6(W3U202),
				.b7(W3U212),
				.b8(W3U222),
				.c(c3222U)
);

ninexnine_unit ninexnine_unit_7651(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3U003),
				.b1(W3U013),
				.b2(W3U023),
				.b3(W3U103),
				.b4(W3U113),
				.b5(W3U123),
				.b6(W3U203),
				.b7(W3U213),
				.b8(W3U223),
				.c(c3322U)
);

ninexnine_unit ninexnine_unit_7652(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3U004),
				.b1(W3U014),
				.b2(W3U024),
				.b3(W3U104),
				.b4(W3U114),
				.b5(W3U124),
				.b6(W3U204),
				.b7(W3U214),
				.b8(W3U224),
				.c(c3422U)
);

ninexnine_unit ninexnine_unit_7653(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3U005),
				.b1(W3U015),
				.b2(W3U025),
				.b3(W3U105),
				.b4(W3U115),
				.b5(W3U125),
				.b6(W3U205),
				.b7(W3U215),
				.b8(W3U225),
				.c(c3522U)
);

ninexnine_unit ninexnine_unit_7654(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3U006),
				.b1(W3U016),
				.b2(W3U026),
				.b3(W3U106),
				.b4(W3U116),
				.b5(W3U126),
				.b6(W3U206),
				.b7(W3U216),
				.b8(W3U226),
				.c(c3622U)
);

ninexnine_unit ninexnine_unit_7655(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3U007),
				.b1(W3U017),
				.b2(W3U027),
				.b3(W3U107),
				.b4(W3U117),
				.b5(W3U127),
				.b6(W3U207),
				.b7(W3U217),
				.b8(W3U227),
				.c(c3722U)
);

ninexnine_unit ninexnine_unit_7656(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3U008),
				.b1(W3U018),
				.b2(W3U028),
				.b3(W3U108),
				.b4(W3U118),
				.b5(W3U128),
				.b6(W3U208),
				.b7(W3U218),
				.b8(W3U228),
				.c(c3822U)
);

ninexnine_unit ninexnine_unit_7657(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3U009),
				.b1(W3U019),
				.b2(W3U029),
				.b3(W3U109),
				.b4(W3U119),
				.b5(W3U129),
				.b6(W3U209),
				.b7(W3U219),
				.b8(W3U229),
				.c(c3922U)
);

ninexnine_unit ninexnine_unit_7658(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3U00A),
				.b1(W3U01A),
				.b2(W3U02A),
				.b3(W3U10A),
				.b4(W3U11A),
				.b5(W3U12A),
				.b6(W3U20A),
				.b7(W3U21A),
				.b8(W3U22A),
				.c(c3A22U)
);

ninexnine_unit ninexnine_unit_7659(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3U00B),
				.b1(W3U01B),
				.b2(W3U02B),
				.b3(W3U10B),
				.b4(W3U11B),
				.b5(W3U12B),
				.b6(W3U20B),
				.b7(W3U21B),
				.b8(W3U22B),
				.c(c3B22U)
);

ninexnine_unit ninexnine_unit_7660(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3U00C),
				.b1(W3U01C),
				.b2(W3U02C),
				.b3(W3U10C),
				.b4(W3U11C),
				.b5(W3U12C),
				.b6(W3U20C),
				.b7(W3U21C),
				.b8(W3U22C),
				.c(c3C22U)
);

ninexnine_unit ninexnine_unit_7661(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3U00D),
				.b1(W3U01D),
				.b2(W3U02D),
				.b3(W3U10D),
				.b4(W3U11D),
				.b5(W3U12D),
				.b6(W3U20D),
				.b7(W3U21D),
				.b8(W3U22D),
				.c(c3D22U)
);

ninexnine_unit ninexnine_unit_7662(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3U00E),
				.b1(W3U01E),
				.b2(W3U02E),
				.b3(W3U10E),
				.b4(W3U11E),
				.b5(W3U12E),
				.b6(W3U20E),
				.b7(W3U21E),
				.b8(W3U22E),
				.c(c3E22U)
);

ninexnine_unit ninexnine_unit_7663(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3U00F),
				.b1(W3U01F),
				.b2(W3U02F),
				.b3(W3U10F),
				.b4(W3U11F),
				.b5(W3U12F),
				.b6(W3U20F),
				.b7(W3U21F),
				.b8(W3U22F),
				.c(c3F22U)
);

assign C322U=c3022U+c3122U+c3222U+c3322U+c3422U+c3522U+c3622U+c3722U+c3822U+c3922U+c3A22U+c3B22U+c3C22U+c3D22U+c3E22U+c3F22U;
assign A322U=(C322U>=0)?1:0;

assign P422U=A322U;

ninexnine_unit ninexnine_unit_7664(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3000V)
);

ninexnine_unit ninexnine_unit_7665(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3100V)
);

ninexnine_unit ninexnine_unit_7666(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3200V)
);

ninexnine_unit ninexnine_unit_7667(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3300V)
);

ninexnine_unit ninexnine_unit_7668(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3400V)
);

ninexnine_unit ninexnine_unit_7669(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3500V)
);

ninexnine_unit ninexnine_unit_7670(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3600V)
);

ninexnine_unit ninexnine_unit_7671(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3700V)
);

ninexnine_unit ninexnine_unit_7672(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3800V)
);

ninexnine_unit ninexnine_unit_7673(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3900V)
);

ninexnine_unit ninexnine_unit_7674(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A00V)
);

ninexnine_unit ninexnine_unit_7675(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B00V)
);

ninexnine_unit ninexnine_unit_7676(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C00V)
);

ninexnine_unit ninexnine_unit_7677(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D00V)
);

ninexnine_unit ninexnine_unit_7678(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E00V)
);

ninexnine_unit ninexnine_unit_7679(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F00V)
);

assign C300V=c3000V+c3100V+c3200V+c3300V+c3400V+c3500V+c3600V+c3700V+c3800V+c3900V+c3A00V+c3B00V+c3C00V+c3D00V+c3E00V+c3F00V;
assign A300V=(C300V>=0)?1:0;

assign P400V=A300V;

ninexnine_unit ninexnine_unit_7680(
				.clk(clk),
				.rstn(rstn),
				.a0(P3010),
				.a1(P3020),
				.a2(P3030),
				.a3(P3110),
				.a4(P3120),
				.a5(P3130),
				.a6(P3210),
				.a7(P3220),
				.a8(P3230),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3001V)
);

ninexnine_unit ninexnine_unit_7681(
				.clk(clk),
				.rstn(rstn),
				.a0(P3011),
				.a1(P3021),
				.a2(P3031),
				.a3(P3111),
				.a4(P3121),
				.a5(P3131),
				.a6(P3211),
				.a7(P3221),
				.a8(P3231),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3101V)
);

ninexnine_unit ninexnine_unit_7682(
				.clk(clk),
				.rstn(rstn),
				.a0(P3012),
				.a1(P3022),
				.a2(P3032),
				.a3(P3112),
				.a4(P3122),
				.a5(P3132),
				.a6(P3212),
				.a7(P3222),
				.a8(P3232),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3201V)
);

ninexnine_unit ninexnine_unit_7683(
				.clk(clk),
				.rstn(rstn),
				.a0(P3013),
				.a1(P3023),
				.a2(P3033),
				.a3(P3113),
				.a4(P3123),
				.a5(P3133),
				.a6(P3213),
				.a7(P3223),
				.a8(P3233),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3301V)
);

ninexnine_unit ninexnine_unit_7684(
				.clk(clk),
				.rstn(rstn),
				.a0(P3014),
				.a1(P3024),
				.a2(P3034),
				.a3(P3114),
				.a4(P3124),
				.a5(P3134),
				.a6(P3214),
				.a7(P3224),
				.a8(P3234),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3401V)
);

ninexnine_unit ninexnine_unit_7685(
				.clk(clk),
				.rstn(rstn),
				.a0(P3015),
				.a1(P3025),
				.a2(P3035),
				.a3(P3115),
				.a4(P3125),
				.a5(P3135),
				.a6(P3215),
				.a7(P3225),
				.a8(P3235),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3501V)
);

ninexnine_unit ninexnine_unit_7686(
				.clk(clk),
				.rstn(rstn),
				.a0(P3016),
				.a1(P3026),
				.a2(P3036),
				.a3(P3116),
				.a4(P3126),
				.a5(P3136),
				.a6(P3216),
				.a7(P3226),
				.a8(P3236),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3601V)
);

ninexnine_unit ninexnine_unit_7687(
				.clk(clk),
				.rstn(rstn),
				.a0(P3017),
				.a1(P3027),
				.a2(P3037),
				.a3(P3117),
				.a4(P3127),
				.a5(P3137),
				.a6(P3217),
				.a7(P3227),
				.a8(P3237),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3701V)
);

ninexnine_unit ninexnine_unit_7688(
				.clk(clk),
				.rstn(rstn),
				.a0(P3018),
				.a1(P3028),
				.a2(P3038),
				.a3(P3118),
				.a4(P3128),
				.a5(P3138),
				.a6(P3218),
				.a7(P3228),
				.a8(P3238),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3801V)
);

ninexnine_unit ninexnine_unit_7689(
				.clk(clk),
				.rstn(rstn),
				.a0(P3019),
				.a1(P3029),
				.a2(P3039),
				.a3(P3119),
				.a4(P3129),
				.a5(P3139),
				.a6(P3219),
				.a7(P3229),
				.a8(P3239),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3901V)
);

ninexnine_unit ninexnine_unit_7690(
				.clk(clk),
				.rstn(rstn),
				.a0(P301A),
				.a1(P302A),
				.a2(P303A),
				.a3(P311A),
				.a4(P312A),
				.a5(P313A),
				.a6(P321A),
				.a7(P322A),
				.a8(P323A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A01V)
);

ninexnine_unit ninexnine_unit_7691(
				.clk(clk),
				.rstn(rstn),
				.a0(P301B),
				.a1(P302B),
				.a2(P303B),
				.a3(P311B),
				.a4(P312B),
				.a5(P313B),
				.a6(P321B),
				.a7(P322B),
				.a8(P323B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B01V)
);

ninexnine_unit ninexnine_unit_7692(
				.clk(clk),
				.rstn(rstn),
				.a0(P301C),
				.a1(P302C),
				.a2(P303C),
				.a3(P311C),
				.a4(P312C),
				.a5(P313C),
				.a6(P321C),
				.a7(P322C),
				.a8(P323C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C01V)
);

ninexnine_unit ninexnine_unit_7693(
				.clk(clk),
				.rstn(rstn),
				.a0(P301D),
				.a1(P302D),
				.a2(P303D),
				.a3(P311D),
				.a4(P312D),
				.a5(P313D),
				.a6(P321D),
				.a7(P322D),
				.a8(P323D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D01V)
);

ninexnine_unit ninexnine_unit_7694(
				.clk(clk),
				.rstn(rstn),
				.a0(P301E),
				.a1(P302E),
				.a2(P303E),
				.a3(P311E),
				.a4(P312E),
				.a5(P313E),
				.a6(P321E),
				.a7(P322E),
				.a8(P323E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E01V)
);

ninexnine_unit ninexnine_unit_7695(
				.clk(clk),
				.rstn(rstn),
				.a0(P301F),
				.a1(P302F),
				.a2(P303F),
				.a3(P311F),
				.a4(P312F),
				.a5(P313F),
				.a6(P321F),
				.a7(P322F),
				.a8(P323F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F01V)
);

assign C301V=c3001V+c3101V+c3201V+c3301V+c3401V+c3501V+c3601V+c3701V+c3801V+c3901V+c3A01V+c3B01V+c3C01V+c3D01V+c3E01V+c3F01V;
assign A301V=(C301V>=0)?1:0;

assign P401V=A301V;

ninexnine_unit ninexnine_unit_7696(
				.clk(clk),
				.rstn(rstn),
				.a0(P3020),
				.a1(P3030),
				.a2(P3040),
				.a3(P3120),
				.a4(P3130),
				.a5(P3140),
				.a6(P3220),
				.a7(P3230),
				.a8(P3240),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3002V)
);

ninexnine_unit ninexnine_unit_7697(
				.clk(clk),
				.rstn(rstn),
				.a0(P3021),
				.a1(P3031),
				.a2(P3041),
				.a3(P3121),
				.a4(P3131),
				.a5(P3141),
				.a6(P3221),
				.a7(P3231),
				.a8(P3241),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3102V)
);

ninexnine_unit ninexnine_unit_7698(
				.clk(clk),
				.rstn(rstn),
				.a0(P3022),
				.a1(P3032),
				.a2(P3042),
				.a3(P3122),
				.a4(P3132),
				.a5(P3142),
				.a6(P3222),
				.a7(P3232),
				.a8(P3242),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3202V)
);

ninexnine_unit ninexnine_unit_7699(
				.clk(clk),
				.rstn(rstn),
				.a0(P3023),
				.a1(P3033),
				.a2(P3043),
				.a3(P3123),
				.a4(P3133),
				.a5(P3143),
				.a6(P3223),
				.a7(P3233),
				.a8(P3243),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3302V)
);

ninexnine_unit ninexnine_unit_7700(
				.clk(clk),
				.rstn(rstn),
				.a0(P3024),
				.a1(P3034),
				.a2(P3044),
				.a3(P3124),
				.a4(P3134),
				.a5(P3144),
				.a6(P3224),
				.a7(P3234),
				.a8(P3244),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3402V)
);

ninexnine_unit ninexnine_unit_7701(
				.clk(clk),
				.rstn(rstn),
				.a0(P3025),
				.a1(P3035),
				.a2(P3045),
				.a3(P3125),
				.a4(P3135),
				.a5(P3145),
				.a6(P3225),
				.a7(P3235),
				.a8(P3245),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3502V)
);

ninexnine_unit ninexnine_unit_7702(
				.clk(clk),
				.rstn(rstn),
				.a0(P3026),
				.a1(P3036),
				.a2(P3046),
				.a3(P3126),
				.a4(P3136),
				.a5(P3146),
				.a6(P3226),
				.a7(P3236),
				.a8(P3246),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3602V)
);

ninexnine_unit ninexnine_unit_7703(
				.clk(clk),
				.rstn(rstn),
				.a0(P3027),
				.a1(P3037),
				.a2(P3047),
				.a3(P3127),
				.a4(P3137),
				.a5(P3147),
				.a6(P3227),
				.a7(P3237),
				.a8(P3247),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3702V)
);

ninexnine_unit ninexnine_unit_7704(
				.clk(clk),
				.rstn(rstn),
				.a0(P3028),
				.a1(P3038),
				.a2(P3048),
				.a3(P3128),
				.a4(P3138),
				.a5(P3148),
				.a6(P3228),
				.a7(P3238),
				.a8(P3248),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3802V)
);

ninexnine_unit ninexnine_unit_7705(
				.clk(clk),
				.rstn(rstn),
				.a0(P3029),
				.a1(P3039),
				.a2(P3049),
				.a3(P3129),
				.a4(P3139),
				.a5(P3149),
				.a6(P3229),
				.a7(P3239),
				.a8(P3249),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3902V)
);

ninexnine_unit ninexnine_unit_7706(
				.clk(clk),
				.rstn(rstn),
				.a0(P302A),
				.a1(P303A),
				.a2(P304A),
				.a3(P312A),
				.a4(P313A),
				.a5(P314A),
				.a6(P322A),
				.a7(P323A),
				.a8(P324A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A02V)
);

ninexnine_unit ninexnine_unit_7707(
				.clk(clk),
				.rstn(rstn),
				.a0(P302B),
				.a1(P303B),
				.a2(P304B),
				.a3(P312B),
				.a4(P313B),
				.a5(P314B),
				.a6(P322B),
				.a7(P323B),
				.a8(P324B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B02V)
);

ninexnine_unit ninexnine_unit_7708(
				.clk(clk),
				.rstn(rstn),
				.a0(P302C),
				.a1(P303C),
				.a2(P304C),
				.a3(P312C),
				.a4(P313C),
				.a5(P314C),
				.a6(P322C),
				.a7(P323C),
				.a8(P324C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C02V)
);

ninexnine_unit ninexnine_unit_7709(
				.clk(clk),
				.rstn(rstn),
				.a0(P302D),
				.a1(P303D),
				.a2(P304D),
				.a3(P312D),
				.a4(P313D),
				.a5(P314D),
				.a6(P322D),
				.a7(P323D),
				.a8(P324D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D02V)
);

ninexnine_unit ninexnine_unit_7710(
				.clk(clk),
				.rstn(rstn),
				.a0(P302E),
				.a1(P303E),
				.a2(P304E),
				.a3(P312E),
				.a4(P313E),
				.a5(P314E),
				.a6(P322E),
				.a7(P323E),
				.a8(P324E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E02V)
);

ninexnine_unit ninexnine_unit_7711(
				.clk(clk),
				.rstn(rstn),
				.a0(P302F),
				.a1(P303F),
				.a2(P304F),
				.a3(P312F),
				.a4(P313F),
				.a5(P314F),
				.a6(P322F),
				.a7(P323F),
				.a8(P324F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F02V)
);

assign C302V=c3002V+c3102V+c3202V+c3302V+c3402V+c3502V+c3602V+c3702V+c3802V+c3902V+c3A02V+c3B02V+c3C02V+c3D02V+c3E02V+c3F02V;
assign A302V=(C302V>=0)?1:0;

assign P402V=A302V;

ninexnine_unit ninexnine_unit_7712(
				.clk(clk),
				.rstn(rstn),
				.a0(P3100),
				.a1(P3110),
				.a2(P3120),
				.a3(P3200),
				.a4(P3210),
				.a5(P3220),
				.a6(P3300),
				.a7(P3310),
				.a8(P3320),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3010V)
);

ninexnine_unit ninexnine_unit_7713(
				.clk(clk),
				.rstn(rstn),
				.a0(P3101),
				.a1(P3111),
				.a2(P3121),
				.a3(P3201),
				.a4(P3211),
				.a5(P3221),
				.a6(P3301),
				.a7(P3311),
				.a8(P3321),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3110V)
);

ninexnine_unit ninexnine_unit_7714(
				.clk(clk),
				.rstn(rstn),
				.a0(P3102),
				.a1(P3112),
				.a2(P3122),
				.a3(P3202),
				.a4(P3212),
				.a5(P3222),
				.a6(P3302),
				.a7(P3312),
				.a8(P3322),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3210V)
);

ninexnine_unit ninexnine_unit_7715(
				.clk(clk),
				.rstn(rstn),
				.a0(P3103),
				.a1(P3113),
				.a2(P3123),
				.a3(P3203),
				.a4(P3213),
				.a5(P3223),
				.a6(P3303),
				.a7(P3313),
				.a8(P3323),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3310V)
);

ninexnine_unit ninexnine_unit_7716(
				.clk(clk),
				.rstn(rstn),
				.a0(P3104),
				.a1(P3114),
				.a2(P3124),
				.a3(P3204),
				.a4(P3214),
				.a5(P3224),
				.a6(P3304),
				.a7(P3314),
				.a8(P3324),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3410V)
);

ninexnine_unit ninexnine_unit_7717(
				.clk(clk),
				.rstn(rstn),
				.a0(P3105),
				.a1(P3115),
				.a2(P3125),
				.a3(P3205),
				.a4(P3215),
				.a5(P3225),
				.a6(P3305),
				.a7(P3315),
				.a8(P3325),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3510V)
);

ninexnine_unit ninexnine_unit_7718(
				.clk(clk),
				.rstn(rstn),
				.a0(P3106),
				.a1(P3116),
				.a2(P3126),
				.a3(P3206),
				.a4(P3216),
				.a5(P3226),
				.a6(P3306),
				.a7(P3316),
				.a8(P3326),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3610V)
);

ninexnine_unit ninexnine_unit_7719(
				.clk(clk),
				.rstn(rstn),
				.a0(P3107),
				.a1(P3117),
				.a2(P3127),
				.a3(P3207),
				.a4(P3217),
				.a5(P3227),
				.a6(P3307),
				.a7(P3317),
				.a8(P3327),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3710V)
);

ninexnine_unit ninexnine_unit_7720(
				.clk(clk),
				.rstn(rstn),
				.a0(P3108),
				.a1(P3118),
				.a2(P3128),
				.a3(P3208),
				.a4(P3218),
				.a5(P3228),
				.a6(P3308),
				.a7(P3318),
				.a8(P3328),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3810V)
);

ninexnine_unit ninexnine_unit_7721(
				.clk(clk),
				.rstn(rstn),
				.a0(P3109),
				.a1(P3119),
				.a2(P3129),
				.a3(P3209),
				.a4(P3219),
				.a5(P3229),
				.a6(P3309),
				.a7(P3319),
				.a8(P3329),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3910V)
);

ninexnine_unit ninexnine_unit_7722(
				.clk(clk),
				.rstn(rstn),
				.a0(P310A),
				.a1(P311A),
				.a2(P312A),
				.a3(P320A),
				.a4(P321A),
				.a5(P322A),
				.a6(P330A),
				.a7(P331A),
				.a8(P332A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A10V)
);

ninexnine_unit ninexnine_unit_7723(
				.clk(clk),
				.rstn(rstn),
				.a0(P310B),
				.a1(P311B),
				.a2(P312B),
				.a3(P320B),
				.a4(P321B),
				.a5(P322B),
				.a6(P330B),
				.a7(P331B),
				.a8(P332B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B10V)
);

ninexnine_unit ninexnine_unit_7724(
				.clk(clk),
				.rstn(rstn),
				.a0(P310C),
				.a1(P311C),
				.a2(P312C),
				.a3(P320C),
				.a4(P321C),
				.a5(P322C),
				.a6(P330C),
				.a7(P331C),
				.a8(P332C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C10V)
);

ninexnine_unit ninexnine_unit_7725(
				.clk(clk),
				.rstn(rstn),
				.a0(P310D),
				.a1(P311D),
				.a2(P312D),
				.a3(P320D),
				.a4(P321D),
				.a5(P322D),
				.a6(P330D),
				.a7(P331D),
				.a8(P332D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D10V)
);

ninexnine_unit ninexnine_unit_7726(
				.clk(clk),
				.rstn(rstn),
				.a0(P310E),
				.a1(P311E),
				.a2(P312E),
				.a3(P320E),
				.a4(P321E),
				.a5(P322E),
				.a6(P330E),
				.a7(P331E),
				.a8(P332E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E10V)
);

ninexnine_unit ninexnine_unit_7727(
				.clk(clk),
				.rstn(rstn),
				.a0(P310F),
				.a1(P311F),
				.a2(P312F),
				.a3(P320F),
				.a4(P321F),
				.a5(P322F),
				.a6(P330F),
				.a7(P331F),
				.a8(P332F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F10V)
);

assign C310V=c3010V+c3110V+c3210V+c3310V+c3410V+c3510V+c3610V+c3710V+c3810V+c3910V+c3A10V+c3B10V+c3C10V+c3D10V+c3E10V+c3F10V;
assign A310V=(C310V>=0)?1:0;

assign P410V=A310V;

ninexnine_unit ninexnine_unit_7728(
				.clk(clk),
				.rstn(rstn),
				.a0(P3110),
				.a1(P3120),
				.a2(P3130),
				.a3(P3210),
				.a4(P3220),
				.a5(P3230),
				.a6(P3310),
				.a7(P3320),
				.a8(P3330),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3011V)
);

ninexnine_unit ninexnine_unit_7729(
				.clk(clk),
				.rstn(rstn),
				.a0(P3111),
				.a1(P3121),
				.a2(P3131),
				.a3(P3211),
				.a4(P3221),
				.a5(P3231),
				.a6(P3311),
				.a7(P3321),
				.a8(P3331),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3111V)
);

ninexnine_unit ninexnine_unit_7730(
				.clk(clk),
				.rstn(rstn),
				.a0(P3112),
				.a1(P3122),
				.a2(P3132),
				.a3(P3212),
				.a4(P3222),
				.a5(P3232),
				.a6(P3312),
				.a7(P3322),
				.a8(P3332),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3211V)
);

ninexnine_unit ninexnine_unit_7731(
				.clk(clk),
				.rstn(rstn),
				.a0(P3113),
				.a1(P3123),
				.a2(P3133),
				.a3(P3213),
				.a4(P3223),
				.a5(P3233),
				.a6(P3313),
				.a7(P3323),
				.a8(P3333),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3311V)
);

ninexnine_unit ninexnine_unit_7732(
				.clk(clk),
				.rstn(rstn),
				.a0(P3114),
				.a1(P3124),
				.a2(P3134),
				.a3(P3214),
				.a4(P3224),
				.a5(P3234),
				.a6(P3314),
				.a7(P3324),
				.a8(P3334),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3411V)
);

ninexnine_unit ninexnine_unit_7733(
				.clk(clk),
				.rstn(rstn),
				.a0(P3115),
				.a1(P3125),
				.a2(P3135),
				.a3(P3215),
				.a4(P3225),
				.a5(P3235),
				.a6(P3315),
				.a7(P3325),
				.a8(P3335),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3511V)
);

ninexnine_unit ninexnine_unit_7734(
				.clk(clk),
				.rstn(rstn),
				.a0(P3116),
				.a1(P3126),
				.a2(P3136),
				.a3(P3216),
				.a4(P3226),
				.a5(P3236),
				.a6(P3316),
				.a7(P3326),
				.a8(P3336),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3611V)
);

ninexnine_unit ninexnine_unit_7735(
				.clk(clk),
				.rstn(rstn),
				.a0(P3117),
				.a1(P3127),
				.a2(P3137),
				.a3(P3217),
				.a4(P3227),
				.a5(P3237),
				.a6(P3317),
				.a7(P3327),
				.a8(P3337),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3711V)
);

ninexnine_unit ninexnine_unit_7736(
				.clk(clk),
				.rstn(rstn),
				.a0(P3118),
				.a1(P3128),
				.a2(P3138),
				.a3(P3218),
				.a4(P3228),
				.a5(P3238),
				.a6(P3318),
				.a7(P3328),
				.a8(P3338),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3811V)
);

ninexnine_unit ninexnine_unit_7737(
				.clk(clk),
				.rstn(rstn),
				.a0(P3119),
				.a1(P3129),
				.a2(P3139),
				.a3(P3219),
				.a4(P3229),
				.a5(P3239),
				.a6(P3319),
				.a7(P3329),
				.a8(P3339),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3911V)
);

ninexnine_unit ninexnine_unit_7738(
				.clk(clk),
				.rstn(rstn),
				.a0(P311A),
				.a1(P312A),
				.a2(P313A),
				.a3(P321A),
				.a4(P322A),
				.a5(P323A),
				.a6(P331A),
				.a7(P332A),
				.a8(P333A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A11V)
);

ninexnine_unit ninexnine_unit_7739(
				.clk(clk),
				.rstn(rstn),
				.a0(P311B),
				.a1(P312B),
				.a2(P313B),
				.a3(P321B),
				.a4(P322B),
				.a5(P323B),
				.a6(P331B),
				.a7(P332B),
				.a8(P333B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B11V)
);

ninexnine_unit ninexnine_unit_7740(
				.clk(clk),
				.rstn(rstn),
				.a0(P311C),
				.a1(P312C),
				.a2(P313C),
				.a3(P321C),
				.a4(P322C),
				.a5(P323C),
				.a6(P331C),
				.a7(P332C),
				.a8(P333C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C11V)
);

ninexnine_unit ninexnine_unit_7741(
				.clk(clk),
				.rstn(rstn),
				.a0(P311D),
				.a1(P312D),
				.a2(P313D),
				.a3(P321D),
				.a4(P322D),
				.a5(P323D),
				.a6(P331D),
				.a7(P332D),
				.a8(P333D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D11V)
);

ninexnine_unit ninexnine_unit_7742(
				.clk(clk),
				.rstn(rstn),
				.a0(P311E),
				.a1(P312E),
				.a2(P313E),
				.a3(P321E),
				.a4(P322E),
				.a5(P323E),
				.a6(P331E),
				.a7(P332E),
				.a8(P333E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E11V)
);

ninexnine_unit ninexnine_unit_7743(
				.clk(clk),
				.rstn(rstn),
				.a0(P311F),
				.a1(P312F),
				.a2(P313F),
				.a3(P321F),
				.a4(P322F),
				.a5(P323F),
				.a6(P331F),
				.a7(P332F),
				.a8(P333F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F11V)
);

assign C311V=c3011V+c3111V+c3211V+c3311V+c3411V+c3511V+c3611V+c3711V+c3811V+c3911V+c3A11V+c3B11V+c3C11V+c3D11V+c3E11V+c3F11V;
assign A311V=(C311V>=0)?1:0;

assign P411V=A311V;

ninexnine_unit ninexnine_unit_7744(
				.clk(clk),
				.rstn(rstn),
				.a0(P3120),
				.a1(P3130),
				.a2(P3140),
				.a3(P3220),
				.a4(P3230),
				.a5(P3240),
				.a6(P3320),
				.a7(P3330),
				.a8(P3340),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3012V)
);

ninexnine_unit ninexnine_unit_7745(
				.clk(clk),
				.rstn(rstn),
				.a0(P3121),
				.a1(P3131),
				.a2(P3141),
				.a3(P3221),
				.a4(P3231),
				.a5(P3241),
				.a6(P3321),
				.a7(P3331),
				.a8(P3341),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3112V)
);

ninexnine_unit ninexnine_unit_7746(
				.clk(clk),
				.rstn(rstn),
				.a0(P3122),
				.a1(P3132),
				.a2(P3142),
				.a3(P3222),
				.a4(P3232),
				.a5(P3242),
				.a6(P3322),
				.a7(P3332),
				.a8(P3342),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3212V)
);

ninexnine_unit ninexnine_unit_7747(
				.clk(clk),
				.rstn(rstn),
				.a0(P3123),
				.a1(P3133),
				.a2(P3143),
				.a3(P3223),
				.a4(P3233),
				.a5(P3243),
				.a6(P3323),
				.a7(P3333),
				.a8(P3343),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3312V)
);

ninexnine_unit ninexnine_unit_7748(
				.clk(clk),
				.rstn(rstn),
				.a0(P3124),
				.a1(P3134),
				.a2(P3144),
				.a3(P3224),
				.a4(P3234),
				.a5(P3244),
				.a6(P3324),
				.a7(P3334),
				.a8(P3344),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3412V)
);

ninexnine_unit ninexnine_unit_7749(
				.clk(clk),
				.rstn(rstn),
				.a0(P3125),
				.a1(P3135),
				.a2(P3145),
				.a3(P3225),
				.a4(P3235),
				.a5(P3245),
				.a6(P3325),
				.a7(P3335),
				.a8(P3345),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3512V)
);

ninexnine_unit ninexnine_unit_7750(
				.clk(clk),
				.rstn(rstn),
				.a0(P3126),
				.a1(P3136),
				.a2(P3146),
				.a3(P3226),
				.a4(P3236),
				.a5(P3246),
				.a6(P3326),
				.a7(P3336),
				.a8(P3346),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3612V)
);

ninexnine_unit ninexnine_unit_7751(
				.clk(clk),
				.rstn(rstn),
				.a0(P3127),
				.a1(P3137),
				.a2(P3147),
				.a3(P3227),
				.a4(P3237),
				.a5(P3247),
				.a6(P3327),
				.a7(P3337),
				.a8(P3347),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3712V)
);

ninexnine_unit ninexnine_unit_7752(
				.clk(clk),
				.rstn(rstn),
				.a0(P3128),
				.a1(P3138),
				.a2(P3148),
				.a3(P3228),
				.a4(P3238),
				.a5(P3248),
				.a6(P3328),
				.a7(P3338),
				.a8(P3348),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3812V)
);

ninexnine_unit ninexnine_unit_7753(
				.clk(clk),
				.rstn(rstn),
				.a0(P3129),
				.a1(P3139),
				.a2(P3149),
				.a3(P3229),
				.a4(P3239),
				.a5(P3249),
				.a6(P3329),
				.a7(P3339),
				.a8(P3349),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3912V)
);

ninexnine_unit ninexnine_unit_7754(
				.clk(clk),
				.rstn(rstn),
				.a0(P312A),
				.a1(P313A),
				.a2(P314A),
				.a3(P322A),
				.a4(P323A),
				.a5(P324A),
				.a6(P332A),
				.a7(P333A),
				.a8(P334A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A12V)
);

ninexnine_unit ninexnine_unit_7755(
				.clk(clk),
				.rstn(rstn),
				.a0(P312B),
				.a1(P313B),
				.a2(P314B),
				.a3(P322B),
				.a4(P323B),
				.a5(P324B),
				.a6(P332B),
				.a7(P333B),
				.a8(P334B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B12V)
);

ninexnine_unit ninexnine_unit_7756(
				.clk(clk),
				.rstn(rstn),
				.a0(P312C),
				.a1(P313C),
				.a2(P314C),
				.a3(P322C),
				.a4(P323C),
				.a5(P324C),
				.a6(P332C),
				.a7(P333C),
				.a8(P334C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C12V)
);

ninexnine_unit ninexnine_unit_7757(
				.clk(clk),
				.rstn(rstn),
				.a0(P312D),
				.a1(P313D),
				.a2(P314D),
				.a3(P322D),
				.a4(P323D),
				.a5(P324D),
				.a6(P332D),
				.a7(P333D),
				.a8(P334D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D12V)
);

ninexnine_unit ninexnine_unit_7758(
				.clk(clk),
				.rstn(rstn),
				.a0(P312E),
				.a1(P313E),
				.a2(P314E),
				.a3(P322E),
				.a4(P323E),
				.a5(P324E),
				.a6(P332E),
				.a7(P333E),
				.a8(P334E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E12V)
);

ninexnine_unit ninexnine_unit_7759(
				.clk(clk),
				.rstn(rstn),
				.a0(P312F),
				.a1(P313F),
				.a2(P314F),
				.a3(P322F),
				.a4(P323F),
				.a5(P324F),
				.a6(P332F),
				.a7(P333F),
				.a8(P334F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F12V)
);

assign C312V=c3012V+c3112V+c3212V+c3312V+c3412V+c3512V+c3612V+c3712V+c3812V+c3912V+c3A12V+c3B12V+c3C12V+c3D12V+c3E12V+c3F12V;
assign A312V=(C312V>=0)?1:0;

assign P412V=A312V;

ninexnine_unit ninexnine_unit_7760(
				.clk(clk),
				.rstn(rstn),
				.a0(P3200),
				.a1(P3210),
				.a2(P3220),
				.a3(P3300),
				.a4(P3310),
				.a5(P3320),
				.a6(P3400),
				.a7(P3410),
				.a8(P3420),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3020V)
);

ninexnine_unit ninexnine_unit_7761(
				.clk(clk),
				.rstn(rstn),
				.a0(P3201),
				.a1(P3211),
				.a2(P3221),
				.a3(P3301),
				.a4(P3311),
				.a5(P3321),
				.a6(P3401),
				.a7(P3411),
				.a8(P3421),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3120V)
);

ninexnine_unit ninexnine_unit_7762(
				.clk(clk),
				.rstn(rstn),
				.a0(P3202),
				.a1(P3212),
				.a2(P3222),
				.a3(P3302),
				.a4(P3312),
				.a5(P3322),
				.a6(P3402),
				.a7(P3412),
				.a8(P3422),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3220V)
);

ninexnine_unit ninexnine_unit_7763(
				.clk(clk),
				.rstn(rstn),
				.a0(P3203),
				.a1(P3213),
				.a2(P3223),
				.a3(P3303),
				.a4(P3313),
				.a5(P3323),
				.a6(P3403),
				.a7(P3413),
				.a8(P3423),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3320V)
);

ninexnine_unit ninexnine_unit_7764(
				.clk(clk),
				.rstn(rstn),
				.a0(P3204),
				.a1(P3214),
				.a2(P3224),
				.a3(P3304),
				.a4(P3314),
				.a5(P3324),
				.a6(P3404),
				.a7(P3414),
				.a8(P3424),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3420V)
);

ninexnine_unit ninexnine_unit_7765(
				.clk(clk),
				.rstn(rstn),
				.a0(P3205),
				.a1(P3215),
				.a2(P3225),
				.a3(P3305),
				.a4(P3315),
				.a5(P3325),
				.a6(P3405),
				.a7(P3415),
				.a8(P3425),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3520V)
);

ninexnine_unit ninexnine_unit_7766(
				.clk(clk),
				.rstn(rstn),
				.a0(P3206),
				.a1(P3216),
				.a2(P3226),
				.a3(P3306),
				.a4(P3316),
				.a5(P3326),
				.a6(P3406),
				.a7(P3416),
				.a8(P3426),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3620V)
);

ninexnine_unit ninexnine_unit_7767(
				.clk(clk),
				.rstn(rstn),
				.a0(P3207),
				.a1(P3217),
				.a2(P3227),
				.a3(P3307),
				.a4(P3317),
				.a5(P3327),
				.a6(P3407),
				.a7(P3417),
				.a8(P3427),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3720V)
);

ninexnine_unit ninexnine_unit_7768(
				.clk(clk),
				.rstn(rstn),
				.a0(P3208),
				.a1(P3218),
				.a2(P3228),
				.a3(P3308),
				.a4(P3318),
				.a5(P3328),
				.a6(P3408),
				.a7(P3418),
				.a8(P3428),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3820V)
);

ninexnine_unit ninexnine_unit_7769(
				.clk(clk),
				.rstn(rstn),
				.a0(P3209),
				.a1(P3219),
				.a2(P3229),
				.a3(P3309),
				.a4(P3319),
				.a5(P3329),
				.a6(P3409),
				.a7(P3419),
				.a8(P3429),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3920V)
);

ninexnine_unit ninexnine_unit_7770(
				.clk(clk),
				.rstn(rstn),
				.a0(P320A),
				.a1(P321A),
				.a2(P322A),
				.a3(P330A),
				.a4(P331A),
				.a5(P332A),
				.a6(P340A),
				.a7(P341A),
				.a8(P342A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A20V)
);

ninexnine_unit ninexnine_unit_7771(
				.clk(clk),
				.rstn(rstn),
				.a0(P320B),
				.a1(P321B),
				.a2(P322B),
				.a3(P330B),
				.a4(P331B),
				.a5(P332B),
				.a6(P340B),
				.a7(P341B),
				.a8(P342B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B20V)
);

ninexnine_unit ninexnine_unit_7772(
				.clk(clk),
				.rstn(rstn),
				.a0(P320C),
				.a1(P321C),
				.a2(P322C),
				.a3(P330C),
				.a4(P331C),
				.a5(P332C),
				.a6(P340C),
				.a7(P341C),
				.a8(P342C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C20V)
);

ninexnine_unit ninexnine_unit_7773(
				.clk(clk),
				.rstn(rstn),
				.a0(P320D),
				.a1(P321D),
				.a2(P322D),
				.a3(P330D),
				.a4(P331D),
				.a5(P332D),
				.a6(P340D),
				.a7(P341D),
				.a8(P342D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D20V)
);

ninexnine_unit ninexnine_unit_7774(
				.clk(clk),
				.rstn(rstn),
				.a0(P320E),
				.a1(P321E),
				.a2(P322E),
				.a3(P330E),
				.a4(P331E),
				.a5(P332E),
				.a6(P340E),
				.a7(P341E),
				.a8(P342E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E20V)
);

ninexnine_unit ninexnine_unit_7775(
				.clk(clk),
				.rstn(rstn),
				.a0(P320F),
				.a1(P321F),
				.a2(P322F),
				.a3(P330F),
				.a4(P331F),
				.a5(P332F),
				.a6(P340F),
				.a7(P341F),
				.a8(P342F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F20V)
);

assign C320V=c3020V+c3120V+c3220V+c3320V+c3420V+c3520V+c3620V+c3720V+c3820V+c3920V+c3A20V+c3B20V+c3C20V+c3D20V+c3E20V+c3F20V;
assign A320V=(C320V>=0)?1:0;

assign P420V=A320V;

ninexnine_unit ninexnine_unit_7776(
				.clk(clk),
				.rstn(rstn),
				.a0(P3210),
				.a1(P3220),
				.a2(P3230),
				.a3(P3310),
				.a4(P3320),
				.a5(P3330),
				.a6(P3410),
				.a7(P3420),
				.a8(P3430),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3021V)
);

ninexnine_unit ninexnine_unit_7777(
				.clk(clk),
				.rstn(rstn),
				.a0(P3211),
				.a1(P3221),
				.a2(P3231),
				.a3(P3311),
				.a4(P3321),
				.a5(P3331),
				.a6(P3411),
				.a7(P3421),
				.a8(P3431),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3121V)
);

ninexnine_unit ninexnine_unit_7778(
				.clk(clk),
				.rstn(rstn),
				.a0(P3212),
				.a1(P3222),
				.a2(P3232),
				.a3(P3312),
				.a4(P3322),
				.a5(P3332),
				.a6(P3412),
				.a7(P3422),
				.a8(P3432),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3221V)
);

ninexnine_unit ninexnine_unit_7779(
				.clk(clk),
				.rstn(rstn),
				.a0(P3213),
				.a1(P3223),
				.a2(P3233),
				.a3(P3313),
				.a4(P3323),
				.a5(P3333),
				.a6(P3413),
				.a7(P3423),
				.a8(P3433),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3321V)
);

ninexnine_unit ninexnine_unit_7780(
				.clk(clk),
				.rstn(rstn),
				.a0(P3214),
				.a1(P3224),
				.a2(P3234),
				.a3(P3314),
				.a4(P3324),
				.a5(P3334),
				.a6(P3414),
				.a7(P3424),
				.a8(P3434),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3421V)
);

ninexnine_unit ninexnine_unit_7781(
				.clk(clk),
				.rstn(rstn),
				.a0(P3215),
				.a1(P3225),
				.a2(P3235),
				.a3(P3315),
				.a4(P3325),
				.a5(P3335),
				.a6(P3415),
				.a7(P3425),
				.a8(P3435),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3521V)
);

ninexnine_unit ninexnine_unit_7782(
				.clk(clk),
				.rstn(rstn),
				.a0(P3216),
				.a1(P3226),
				.a2(P3236),
				.a3(P3316),
				.a4(P3326),
				.a5(P3336),
				.a6(P3416),
				.a7(P3426),
				.a8(P3436),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3621V)
);

ninexnine_unit ninexnine_unit_7783(
				.clk(clk),
				.rstn(rstn),
				.a0(P3217),
				.a1(P3227),
				.a2(P3237),
				.a3(P3317),
				.a4(P3327),
				.a5(P3337),
				.a6(P3417),
				.a7(P3427),
				.a8(P3437),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3721V)
);

ninexnine_unit ninexnine_unit_7784(
				.clk(clk),
				.rstn(rstn),
				.a0(P3218),
				.a1(P3228),
				.a2(P3238),
				.a3(P3318),
				.a4(P3328),
				.a5(P3338),
				.a6(P3418),
				.a7(P3428),
				.a8(P3438),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3821V)
);

ninexnine_unit ninexnine_unit_7785(
				.clk(clk),
				.rstn(rstn),
				.a0(P3219),
				.a1(P3229),
				.a2(P3239),
				.a3(P3319),
				.a4(P3329),
				.a5(P3339),
				.a6(P3419),
				.a7(P3429),
				.a8(P3439),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3921V)
);

ninexnine_unit ninexnine_unit_7786(
				.clk(clk),
				.rstn(rstn),
				.a0(P321A),
				.a1(P322A),
				.a2(P323A),
				.a3(P331A),
				.a4(P332A),
				.a5(P333A),
				.a6(P341A),
				.a7(P342A),
				.a8(P343A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A21V)
);

ninexnine_unit ninexnine_unit_7787(
				.clk(clk),
				.rstn(rstn),
				.a0(P321B),
				.a1(P322B),
				.a2(P323B),
				.a3(P331B),
				.a4(P332B),
				.a5(P333B),
				.a6(P341B),
				.a7(P342B),
				.a8(P343B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B21V)
);

ninexnine_unit ninexnine_unit_7788(
				.clk(clk),
				.rstn(rstn),
				.a0(P321C),
				.a1(P322C),
				.a2(P323C),
				.a3(P331C),
				.a4(P332C),
				.a5(P333C),
				.a6(P341C),
				.a7(P342C),
				.a8(P343C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C21V)
);

ninexnine_unit ninexnine_unit_7789(
				.clk(clk),
				.rstn(rstn),
				.a0(P321D),
				.a1(P322D),
				.a2(P323D),
				.a3(P331D),
				.a4(P332D),
				.a5(P333D),
				.a6(P341D),
				.a7(P342D),
				.a8(P343D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D21V)
);

ninexnine_unit ninexnine_unit_7790(
				.clk(clk),
				.rstn(rstn),
				.a0(P321E),
				.a1(P322E),
				.a2(P323E),
				.a3(P331E),
				.a4(P332E),
				.a5(P333E),
				.a6(P341E),
				.a7(P342E),
				.a8(P343E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E21V)
);

ninexnine_unit ninexnine_unit_7791(
				.clk(clk),
				.rstn(rstn),
				.a0(P321F),
				.a1(P322F),
				.a2(P323F),
				.a3(P331F),
				.a4(P332F),
				.a5(P333F),
				.a6(P341F),
				.a7(P342F),
				.a8(P343F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F21V)
);

assign C321V=c3021V+c3121V+c3221V+c3321V+c3421V+c3521V+c3621V+c3721V+c3821V+c3921V+c3A21V+c3B21V+c3C21V+c3D21V+c3E21V+c3F21V;
assign A321V=(C321V>=0)?1:0;

assign P421V=A321V;

ninexnine_unit ninexnine_unit_7792(
				.clk(clk),
				.rstn(rstn),
				.a0(P3220),
				.a1(P3230),
				.a2(P3240),
				.a3(P3320),
				.a4(P3330),
				.a5(P3340),
				.a6(P3420),
				.a7(P3430),
				.a8(P3440),
				.b0(W3V000),
				.b1(W3V010),
				.b2(W3V020),
				.b3(W3V100),
				.b4(W3V110),
				.b5(W3V120),
				.b6(W3V200),
				.b7(W3V210),
				.b8(W3V220),
				.c(c3022V)
);

ninexnine_unit ninexnine_unit_7793(
				.clk(clk),
				.rstn(rstn),
				.a0(P3221),
				.a1(P3231),
				.a2(P3241),
				.a3(P3321),
				.a4(P3331),
				.a5(P3341),
				.a6(P3421),
				.a7(P3431),
				.a8(P3441),
				.b0(W3V001),
				.b1(W3V011),
				.b2(W3V021),
				.b3(W3V101),
				.b4(W3V111),
				.b5(W3V121),
				.b6(W3V201),
				.b7(W3V211),
				.b8(W3V221),
				.c(c3122V)
);

ninexnine_unit ninexnine_unit_7794(
				.clk(clk),
				.rstn(rstn),
				.a0(P3222),
				.a1(P3232),
				.a2(P3242),
				.a3(P3322),
				.a4(P3332),
				.a5(P3342),
				.a6(P3422),
				.a7(P3432),
				.a8(P3442),
				.b0(W3V002),
				.b1(W3V012),
				.b2(W3V022),
				.b3(W3V102),
				.b4(W3V112),
				.b5(W3V122),
				.b6(W3V202),
				.b7(W3V212),
				.b8(W3V222),
				.c(c3222V)
);

ninexnine_unit ninexnine_unit_7795(
				.clk(clk),
				.rstn(rstn),
				.a0(P3223),
				.a1(P3233),
				.a2(P3243),
				.a3(P3323),
				.a4(P3333),
				.a5(P3343),
				.a6(P3423),
				.a7(P3433),
				.a8(P3443),
				.b0(W3V003),
				.b1(W3V013),
				.b2(W3V023),
				.b3(W3V103),
				.b4(W3V113),
				.b5(W3V123),
				.b6(W3V203),
				.b7(W3V213),
				.b8(W3V223),
				.c(c3322V)
);

ninexnine_unit ninexnine_unit_7796(
				.clk(clk),
				.rstn(rstn),
				.a0(P3224),
				.a1(P3234),
				.a2(P3244),
				.a3(P3324),
				.a4(P3334),
				.a5(P3344),
				.a6(P3424),
				.a7(P3434),
				.a8(P3444),
				.b0(W3V004),
				.b1(W3V014),
				.b2(W3V024),
				.b3(W3V104),
				.b4(W3V114),
				.b5(W3V124),
				.b6(W3V204),
				.b7(W3V214),
				.b8(W3V224),
				.c(c3422V)
);

ninexnine_unit ninexnine_unit_7797(
				.clk(clk),
				.rstn(rstn),
				.a0(P3225),
				.a1(P3235),
				.a2(P3245),
				.a3(P3325),
				.a4(P3335),
				.a5(P3345),
				.a6(P3425),
				.a7(P3435),
				.a8(P3445),
				.b0(W3V005),
				.b1(W3V015),
				.b2(W3V025),
				.b3(W3V105),
				.b4(W3V115),
				.b5(W3V125),
				.b6(W3V205),
				.b7(W3V215),
				.b8(W3V225),
				.c(c3522V)
);

ninexnine_unit ninexnine_unit_7798(
				.clk(clk),
				.rstn(rstn),
				.a0(P3226),
				.a1(P3236),
				.a2(P3246),
				.a3(P3326),
				.a4(P3336),
				.a5(P3346),
				.a6(P3426),
				.a7(P3436),
				.a8(P3446),
				.b0(W3V006),
				.b1(W3V016),
				.b2(W3V026),
				.b3(W3V106),
				.b4(W3V116),
				.b5(W3V126),
				.b6(W3V206),
				.b7(W3V216),
				.b8(W3V226),
				.c(c3622V)
);

ninexnine_unit ninexnine_unit_7799(
				.clk(clk),
				.rstn(rstn),
				.a0(P3227),
				.a1(P3237),
				.a2(P3247),
				.a3(P3327),
				.a4(P3337),
				.a5(P3347),
				.a6(P3427),
				.a7(P3437),
				.a8(P3447),
				.b0(W3V007),
				.b1(W3V017),
				.b2(W3V027),
				.b3(W3V107),
				.b4(W3V117),
				.b5(W3V127),
				.b6(W3V207),
				.b7(W3V217),
				.b8(W3V227),
				.c(c3722V)
);

ninexnine_unit ninexnine_unit_7800(
				.clk(clk),
				.rstn(rstn),
				.a0(P3228),
				.a1(P3238),
				.a2(P3248),
				.a3(P3328),
				.a4(P3338),
				.a5(P3348),
				.a6(P3428),
				.a7(P3438),
				.a8(P3448),
				.b0(W3V008),
				.b1(W3V018),
				.b2(W3V028),
				.b3(W3V108),
				.b4(W3V118),
				.b5(W3V128),
				.b6(W3V208),
				.b7(W3V218),
				.b8(W3V228),
				.c(c3822V)
);

ninexnine_unit ninexnine_unit_7801(
				.clk(clk),
				.rstn(rstn),
				.a0(P3229),
				.a1(P3239),
				.a2(P3249),
				.a3(P3329),
				.a4(P3339),
				.a5(P3349),
				.a6(P3429),
				.a7(P3439),
				.a8(P3449),
				.b0(W3V009),
				.b1(W3V019),
				.b2(W3V029),
				.b3(W3V109),
				.b4(W3V119),
				.b5(W3V129),
				.b6(W3V209),
				.b7(W3V219),
				.b8(W3V229),
				.c(c3922V)
);

ninexnine_unit ninexnine_unit_7802(
				.clk(clk),
				.rstn(rstn),
				.a0(P322A),
				.a1(P323A),
				.a2(P324A),
				.a3(P332A),
				.a4(P333A),
				.a5(P334A),
				.a6(P342A),
				.a7(P343A),
				.a8(P344A),
				.b0(W3V00A),
				.b1(W3V01A),
				.b2(W3V02A),
				.b3(W3V10A),
				.b4(W3V11A),
				.b5(W3V12A),
				.b6(W3V20A),
				.b7(W3V21A),
				.b8(W3V22A),
				.c(c3A22V)
);

ninexnine_unit ninexnine_unit_7803(
				.clk(clk),
				.rstn(rstn),
				.a0(P322B),
				.a1(P323B),
				.a2(P324B),
				.a3(P332B),
				.a4(P333B),
				.a5(P334B),
				.a6(P342B),
				.a7(P343B),
				.a8(P344B),
				.b0(W3V00B),
				.b1(W3V01B),
				.b2(W3V02B),
				.b3(W3V10B),
				.b4(W3V11B),
				.b5(W3V12B),
				.b6(W3V20B),
				.b7(W3V21B),
				.b8(W3V22B),
				.c(c3B22V)
);

ninexnine_unit ninexnine_unit_7804(
				.clk(clk),
				.rstn(rstn),
				.a0(P322C),
				.a1(P323C),
				.a2(P324C),
				.a3(P332C),
				.a4(P333C),
				.a5(P334C),
				.a6(P342C),
				.a7(P343C),
				.a8(P344C),
				.b0(W3V00C),
				.b1(W3V01C),
				.b2(W3V02C),
				.b3(W3V10C),
				.b4(W3V11C),
				.b5(W3V12C),
				.b6(W3V20C),
				.b7(W3V21C),
				.b8(W3V22C),
				.c(c3C22V)
);

ninexnine_unit ninexnine_unit_7805(
				.clk(clk),
				.rstn(rstn),
				.a0(P322D),
				.a1(P323D),
				.a2(P324D),
				.a3(P332D),
				.a4(P333D),
				.a5(P334D),
				.a6(P342D),
				.a7(P343D),
				.a8(P344D),
				.b0(W3V00D),
				.b1(W3V01D),
				.b2(W3V02D),
				.b3(W3V10D),
				.b4(W3V11D),
				.b5(W3V12D),
				.b6(W3V20D),
				.b7(W3V21D),
				.b8(W3V22D),
				.c(c3D22V)
);

ninexnine_unit ninexnine_unit_7806(
				.clk(clk),
				.rstn(rstn),
				.a0(P322E),
				.a1(P323E),
				.a2(P324E),
				.a3(P332E),
				.a4(P333E),
				.a5(P334E),
				.a6(P342E),
				.a7(P343E),
				.a8(P344E),
				.b0(W3V00E),
				.b1(W3V01E),
				.b2(W3V02E),
				.b3(W3V10E),
				.b4(W3V11E),
				.b5(W3V12E),
				.b6(W3V20E),
				.b7(W3V21E),
				.b8(W3V22E),
				.c(c3E22V)
);

ninexnine_unit ninexnine_unit_7807(
				.clk(clk),
				.rstn(rstn),
				.a0(P322F),
				.a1(P323F),
				.a2(P324F),
				.a3(P332F),
				.a4(P333F),
				.a5(P334F),
				.a6(P342F),
				.a7(P343F),
				.a8(P344F),
				.b0(W3V00F),
				.b1(W3V01F),
				.b2(W3V02F),
				.b3(W3V10F),
				.b4(W3V11F),
				.b5(W3V12F),
				.b6(W3V20F),
				.b7(W3V21F),
				.b8(W3V22F),
				.c(c3F22V)
);

assign C322V=c3022V+c3122V+c3222V+c3322V+c3422V+c3522V+c3622V+c3722V+c3822V+c3922V+c3A22V+c3B22V+c3C22V+c3D22V+c3E22V+c3F22V;
assign A322V=(C322V>=0)?1:0;

assign P422V=A322V;

//layer3 done, begain next layer
(*DONT_TOUCH="true"*) wire P5000;
(*DONT_TOUCH="true"*) wire P5001;
(*DONT_TOUCH="true"*) wire W40000,W40010,W40020,W40100,W40110,W40120,W40200,W40210,W40220;
(*DONT_TOUCH="true"*) wire W40001,W40011,W40021,W40101,W40111,W40121,W40201,W40211,W40221;
(*DONT_TOUCH="true"*) wire W40002,W40012,W40022,W40102,W40112,W40122,W40202,W40212,W40222;
(*DONT_TOUCH="true"*) wire W40003,W40013,W40023,W40103,W40113,W40123,W40203,W40213,W40223;
(*DONT_TOUCH="true"*) wire W40004,W40014,W40024,W40104,W40114,W40124,W40204,W40214,W40224;
(*DONT_TOUCH="true"*) wire W40005,W40015,W40025,W40105,W40115,W40125,W40205,W40215,W40225;
(*DONT_TOUCH="true"*) wire W40006,W40016,W40026,W40106,W40116,W40126,W40206,W40216,W40226;
(*DONT_TOUCH="true"*) wire W40007,W40017,W40027,W40107,W40117,W40127,W40207,W40217,W40227;
(*DONT_TOUCH="true"*) wire W40008,W40018,W40028,W40108,W40118,W40128,W40208,W40218,W40228;
(*DONT_TOUCH="true"*) wire W40009,W40019,W40029,W40109,W40119,W40129,W40209,W40219,W40229;
(*DONT_TOUCH="true"*) wire W4000A,W4001A,W4002A,W4010A,W4011A,W4012A,W4020A,W4021A,W4022A;
(*DONT_TOUCH="true"*) wire W4000B,W4001B,W4002B,W4010B,W4011B,W4012B,W4020B,W4021B,W4022B;
(*DONT_TOUCH="true"*) wire W4000C,W4001C,W4002C,W4010C,W4011C,W4012C,W4020C,W4021C,W4022C;
(*DONT_TOUCH="true"*) wire W4000D,W4001D,W4002D,W4010D,W4011D,W4012D,W4020D,W4021D,W4022D;
(*DONT_TOUCH="true"*) wire W4000E,W4001E,W4002E,W4010E,W4011E,W4012E,W4020E,W4021E,W4022E;
(*DONT_TOUCH="true"*) wire W4000F,W4001F,W4002F,W4010F,W4011F,W4012F,W4020F,W4021F,W4022F;
(*DONT_TOUCH="true"*) wire W4000G,W4001G,W4002G,W4010G,W4011G,W4012G,W4020G,W4021G,W4022G;
(*DONT_TOUCH="true"*) wire W4000H,W4001H,W4002H,W4010H,W4011H,W4012H,W4020H,W4021H,W4022H;
(*DONT_TOUCH="true"*) wire W4000I,W4001I,W4002I,W4010I,W4011I,W4012I,W4020I,W4021I,W4022I;
(*DONT_TOUCH="true"*) wire W4000J,W4001J,W4002J,W4010J,W4011J,W4012J,W4020J,W4021J,W4022J;
(*DONT_TOUCH="true"*) wire W4000K,W4001K,W4002K,W4010K,W4011K,W4012K,W4020K,W4021K,W4022K;
(*DONT_TOUCH="true"*) wire W4000L,W4001L,W4002L,W4010L,W4011L,W4012L,W4020L,W4021L,W4022L;
(*DONT_TOUCH="true"*) wire W4000M,W4001M,W4002M,W4010M,W4011M,W4012M,W4020M,W4021M,W4022M;
(*DONT_TOUCH="true"*) wire W4000N,W4001N,W4002N,W4010N,W4011N,W4012N,W4020N,W4021N,W4022N;
(*DONT_TOUCH="true"*) wire W4000O,W4001O,W4002O,W4010O,W4011O,W4012O,W4020O,W4021O,W4022O;
(*DONT_TOUCH="true"*) wire W4000P,W4001P,W4002P,W4010P,W4011P,W4012P,W4020P,W4021P,W4022P;
(*DONT_TOUCH="true"*) wire W4000Q,W4001Q,W4002Q,W4010Q,W4011Q,W4012Q,W4020Q,W4021Q,W4022Q;
(*DONT_TOUCH="true"*) wire W4000R,W4001R,W4002R,W4010R,W4011R,W4012R,W4020R,W4021R,W4022R;
(*DONT_TOUCH="true"*) wire W4000S,W4001S,W4002S,W4010S,W4011S,W4012S,W4020S,W4021S,W4022S;
(*DONT_TOUCH="true"*) wire W4000T,W4001T,W4002T,W4010T,W4011T,W4012T,W4020T,W4021T,W4022T;
(*DONT_TOUCH="true"*) wire W4000U,W4001U,W4002U,W4010U,W4011U,W4012U,W4020U,W4021U,W4022U;
(*DONT_TOUCH="true"*) wire W4000V,W4001V,W4002V,W4010V,W4011V,W4012V,W4020V,W4021V,W4022V;
(*DONT_TOUCH="true"*) wire W41000,W41010,W41020,W41100,W41110,W41120,W41200,W41210,W41220;
(*DONT_TOUCH="true"*) wire W41001,W41011,W41021,W41101,W41111,W41121,W41201,W41211,W41221;
(*DONT_TOUCH="true"*) wire W41002,W41012,W41022,W41102,W41112,W41122,W41202,W41212,W41222;
(*DONT_TOUCH="true"*) wire W41003,W41013,W41023,W41103,W41113,W41123,W41203,W41213,W41223;
(*DONT_TOUCH="true"*) wire W41004,W41014,W41024,W41104,W41114,W41124,W41204,W41214,W41224;
(*DONT_TOUCH="true"*) wire W41005,W41015,W41025,W41105,W41115,W41125,W41205,W41215,W41225;
(*DONT_TOUCH="true"*) wire W41006,W41016,W41026,W41106,W41116,W41126,W41206,W41216,W41226;
(*DONT_TOUCH="true"*) wire W41007,W41017,W41027,W41107,W41117,W41127,W41207,W41217,W41227;
(*DONT_TOUCH="true"*) wire W41008,W41018,W41028,W41108,W41118,W41128,W41208,W41218,W41228;
(*DONT_TOUCH="true"*) wire W41009,W41019,W41029,W41109,W41119,W41129,W41209,W41219,W41229;
(*DONT_TOUCH="true"*) wire W4100A,W4101A,W4102A,W4110A,W4111A,W4112A,W4120A,W4121A,W4122A;
(*DONT_TOUCH="true"*) wire W4100B,W4101B,W4102B,W4110B,W4111B,W4112B,W4120B,W4121B,W4122B;
(*DONT_TOUCH="true"*) wire W4100C,W4101C,W4102C,W4110C,W4111C,W4112C,W4120C,W4121C,W4122C;
(*DONT_TOUCH="true"*) wire W4100D,W4101D,W4102D,W4110D,W4111D,W4112D,W4120D,W4121D,W4122D;
(*DONT_TOUCH="true"*) wire W4100E,W4101E,W4102E,W4110E,W4111E,W4112E,W4120E,W4121E,W4122E;
(*DONT_TOUCH="true"*) wire W4100F,W4101F,W4102F,W4110F,W4111F,W4112F,W4120F,W4121F,W4122F;
(*DONT_TOUCH="true"*) wire W4100G,W4101G,W4102G,W4110G,W4111G,W4112G,W4120G,W4121G,W4122G;
(*DONT_TOUCH="true"*) wire W4100H,W4101H,W4102H,W4110H,W4111H,W4112H,W4120H,W4121H,W4122H;
(*DONT_TOUCH="true"*) wire W4100I,W4101I,W4102I,W4110I,W4111I,W4112I,W4120I,W4121I,W4122I;
(*DONT_TOUCH="true"*) wire W4100J,W4101J,W4102J,W4110J,W4111J,W4112J,W4120J,W4121J,W4122J;
(*DONT_TOUCH="true"*) wire W4100K,W4101K,W4102K,W4110K,W4111K,W4112K,W4120K,W4121K,W4122K;
(*DONT_TOUCH="true"*) wire W4100L,W4101L,W4102L,W4110L,W4111L,W4112L,W4120L,W4121L,W4122L;
(*DONT_TOUCH="true"*) wire W4100M,W4101M,W4102M,W4110M,W4111M,W4112M,W4120M,W4121M,W4122M;
(*DONT_TOUCH="true"*) wire W4100N,W4101N,W4102N,W4110N,W4111N,W4112N,W4120N,W4121N,W4122N;
(*DONT_TOUCH="true"*) wire W4100O,W4101O,W4102O,W4110O,W4111O,W4112O,W4120O,W4121O,W4122O;
(*DONT_TOUCH="true"*) wire W4100P,W4101P,W4102P,W4110P,W4111P,W4112P,W4120P,W4121P,W4122P;
(*DONT_TOUCH="true"*) wire W4100Q,W4101Q,W4102Q,W4110Q,W4111Q,W4112Q,W4120Q,W4121Q,W4122Q;
(*DONT_TOUCH="true"*) wire W4100R,W4101R,W4102R,W4110R,W4111R,W4112R,W4120R,W4121R,W4122R;
(*DONT_TOUCH="true"*) wire W4100S,W4101S,W4102S,W4110S,W4111S,W4112S,W4120S,W4121S,W4122S;
(*DONT_TOUCH="true"*) wire W4100T,W4101T,W4102T,W4110T,W4111T,W4112T,W4120T,W4121T,W4122T;
(*DONT_TOUCH="true"*) wire W4100U,W4101U,W4102U,W4110U,W4111U,W4112U,W4120U,W4121U,W4122U;
(*DONT_TOUCH="true"*) wire W4100V,W4101V,W4102V,W4110V,W4111V,W4112V,W4120V,W4121V,W4122V;
(*DONT_TOUCH="true"*) wire signed [4:0] c40000,c41000,c42000,c43000,c44000,c45000,c46000,c47000,c48000,c49000,c4A000,c4B000,c4C000,c4D000,c4E000,c4F000,c4G000,c4H000,c4I000,c4J000,c4K000,c4L000,c4M000,c4N000,c4O000,c4P000,c4Q000,c4R000,c4S000,c4T000,c4U000,c4V000;
(*DONT_TOUCH="true"*) wire signed [4:0] c40001,c41001,c42001,c43001,c44001,c45001,c46001,c47001,c48001,c49001,c4A001,c4B001,c4C001,c4D001,c4E001,c4F001,c4G001,c4H001,c4I001,c4J001,c4K001,c4L001,c4M001,c4N001,c4O001,c4P001,c4Q001,c4R001,c4S001,c4T001,c4U001,c4V001;
(*DONT_TOUCH="true"*) wire signed [9:0] C4000;
(*DONT_TOUCH="true"*) wire A4000;
(*DONT_TOUCH="true"*) wire signed [9:0] C4001;
(*DONT_TOUCH="true"*) wire A4001;
DFF_save_fm DFF_W5760(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40000));
DFF_save_fm DFF_W5761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40010));
DFF_save_fm DFF_W5762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40020));
DFF_save_fm DFF_W5763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40100));
DFF_save_fm DFF_W5764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40110));
DFF_save_fm DFF_W5765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40120));
DFF_save_fm DFF_W5766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40200));
DFF_save_fm DFF_W5767(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40210));
DFF_save_fm DFF_W5768(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40220));
DFF_save_fm DFF_W5769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40001));
DFF_save_fm DFF_W5770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40011));
DFF_save_fm DFF_W5771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40021));
DFF_save_fm DFF_W5772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40101));
DFF_save_fm DFF_W5773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40111));
DFF_save_fm DFF_W5774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40121));
DFF_save_fm DFF_W5775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40201));
DFF_save_fm DFF_W5776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40211));
DFF_save_fm DFF_W5777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40221));
DFF_save_fm DFF_W5778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40002));
DFF_save_fm DFF_W5779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40012));
DFF_save_fm DFF_W5780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40022));
DFF_save_fm DFF_W5781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40102));
DFF_save_fm DFF_W5782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40112));
DFF_save_fm DFF_W5783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40122));
DFF_save_fm DFF_W5784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40202));
DFF_save_fm DFF_W5785(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40212));
DFF_save_fm DFF_W5786(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40222));
DFF_save_fm DFF_W5787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40003));
DFF_save_fm DFF_W5788(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40013));
DFF_save_fm DFF_W5789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40023));
DFF_save_fm DFF_W5790(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40103));
DFF_save_fm DFF_W5791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40113));
DFF_save_fm DFF_W5792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40123));
DFF_save_fm DFF_W5793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40203));
DFF_save_fm DFF_W5794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40213));
DFF_save_fm DFF_W5795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40223));
DFF_save_fm DFF_W5796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40004));
DFF_save_fm DFF_W5797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40014));
DFF_save_fm DFF_W5798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40024));
DFF_save_fm DFF_W5799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40104));
DFF_save_fm DFF_W5800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40114));
DFF_save_fm DFF_W5801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40124));
DFF_save_fm DFF_W5802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40204));
DFF_save_fm DFF_W5803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40214));
DFF_save_fm DFF_W5804(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40224));
DFF_save_fm DFF_W5805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40005));
DFF_save_fm DFF_W5806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40015));
DFF_save_fm DFF_W5807(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40025));
DFF_save_fm DFF_W5808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40105));
DFF_save_fm DFF_W5809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40115));
DFF_save_fm DFF_W5810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40125));
DFF_save_fm DFF_W5811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40205));
DFF_save_fm DFF_W5812(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40215));
DFF_save_fm DFF_W5813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40225));
DFF_save_fm DFF_W5814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40006));
DFF_save_fm DFF_W5815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40016));
DFF_save_fm DFF_W5816(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40026));
DFF_save_fm DFF_W5817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40106));
DFF_save_fm DFF_W5818(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40116));
DFF_save_fm DFF_W5819(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40126));
DFF_save_fm DFF_W5820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40206));
DFF_save_fm DFF_W5821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40216));
DFF_save_fm DFF_W5822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40226));
DFF_save_fm DFF_W5823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40007));
DFF_save_fm DFF_W5824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40017));
DFF_save_fm DFF_W5825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40027));
DFF_save_fm DFF_W5826(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40107));
DFF_save_fm DFF_W5827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40117));
DFF_save_fm DFF_W5828(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40127));
DFF_save_fm DFF_W5829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40207));
DFF_save_fm DFF_W5830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40217));
DFF_save_fm DFF_W5831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40227));
DFF_save_fm DFF_W5832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40008));
DFF_save_fm DFF_W5833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40018));
DFF_save_fm DFF_W5834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40028));
DFF_save_fm DFF_W5835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40108));
DFF_save_fm DFF_W5836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40118));
DFF_save_fm DFF_W5837(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40128));
DFF_save_fm DFF_W5838(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40208));
DFF_save_fm DFF_W5839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40218));
DFF_save_fm DFF_W5840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40228));
DFF_save_fm DFF_W5841(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40009));
DFF_save_fm DFF_W5842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40019));
DFF_save_fm DFF_W5843(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40029));
DFF_save_fm DFF_W5844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40109));
DFF_save_fm DFF_W5845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40119));
DFF_save_fm DFF_W5846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40129));
DFF_save_fm DFF_W5847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40209));
DFF_save_fm DFF_W5848(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40219));
DFF_save_fm DFF_W5849(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40229));
DFF_save_fm DFF_W5850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000A));
DFF_save_fm DFF_W5851(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001A));
DFF_save_fm DFF_W5852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002A));
DFF_save_fm DFF_W5853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010A));
DFF_save_fm DFF_W5854(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011A));
DFF_save_fm DFF_W5855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012A));
DFF_save_fm DFF_W5856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020A));
DFF_save_fm DFF_W5857(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021A));
DFF_save_fm DFF_W5858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022A));
DFF_save_fm DFF_W5859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000B));
DFF_save_fm DFF_W5860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001B));
DFF_save_fm DFF_W5861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002B));
DFF_save_fm DFF_W5862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010B));
DFF_save_fm DFF_W5863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011B));
DFF_save_fm DFF_W5864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012B));
DFF_save_fm DFF_W5865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020B));
DFF_save_fm DFF_W5866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021B));
DFF_save_fm DFF_W5867(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022B));
DFF_save_fm DFF_W5868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000C));
DFF_save_fm DFF_W5869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001C));
DFF_save_fm DFF_W5870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002C));
DFF_save_fm DFF_W5871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010C));
DFF_save_fm DFF_W5872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011C));
DFF_save_fm DFF_W5873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012C));
DFF_save_fm DFF_W5874(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020C));
DFF_save_fm DFF_W5875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021C));
DFF_save_fm DFF_W5876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022C));
DFF_save_fm DFF_W5877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000D));
DFF_save_fm DFF_W5878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001D));
DFF_save_fm DFF_W5879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002D));
DFF_save_fm DFF_W5880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010D));
DFF_save_fm DFF_W5881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011D));
DFF_save_fm DFF_W5882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012D));
DFF_save_fm DFF_W5883(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020D));
DFF_save_fm DFF_W5884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021D));
DFF_save_fm DFF_W5885(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022D));
DFF_save_fm DFF_W5886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000E));
DFF_save_fm DFF_W5887(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001E));
DFF_save_fm DFF_W5888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002E));
DFF_save_fm DFF_W5889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010E));
DFF_save_fm DFF_W5890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011E));
DFF_save_fm DFF_W5891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012E));
DFF_save_fm DFF_W5892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020E));
DFF_save_fm DFF_W5893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021E));
DFF_save_fm DFF_W5894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022E));
DFF_save_fm DFF_W5895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000F));
DFF_save_fm DFF_W5896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001F));
DFF_save_fm DFF_W5897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002F));
DFF_save_fm DFF_W5898(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010F));
DFF_save_fm DFF_W5899(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011F));
DFF_save_fm DFF_W5900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012F));
DFF_save_fm DFF_W5901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020F));
DFF_save_fm DFF_W5902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021F));
DFF_save_fm DFF_W5903(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022F));
DFF_save_fm DFF_W5904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000G));
DFF_save_fm DFF_W5905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001G));
DFF_save_fm DFF_W5906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002G));
DFF_save_fm DFF_W5907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010G));
DFF_save_fm DFF_W5908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011G));
DFF_save_fm DFF_W5909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012G));
DFF_save_fm DFF_W5910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020G));
DFF_save_fm DFF_W5911(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021G));
DFF_save_fm DFF_W5912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022G));
DFF_save_fm DFF_W5913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000H));
DFF_save_fm DFF_W5914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001H));
DFF_save_fm DFF_W5915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002H));
DFF_save_fm DFF_W5916(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010H));
DFF_save_fm DFF_W5917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011H));
DFF_save_fm DFF_W5918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012H));
DFF_save_fm DFF_W5919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020H));
DFF_save_fm DFF_W5920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021H));
DFF_save_fm DFF_W5921(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022H));
DFF_save_fm DFF_W5922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000I));
DFF_save_fm DFF_W5923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001I));
DFF_save_fm DFF_W5924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002I));
DFF_save_fm DFF_W5925(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010I));
DFF_save_fm DFF_W5926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011I));
DFF_save_fm DFF_W5927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012I));
DFF_save_fm DFF_W5928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020I));
DFF_save_fm DFF_W5929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021I));
DFF_save_fm DFF_W5930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022I));
DFF_save_fm DFF_W5931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000J));
DFF_save_fm DFF_W5932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001J));
DFF_save_fm DFF_W5933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002J));
DFF_save_fm DFF_W5934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010J));
DFF_save_fm DFF_W5935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011J));
DFF_save_fm DFF_W5936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012J));
DFF_save_fm DFF_W5937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020J));
DFF_save_fm DFF_W5938(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021J));
DFF_save_fm DFF_W5939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022J));
DFF_save_fm DFF_W5940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000K));
DFF_save_fm DFF_W5941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001K));
DFF_save_fm DFF_W5942(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002K));
DFF_save_fm DFF_W5943(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010K));
DFF_save_fm DFF_W5944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011K));
DFF_save_fm DFF_W5945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012K));
DFF_save_fm DFF_W5946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020K));
DFF_save_fm DFF_W5947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021K));
DFF_save_fm DFF_W5948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022K));
DFF_save_fm DFF_W5949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000L));
DFF_save_fm DFF_W5950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001L));
DFF_save_fm DFF_W5951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002L));
DFF_save_fm DFF_W5952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010L));
DFF_save_fm DFF_W5953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011L));
DFF_save_fm DFF_W5954(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012L));
DFF_save_fm DFF_W5955(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020L));
DFF_save_fm DFF_W5956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021L));
DFF_save_fm DFF_W5957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022L));
DFF_save_fm DFF_W5958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000M));
DFF_save_fm DFF_W5959(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001M));
DFF_save_fm DFF_W5960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002M));
DFF_save_fm DFF_W5961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010M));
DFF_save_fm DFF_W5962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011M));
DFF_save_fm DFF_W5963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012M));
DFF_save_fm DFF_W5964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020M));
DFF_save_fm DFF_W5965(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021M));
DFF_save_fm DFF_W5966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022M));
DFF_save_fm DFF_W5967(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000N));
DFF_save_fm DFF_W5968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001N));
DFF_save_fm DFF_W5969(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002N));
DFF_save_fm DFF_W5970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010N));
DFF_save_fm DFF_W5971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011N));
DFF_save_fm DFF_W5972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012N));
DFF_save_fm DFF_W5973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020N));
DFF_save_fm DFF_W5974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021N));
DFF_save_fm DFF_W5975(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022N));
DFF_save_fm DFF_W5976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000O));
DFF_save_fm DFF_W5977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001O));
DFF_save_fm DFF_W5978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002O));
DFF_save_fm DFF_W5979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010O));
DFF_save_fm DFF_W5980(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011O));
DFF_save_fm DFF_W5981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012O));
DFF_save_fm DFF_W5982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020O));
DFF_save_fm DFF_W5983(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021O));
DFF_save_fm DFF_W5984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022O));
DFF_save_fm DFF_W5985(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000P));
DFF_save_fm DFF_W5986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001P));
DFF_save_fm DFF_W5987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002P));
DFF_save_fm DFF_W5988(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010P));
DFF_save_fm DFF_W5989(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011P));
DFF_save_fm DFF_W5990(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012P));
DFF_save_fm DFF_W5991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020P));
DFF_save_fm DFF_W5992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021P));
DFF_save_fm DFF_W5993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022P));
DFF_save_fm DFF_W5994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000Q));
DFF_save_fm DFF_W5995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001Q));
DFF_save_fm DFF_W5996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002Q));
DFF_save_fm DFF_W5997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010Q));
DFF_save_fm DFF_W5998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011Q));
DFF_save_fm DFF_W5999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012Q));
DFF_save_fm DFF_W6000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020Q));
DFF_save_fm DFF_W6001(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021Q));
DFF_save_fm DFF_W6002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022Q));
DFF_save_fm DFF_W6003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000R));
DFF_save_fm DFF_W6004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001R));
DFF_save_fm DFF_W6005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002R));
DFF_save_fm DFF_W6006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010R));
DFF_save_fm DFF_W6007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011R));
DFF_save_fm DFF_W6008(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012R));
DFF_save_fm DFF_W6009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020R));
DFF_save_fm DFF_W6010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021R));
DFF_save_fm DFF_W6011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022R));
DFF_save_fm DFF_W6012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000S));
DFF_save_fm DFF_W6013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001S));
DFF_save_fm DFF_W6014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002S));
DFF_save_fm DFF_W6015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010S));
DFF_save_fm DFF_W6016(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011S));
DFF_save_fm DFF_W6017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012S));
DFF_save_fm DFF_W6018(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020S));
DFF_save_fm DFF_W6019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021S));
DFF_save_fm DFF_W6020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022S));
DFF_save_fm DFF_W6021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000T));
DFF_save_fm DFF_W6022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001T));
DFF_save_fm DFF_W6023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002T));
DFF_save_fm DFF_W6024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010T));
DFF_save_fm DFF_W6025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011T));
DFF_save_fm DFF_W6026(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012T));
DFF_save_fm DFF_W6027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020T));
DFF_save_fm DFF_W6028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021T));
DFF_save_fm DFF_W6029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022T));
DFF_save_fm DFF_W6030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000U));
DFF_save_fm DFF_W6031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001U));
DFF_save_fm DFF_W6032(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002U));
DFF_save_fm DFF_W6033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010U));
DFF_save_fm DFF_W6034(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011U));
DFF_save_fm DFF_W6035(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012U));
DFF_save_fm DFF_W6036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020U));
DFF_save_fm DFF_W6037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021U));
DFF_save_fm DFF_W6038(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022U));
DFF_save_fm DFF_W6039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000V));
DFF_save_fm DFF_W6040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001V));
DFF_save_fm DFF_W6041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002V));
DFF_save_fm DFF_W6042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010V));
DFF_save_fm DFF_W6043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011V));
DFF_save_fm DFF_W6044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012V));
DFF_save_fm DFF_W6045(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020V));
DFF_save_fm DFF_W6046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021V));
DFF_save_fm DFF_W6047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022V));
DFF_save_fm DFF_W6048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41000));
DFF_save_fm DFF_W6049(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41010));
DFF_save_fm DFF_W6050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41020));
DFF_save_fm DFF_W6051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41100));
DFF_save_fm DFF_W6052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41110));
DFF_save_fm DFF_W6053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41120));
DFF_save_fm DFF_W6054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41200));
DFF_save_fm DFF_W6055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41210));
DFF_save_fm DFF_W6056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41220));
DFF_save_fm DFF_W6057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41001));
DFF_save_fm DFF_W6058(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41011));
DFF_save_fm DFF_W6059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41021));
DFF_save_fm DFF_W6060(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41101));
DFF_save_fm DFF_W6061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41111));
DFF_save_fm DFF_W6062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41121));
DFF_save_fm DFF_W6063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41201));
DFF_save_fm DFF_W6064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41211));
DFF_save_fm DFF_W6065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41221));
DFF_save_fm DFF_W6066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41002));
DFF_save_fm DFF_W6067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41012));
DFF_save_fm DFF_W6068(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41022));
DFF_save_fm DFF_W6069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41102));
DFF_save_fm DFF_W6070(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41112));
DFF_save_fm DFF_W6071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41122));
DFF_save_fm DFF_W6072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41202));
DFF_save_fm DFF_W6073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41212));
DFF_save_fm DFF_W6074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41222));
DFF_save_fm DFF_W6075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41003));
DFF_save_fm DFF_W6076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41013));
DFF_save_fm DFF_W6077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41023));
DFF_save_fm DFF_W6078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41103));
DFF_save_fm DFF_W6079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41113));
DFF_save_fm DFF_W6080(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41123));
DFF_save_fm DFF_W6081(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41203));
DFF_save_fm DFF_W6082(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41213));
DFF_save_fm DFF_W6083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41223));
DFF_save_fm DFF_W6084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41004));
DFF_save_fm DFF_W6085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41014));
DFF_save_fm DFF_W6086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41024));
DFF_save_fm DFF_W6087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41104));
DFF_save_fm DFF_W6088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41114));
DFF_save_fm DFF_W6089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41124));
DFF_save_fm DFF_W6090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41204));
DFF_save_fm DFF_W6091(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41214));
DFF_save_fm DFF_W6092(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41224));
DFF_save_fm DFF_W6093(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41005));
DFF_save_fm DFF_W6094(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41015));
DFF_save_fm DFF_W6095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41025));
DFF_save_fm DFF_W6096(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41105));
DFF_save_fm DFF_W6097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41115));
DFF_save_fm DFF_W6098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41125));
DFF_save_fm DFF_W6099(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41205));
DFF_save_fm DFF_W6100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41215));
DFF_save_fm DFF_W6101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41225));
DFF_save_fm DFF_W6102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41006));
DFF_save_fm DFF_W6103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41016));
DFF_save_fm DFF_W6104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41026));
DFF_save_fm DFF_W6105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41106));
DFF_save_fm DFF_W6106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41116));
DFF_save_fm DFF_W6107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41126));
DFF_save_fm DFF_W6108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41206));
DFF_save_fm DFF_W6109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41216));
DFF_save_fm DFF_W6110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41226));
DFF_save_fm DFF_W6111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41007));
DFF_save_fm DFF_W6112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41017));
DFF_save_fm DFF_W6113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41027));
DFF_save_fm DFF_W6114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41107));
DFF_save_fm DFF_W6115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41117));
DFF_save_fm DFF_W6116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41127));
DFF_save_fm DFF_W6117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41207));
DFF_save_fm DFF_W6118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41217));
DFF_save_fm DFF_W6119(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41227));
DFF_save_fm DFF_W6120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41008));
DFF_save_fm DFF_W6121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41018));
DFF_save_fm DFF_W6122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41028));
DFF_save_fm DFF_W6123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41108));
DFF_save_fm DFF_W6124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41118));
DFF_save_fm DFF_W6125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41128));
DFF_save_fm DFF_W6126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41208));
DFF_save_fm DFF_W6127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41218));
DFF_save_fm DFF_W6128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41228));
DFF_save_fm DFF_W6129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41009));
DFF_save_fm DFF_W6130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41019));
DFF_save_fm DFF_W6131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41029));
DFF_save_fm DFF_W6132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41109));
DFF_save_fm DFF_W6133(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41119));
DFF_save_fm DFF_W6134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41129));
DFF_save_fm DFF_W6135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41209));
DFF_save_fm DFF_W6136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41219));
DFF_save_fm DFF_W6137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41229));
DFF_save_fm DFF_W6138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100A));
DFF_save_fm DFF_W6139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101A));
DFF_save_fm DFF_W6140(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102A));
DFF_save_fm DFF_W6141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110A));
DFF_save_fm DFF_W6142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111A));
DFF_save_fm DFF_W6143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112A));
DFF_save_fm DFF_W6144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120A));
DFF_save_fm DFF_W6145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121A));
DFF_save_fm DFF_W6146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122A));
DFF_save_fm DFF_W6147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100B));
DFF_save_fm DFF_W6148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101B));
DFF_save_fm DFF_W6149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102B));
DFF_save_fm DFF_W6150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110B));
DFF_save_fm DFF_W6151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111B));
DFF_save_fm DFF_W6152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112B));
DFF_save_fm DFF_W6153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120B));
DFF_save_fm DFF_W6154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121B));
DFF_save_fm DFF_W6155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122B));
DFF_save_fm DFF_W6156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100C));
DFF_save_fm DFF_W6157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101C));
DFF_save_fm DFF_W6158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102C));
DFF_save_fm DFF_W6159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110C));
DFF_save_fm DFF_W6160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111C));
DFF_save_fm DFF_W6161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112C));
DFF_save_fm DFF_W6162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120C));
DFF_save_fm DFF_W6163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121C));
DFF_save_fm DFF_W6164(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122C));
DFF_save_fm DFF_W6165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100D));
DFF_save_fm DFF_W6166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101D));
DFF_save_fm DFF_W6167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102D));
DFF_save_fm DFF_W6168(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110D));
DFF_save_fm DFF_W6169(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111D));
DFF_save_fm DFF_W6170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112D));
DFF_save_fm DFF_W6171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120D));
DFF_save_fm DFF_W6172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121D));
DFF_save_fm DFF_W6173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122D));
DFF_save_fm DFF_W6174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100E));
DFF_save_fm DFF_W6175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101E));
DFF_save_fm DFF_W6176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102E));
DFF_save_fm DFF_W6177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110E));
DFF_save_fm DFF_W6178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111E));
DFF_save_fm DFF_W6179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112E));
DFF_save_fm DFF_W6180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120E));
DFF_save_fm DFF_W6181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121E));
DFF_save_fm DFF_W6182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122E));
DFF_save_fm DFF_W6183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100F));
DFF_save_fm DFF_W6184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101F));
DFF_save_fm DFF_W6185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102F));
DFF_save_fm DFF_W6186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110F));
DFF_save_fm DFF_W6187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111F));
DFF_save_fm DFF_W6188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112F));
DFF_save_fm DFF_W6189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120F));
DFF_save_fm DFF_W6190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121F));
DFF_save_fm DFF_W6191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122F));
DFF_save_fm DFF_W6192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100G));
DFF_save_fm DFF_W6193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101G));
DFF_save_fm DFF_W6194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102G));
DFF_save_fm DFF_W6195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110G));
DFF_save_fm DFF_W6196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111G));
DFF_save_fm DFF_W6197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112G));
DFF_save_fm DFF_W6198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120G));
DFF_save_fm DFF_W6199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121G));
DFF_save_fm DFF_W6200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122G));
DFF_save_fm DFF_W6201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100H));
DFF_save_fm DFF_W6202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101H));
DFF_save_fm DFF_W6203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102H));
DFF_save_fm DFF_W6204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110H));
DFF_save_fm DFF_W6205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111H));
DFF_save_fm DFF_W6206(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112H));
DFF_save_fm DFF_W6207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120H));
DFF_save_fm DFF_W6208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121H));
DFF_save_fm DFF_W6209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122H));
DFF_save_fm DFF_W6210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100I));
DFF_save_fm DFF_W6211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101I));
DFF_save_fm DFF_W6212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102I));
DFF_save_fm DFF_W6213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110I));
DFF_save_fm DFF_W6214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111I));
DFF_save_fm DFF_W6215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112I));
DFF_save_fm DFF_W6216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120I));
DFF_save_fm DFF_W6217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121I));
DFF_save_fm DFF_W6218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122I));
DFF_save_fm DFF_W6219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100J));
DFF_save_fm DFF_W6220(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101J));
DFF_save_fm DFF_W6221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102J));
DFF_save_fm DFF_W6222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110J));
DFF_save_fm DFF_W6223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111J));
DFF_save_fm DFF_W6224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112J));
DFF_save_fm DFF_W6225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120J));
DFF_save_fm DFF_W6226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121J));
DFF_save_fm DFF_W6227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122J));
DFF_save_fm DFF_W6228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100K));
DFF_save_fm DFF_W6229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101K));
DFF_save_fm DFF_W6230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102K));
DFF_save_fm DFF_W6231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110K));
DFF_save_fm DFF_W6232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111K));
DFF_save_fm DFF_W6233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112K));
DFF_save_fm DFF_W6234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120K));
DFF_save_fm DFF_W6235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121K));
DFF_save_fm DFF_W6236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122K));
DFF_save_fm DFF_W6237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100L));
DFF_save_fm DFF_W6238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101L));
DFF_save_fm DFF_W6239(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102L));
DFF_save_fm DFF_W6240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110L));
DFF_save_fm DFF_W6241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111L));
DFF_save_fm DFF_W6242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112L));
DFF_save_fm DFF_W6243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120L));
DFF_save_fm DFF_W6244(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121L));
DFF_save_fm DFF_W6245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122L));
DFF_save_fm DFF_W6246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100M));
DFF_save_fm DFF_W6247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101M));
DFF_save_fm DFF_W6248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102M));
DFF_save_fm DFF_W6249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110M));
DFF_save_fm DFF_W6250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111M));
DFF_save_fm DFF_W6251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112M));
DFF_save_fm DFF_W6252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120M));
DFF_save_fm DFF_W6253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121M));
DFF_save_fm DFF_W6254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122M));
DFF_save_fm DFF_W6255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100N));
DFF_save_fm DFF_W6256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101N));
DFF_save_fm DFF_W6257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102N));
DFF_save_fm DFF_W6258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110N));
DFF_save_fm DFF_W6259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111N));
DFF_save_fm DFF_W6260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112N));
DFF_save_fm DFF_W6261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120N));
DFF_save_fm DFF_W6262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121N));
DFF_save_fm DFF_W6263(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122N));
DFF_save_fm DFF_W6264(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100O));
DFF_save_fm DFF_W6265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101O));
DFF_save_fm DFF_W6266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102O));
DFF_save_fm DFF_W6267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110O));
DFF_save_fm DFF_W6268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111O));
DFF_save_fm DFF_W6269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112O));
DFF_save_fm DFF_W6270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120O));
DFF_save_fm DFF_W6271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121O));
DFF_save_fm DFF_W6272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122O));
DFF_save_fm DFF_W6273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100P));
DFF_save_fm DFF_W6274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101P));
DFF_save_fm DFF_W6275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102P));
DFF_save_fm DFF_W6276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110P));
DFF_save_fm DFF_W6277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111P));
DFF_save_fm DFF_W6278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112P));
DFF_save_fm DFF_W6279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120P));
DFF_save_fm DFF_W6280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121P));
DFF_save_fm DFF_W6281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122P));
DFF_save_fm DFF_W6282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100Q));
DFF_save_fm DFF_W6283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101Q));
DFF_save_fm DFF_W6284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102Q));
DFF_save_fm DFF_W6285(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110Q));
DFF_save_fm DFF_W6286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111Q));
DFF_save_fm DFF_W6287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112Q));
DFF_save_fm DFF_W6288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120Q));
DFF_save_fm DFF_W6289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121Q));
DFF_save_fm DFF_W6290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122Q));
DFF_save_fm DFF_W6291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100R));
DFF_save_fm DFF_W6292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101R));
DFF_save_fm DFF_W6293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102R));
DFF_save_fm DFF_W6294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110R));
DFF_save_fm DFF_W6295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111R));
DFF_save_fm DFF_W6296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112R));
DFF_save_fm DFF_W6297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120R));
DFF_save_fm DFF_W6298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121R));
DFF_save_fm DFF_W6299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122R));
DFF_save_fm DFF_W6300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100S));
DFF_save_fm DFF_W6301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101S));
DFF_save_fm DFF_W6302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102S));
DFF_save_fm DFF_W6303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110S));
DFF_save_fm DFF_W6304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111S));
DFF_save_fm DFF_W6305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112S));
DFF_save_fm DFF_W6306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120S));
DFF_save_fm DFF_W6307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121S));
DFF_save_fm DFF_W6308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122S));
DFF_save_fm DFF_W6309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100T));
DFF_save_fm DFF_W6310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101T));
DFF_save_fm DFF_W6311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102T));
DFF_save_fm DFF_W6312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110T));
DFF_save_fm DFF_W6313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111T));
DFF_save_fm DFF_W6314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112T));
DFF_save_fm DFF_W6315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120T));
DFF_save_fm DFF_W6316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121T));
DFF_save_fm DFF_W6317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122T));
DFF_save_fm DFF_W6318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100U));
DFF_save_fm DFF_W6319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101U));
DFF_save_fm DFF_W6320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102U));
DFF_save_fm DFF_W6321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110U));
DFF_save_fm DFF_W6322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111U));
DFF_save_fm DFF_W6323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112U));
DFF_save_fm DFF_W6324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120U));
DFF_save_fm DFF_W6325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121U));
DFF_save_fm DFF_W6326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122U));
DFF_save_fm DFF_W6327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100V));
DFF_save_fm DFF_W6328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101V));
DFF_save_fm DFF_W6329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102V));
DFF_save_fm DFF_W6330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110V));
DFF_save_fm DFF_W6331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111V));
DFF_save_fm DFF_W6332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112V));
DFF_save_fm DFF_W6333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120V));
DFF_save_fm DFF_W6334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121V));
DFF_save_fm DFF_W6335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122V));
ninexnine_unit ninexnine_unit_7808(
				.clk(clk),
				.rstn(rstn),
				.a0(P4000),
				.a1(P4010),
				.a2(P4020),
				.a3(P4100),
				.a4(P4110),
				.a5(P4120),
				.a6(P4200),
				.a7(P4210),
				.a8(P4220),
				.b0(W40000),
				.b1(W40010),
				.b2(W40020),
				.b3(W40100),
				.b4(W40110),
				.b5(W40120),
				.b6(W40200),
				.b7(W40210),
				.b8(W40220),
				.c(c40000)
);

ninexnine_unit ninexnine_unit_7809(
				.clk(clk),
				.rstn(rstn),
				.a0(P4001),
				.a1(P4011),
				.a2(P4021),
				.a3(P4101),
				.a4(P4111),
				.a5(P4121),
				.a6(P4201),
				.a7(P4211),
				.a8(P4221),
				.b0(W40001),
				.b1(W40011),
				.b2(W40021),
				.b3(W40101),
				.b4(W40111),
				.b5(W40121),
				.b6(W40201),
				.b7(W40211),
				.b8(W40221),
				.c(c41000)
);

ninexnine_unit ninexnine_unit_7810(
				.clk(clk),
				.rstn(rstn),
				.a0(P4002),
				.a1(P4012),
				.a2(P4022),
				.a3(P4102),
				.a4(P4112),
				.a5(P4122),
				.a6(P4202),
				.a7(P4212),
				.a8(P4222),
				.b0(W40002),
				.b1(W40012),
				.b2(W40022),
				.b3(W40102),
				.b4(W40112),
				.b5(W40122),
				.b6(W40202),
				.b7(W40212),
				.b8(W40222),
				.c(c42000)
);

ninexnine_unit ninexnine_unit_7811(
				.clk(clk),
				.rstn(rstn),
				.a0(P4003),
				.a1(P4013),
				.a2(P4023),
				.a3(P4103),
				.a4(P4113),
				.a5(P4123),
				.a6(P4203),
				.a7(P4213),
				.a8(P4223),
				.b0(W40003),
				.b1(W40013),
				.b2(W40023),
				.b3(W40103),
				.b4(W40113),
				.b5(W40123),
				.b6(W40203),
				.b7(W40213),
				.b8(W40223),
				.c(c43000)
);

ninexnine_unit ninexnine_unit_7812(
				.clk(clk),
				.rstn(rstn),
				.a0(P4004),
				.a1(P4014),
				.a2(P4024),
				.a3(P4104),
				.a4(P4114),
				.a5(P4124),
				.a6(P4204),
				.a7(P4214),
				.a8(P4224),
				.b0(W40004),
				.b1(W40014),
				.b2(W40024),
				.b3(W40104),
				.b4(W40114),
				.b5(W40124),
				.b6(W40204),
				.b7(W40214),
				.b8(W40224),
				.c(c44000)
);

ninexnine_unit ninexnine_unit_7813(
				.clk(clk),
				.rstn(rstn),
				.a0(P4005),
				.a1(P4015),
				.a2(P4025),
				.a3(P4105),
				.a4(P4115),
				.a5(P4125),
				.a6(P4205),
				.a7(P4215),
				.a8(P4225),
				.b0(W40005),
				.b1(W40015),
				.b2(W40025),
				.b3(W40105),
				.b4(W40115),
				.b5(W40125),
				.b6(W40205),
				.b7(W40215),
				.b8(W40225),
				.c(c45000)
);

ninexnine_unit ninexnine_unit_7814(
				.clk(clk),
				.rstn(rstn),
				.a0(P4006),
				.a1(P4016),
				.a2(P4026),
				.a3(P4106),
				.a4(P4116),
				.a5(P4126),
				.a6(P4206),
				.a7(P4216),
				.a8(P4226),
				.b0(W40006),
				.b1(W40016),
				.b2(W40026),
				.b3(W40106),
				.b4(W40116),
				.b5(W40126),
				.b6(W40206),
				.b7(W40216),
				.b8(W40226),
				.c(c46000)
);

ninexnine_unit ninexnine_unit_7815(
				.clk(clk),
				.rstn(rstn),
				.a0(P4007),
				.a1(P4017),
				.a2(P4027),
				.a3(P4107),
				.a4(P4117),
				.a5(P4127),
				.a6(P4207),
				.a7(P4217),
				.a8(P4227),
				.b0(W40007),
				.b1(W40017),
				.b2(W40027),
				.b3(W40107),
				.b4(W40117),
				.b5(W40127),
				.b6(W40207),
				.b7(W40217),
				.b8(W40227),
				.c(c47000)
);

ninexnine_unit ninexnine_unit_7816(
				.clk(clk),
				.rstn(rstn),
				.a0(P4008),
				.a1(P4018),
				.a2(P4028),
				.a3(P4108),
				.a4(P4118),
				.a5(P4128),
				.a6(P4208),
				.a7(P4218),
				.a8(P4228),
				.b0(W40008),
				.b1(W40018),
				.b2(W40028),
				.b3(W40108),
				.b4(W40118),
				.b5(W40128),
				.b6(W40208),
				.b7(W40218),
				.b8(W40228),
				.c(c48000)
);

ninexnine_unit ninexnine_unit_7817(
				.clk(clk),
				.rstn(rstn),
				.a0(P4009),
				.a1(P4019),
				.a2(P4029),
				.a3(P4109),
				.a4(P4119),
				.a5(P4129),
				.a6(P4209),
				.a7(P4219),
				.a8(P4229),
				.b0(W40009),
				.b1(W40019),
				.b2(W40029),
				.b3(W40109),
				.b4(W40119),
				.b5(W40129),
				.b6(W40209),
				.b7(W40219),
				.b8(W40229),
				.c(c49000)
);

ninexnine_unit ninexnine_unit_7818(
				.clk(clk),
				.rstn(rstn),
				.a0(P400A),
				.a1(P401A),
				.a2(P402A),
				.a3(P410A),
				.a4(P411A),
				.a5(P412A),
				.a6(P420A),
				.a7(P421A),
				.a8(P422A),
				.b0(W4000A),
				.b1(W4001A),
				.b2(W4002A),
				.b3(W4010A),
				.b4(W4011A),
				.b5(W4012A),
				.b6(W4020A),
				.b7(W4021A),
				.b8(W4022A),
				.c(c4A000)
);

ninexnine_unit ninexnine_unit_7819(
				.clk(clk),
				.rstn(rstn),
				.a0(P400B),
				.a1(P401B),
				.a2(P402B),
				.a3(P410B),
				.a4(P411B),
				.a5(P412B),
				.a6(P420B),
				.a7(P421B),
				.a8(P422B),
				.b0(W4000B),
				.b1(W4001B),
				.b2(W4002B),
				.b3(W4010B),
				.b4(W4011B),
				.b5(W4012B),
				.b6(W4020B),
				.b7(W4021B),
				.b8(W4022B),
				.c(c4B000)
);

ninexnine_unit ninexnine_unit_7820(
				.clk(clk),
				.rstn(rstn),
				.a0(P400C),
				.a1(P401C),
				.a2(P402C),
				.a3(P410C),
				.a4(P411C),
				.a5(P412C),
				.a6(P420C),
				.a7(P421C),
				.a8(P422C),
				.b0(W4000C),
				.b1(W4001C),
				.b2(W4002C),
				.b3(W4010C),
				.b4(W4011C),
				.b5(W4012C),
				.b6(W4020C),
				.b7(W4021C),
				.b8(W4022C),
				.c(c4C000)
);

ninexnine_unit ninexnine_unit_7821(
				.clk(clk),
				.rstn(rstn),
				.a0(P400D),
				.a1(P401D),
				.a2(P402D),
				.a3(P410D),
				.a4(P411D),
				.a5(P412D),
				.a6(P420D),
				.a7(P421D),
				.a8(P422D),
				.b0(W4000D),
				.b1(W4001D),
				.b2(W4002D),
				.b3(W4010D),
				.b4(W4011D),
				.b5(W4012D),
				.b6(W4020D),
				.b7(W4021D),
				.b8(W4022D),
				.c(c4D000)
);

ninexnine_unit ninexnine_unit_7822(
				.clk(clk),
				.rstn(rstn),
				.a0(P400E),
				.a1(P401E),
				.a2(P402E),
				.a3(P410E),
				.a4(P411E),
				.a5(P412E),
				.a6(P420E),
				.a7(P421E),
				.a8(P422E),
				.b0(W4000E),
				.b1(W4001E),
				.b2(W4002E),
				.b3(W4010E),
				.b4(W4011E),
				.b5(W4012E),
				.b6(W4020E),
				.b7(W4021E),
				.b8(W4022E),
				.c(c4E000)
);

ninexnine_unit ninexnine_unit_7823(
				.clk(clk),
				.rstn(rstn),
				.a0(P400F),
				.a1(P401F),
				.a2(P402F),
				.a3(P410F),
				.a4(P411F),
				.a5(P412F),
				.a6(P420F),
				.a7(P421F),
				.a8(P422F),
				.b0(W4000F),
				.b1(W4001F),
				.b2(W4002F),
				.b3(W4010F),
				.b4(W4011F),
				.b5(W4012F),
				.b6(W4020F),
				.b7(W4021F),
				.b8(W4022F),
				.c(c4F000)
);

ninexnine_unit ninexnine_unit_7824(
				.clk(clk),
				.rstn(rstn),
				.a0(P400G),
				.a1(P401G),
				.a2(P402G),
				.a3(P410G),
				.a4(P411G),
				.a5(P412G),
				.a6(P420G),
				.a7(P421G),
				.a8(P422G),
				.b0(W4000G),
				.b1(W4001G),
				.b2(W4002G),
				.b3(W4010G),
				.b4(W4011G),
				.b5(W4012G),
				.b6(W4020G),
				.b7(W4021G),
				.b8(W4022G),
				.c(c4G000)
);

ninexnine_unit ninexnine_unit_7825(
				.clk(clk),
				.rstn(rstn),
				.a0(P400H),
				.a1(P401H),
				.a2(P402H),
				.a3(P410H),
				.a4(P411H),
				.a5(P412H),
				.a6(P420H),
				.a7(P421H),
				.a8(P422H),
				.b0(W4000H),
				.b1(W4001H),
				.b2(W4002H),
				.b3(W4010H),
				.b4(W4011H),
				.b5(W4012H),
				.b6(W4020H),
				.b7(W4021H),
				.b8(W4022H),
				.c(c4H000)
);

ninexnine_unit ninexnine_unit_7826(
				.clk(clk),
				.rstn(rstn),
				.a0(P400I),
				.a1(P401I),
				.a2(P402I),
				.a3(P410I),
				.a4(P411I),
				.a5(P412I),
				.a6(P420I),
				.a7(P421I),
				.a8(P422I),
				.b0(W4000I),
				.b1(W4001I),
				.b2(W4002I),
				.b3(W4010I),
				.b4(W4011I),
				.b5(W4012I),
				.b6(W4020I),
				.b7(W4021I),
				.b8(W4022I),
				.c(c4I000)
);

ninexnine_unit ninexnine_unit_7827(
				.clk(clk),
				.rstn(rstn),
				.a0(P400J),
				.a1(P401J),
				.a2(P402J),
				.a3(P410J),
				.a4(P411J),
				.a5(P412J),
				.a6(P420J),
				.a7(P421J),
				.a8(P422J),
				.b0(W4000J),
				.b1(W4001J),
				.b2(W4002J),
				.b3(W4010J),
				.b4(W4011J),
				.b5(W4012J),
				.b6(W4020J),
				.b7(W4021J),
				.b8(W4022J),
				.c(c4J000)
);

ninexnine_unit ninexnine_unit_7828(
				.clk(clk),
				.rstn(rstn),
				.a0(P400K),
				.a1(P401K),
				.a2(P402K),
				.a3(P410K),
				.a4(P411K),
				.a5(P412K),
				.a6(P420K),
				.a7(P421K),
				.a8(P422K),
				.b0(W4000K),
				.b1(W4001K),
				.b2(W4002K),
				.b3(W4010K),
				.b4(W4011K),
				.b5(W4012K),
				.b6(W4020K),
				.b7(W4021K),
				.b8(W4022K),
				.c(c4K000)
);

ninexnine_unit ninexnine_unit_7829(
				.clk(clk),
				.rstn(rstn),
				.a0(P400L),
				.a1(P401L),
				.a2(P402L),
				.a3(P410L),
				.a4(P411L),
				.a5(P412L),
				.a6(P420L),
				.a7(P421L),
				.a8(P422L),
				.b0(W4000L),
				.b1(W4001L),
				.b2(W4002L),
				.b3(W4010L),
				.b4(W4011L),
				.b5(W4012L),
				.b6(W4020L),
				.b7(W4021L),
				.b8(W4022L),
				.c(c4L000)
);

ninexnine_unit ninexnine_unit_7830(
				.clk(clk),
				.rstn(rstn),
				.a0(P400M),
				.a1(P401M),
				.a2(P402M),
				.a3(P410M),
				.a4(P411M),
				.a5(P412M),
				.a6(P420M),
				.a7(P421M),
				.a8(P422M),
				.b0(W4000M),
				.b1(W4001M),
				.b2(W4002M),
				.b3(W4010M),
				.b4(W4011M),
				.b5(W4012M),
				.b6(W4020M),
				.b7(W4021M),
				.b8(W4022M),
				.c(c4M000)
);

ninexnine_unit ninexnine_unit_7831(
				.clk(clk),
				.rstn(rstn),
				.a0(P400N),
				.a1(P401N),
				.a2(P402N),
				.a3(P410N),
				.a4(P411N),
				.a5(P412N),
				.a6(P420N),
				.a7(P421N),
				.a8(P422N),
				.b0(W4000N),
				.b1(W4001N),
				.b2(W4002N),
				.b3(W4010N),
				.b4(W4011N),
				.b5(W4012N),
				.b6(W4020N),
				.b7(W4021N),
				.b8(W4022N),
				.c(c4N000)
);

ninexnine_unit ninexnine_unit_7832(
				.clk(clk),
				.rstn(rstn),
				.a0(P400O),
				.a1(P401O),
				.a2(P402O),
				.a3(P410O),
				.a4(P411O),
				.a5(P412O),
				.a6(P420O),
				.a7(P421O),
				.a8(P422O),
				.b0(W4000O),
				.b1(W4001O),
				.b2(W4002O),
				.b3(W4010O),
				.b4(W4011O),
				.b5(W4012O),
				.b6(W4020O),
				.b7(W4021O),
				.b8(W4022O),
				.c(c4O000)
);

ninexnine_unit ninexnine_unit_7833(
				.clk(clk),
				.rstn(rstn),
				.a0(P400P),
				.a1(P401P),
				.a2(P402P),
				.a3(P410P),
				.a4(P411P),
				.a5(P412P),
				.a6(P420P),
				.a7(P421P),
				.a8(P422P),
				.b0(W4000P),
				.b1(W4001P),
				.b2(W4002P),
				.b3(W4010P),
				.b4(W4011P),
				.b5(W4012P),
				.b6(W4020P),
				.b7(W4021P),
				.b8(W4022P),
				.c(c4P000)
);

ninexnine_unit ninexnine_unit_7834(
				.clk(clk),
				.rstn(rstn),
				.a0(P400Q),
				.a1(P401Q),
				.a2(P402Q),
				.a3(P410Q),
				.a4(P411Q),
				.a5(P412Q),
				.a6(P420Q),
				.a7(P421Q),
				.a8(P422Q),
				.b0(W4000Q),
				.b1(W4001Q),
				.b2(W4002Q),
				.b3(W4010Q),
				.b4(W4011Q),
				.b5(W4012Q),
				.b6(W4020Q),
				.b7(W4021Q),
				.b8(W4022Q),
				.c(c4Q000)
);

ninexnine_unit ninexnine_unit_7835(
				.clk(clk),
				.rstn(rstn),
				.a0(P400R),
				.a1(P401R),
				.a2(P402R),
				.a3(P410R),
				.a4(P411R),
				.a5(P412R),
				.a6(P420R),
				.a7(P421R),
				.a8(P422R),
				.b0(W4000R),
				.b1(W4001R),
				.b2(W4002R),
				.b3(W4010R),
				.b4(W4011R),
				.b5(W4012R),
				.b6(W4020R),
				.b7(W4021R),
				.b8(W4022R),
				.c(c4R000)
);

ninexnine_unit ninexnine_unit_7836(
				.clk(clk),
				.rstn(rstn),
				.a0(P400S),
				.a1(P401S),
				.a2(P402S),
				.a3(P410S),
				.a4(P411S),
				.a5(P412S),
				.a6(P420S),
				.a7(P421S),
				.a8(P422S),
				.b0(W4000S),
				.b1(W4001S),
				.b2(W4002S),
				.b3(W4010S),
				.b4(W4011S),
				.b5(W4012S),
				.b6(W4020S),
				.b7(W4021S),
				.b8(W4022S),
				.c(c4S000)
);

ninexnine_unit ninexnine_unit_7837(
				.clk(clk),
				.rstn(rstn),
				.a0(P400T),
				.a1(P401T),
				.a2(P402T),
				.a3(P410T),
				.a4(P411T),
				.a5(P412T),
				.a6(P420T),
				.a7(P421T),
				.a8(P422T),
				.b0(W4000T),
				.b1(W4001T),
				.b2(W4002T),
				.b3(W4010T),
				.b4(W4011T),
				.b5(W4012T),
				.b6(W4020T),
				.b7(W4021T),
				.b8(W4022T),
				.c(c4T000)
);

ninexnine_unit ninexnine_unit_7838(
				.clk(clk),
				.rstn(rstn),
				.a0(P400U),
				.a1(P401U),
				.a2(P402U),
				.a3(P410U),
				.a4(P411U),
				.a5(P412U),
				.a6(P420U),
				.a7(P421U),
				.a8(P422U),
				.b0(W4000U),
				.b1(W4001U),
				.b2(W4002U),
				.b3(W4010U),
				.b4(W4011U),
				.b5(W4012U),
				.b6(W4020U),
				.b7(W4021U),
				.b8(W4022U),
				.c(c4U000)
);

ninexnine_unit ninexnine_unit_7839(
				.clk(clk),
				.rstn(rstn),
				.a0(P400V),
				.a1(P401V),
				.a2(P402V),
				.a3(P410V),
				.a4(P411V),
				.a5(P412V),
				.a6(P420V),
				.a7(P421V),
				.a8(P422V),
				.b0(W4000V),
				.b1(W4001V),
				.b2(W4002V),
				.b3(W4010V),
				.b4(W4011V),
				.b5(W4012V),
				.b6(W4020V),
				.b7(W4021V),
				.b8(W4022V),
				.c(c4V000)
);

assign C4000=c40000+c41000+c42000+c43000+c44000+c45000+c46000+c47000+c48000+c49000+c4A000+c4B000+c4C000+c4D000+c4E000+c4F000+c4G000+c4H000+c4I000+c4J000+c4K000+c4L000+c4M000+c4N000+c4O000+c4P000+c4Q000+c4R000+c4S000+c4T000+c4U000+c4V000;
assign A4000=(C4000>=0)?1:0;

assign P5000=A4000;

ninexnine_unit ninexnine_unit_7840(
				.clk(clk),
				.rstn(rstn),
				.a0(P4000),
				.a1(P4010),
				.a2(P4020),
				.a3(P4100),
				.a4(P4110),
				.a5(P4120),
				.a6(P4200),
				.a7(P4210),
				.a8(P4220),
				.b0(W41000),
				.b1(W41010),
				.b2(W41020),
				.b3(W41100),
				.b4(W41110),
				.b5(W41120),
				.b6(W41200),
				.b7(W41210),
				.b8(W41220),
				.c(c40001)
);

ninexnine_unit ninexnine_unit_7841(
				.clk(clk),
				.rstn(rstn),
				.a0(P4001),
				.a1(P4011),
				.a2(P4021),
				.a3(P4101),
				.a4(P4111),
				.a5(P4121),
				.a6(P4201),
				.a7(P4211),
				.a8(P4221),
				.b0(W41001),
				.b1(W41011),
				.b2(W41021),
				.b3(W41101),
				.b4(W41111),
				.b5(W41121),
				.b6(W41201),
				.b7(W41211),
				.b8(W41221),
				.c(c41001)
);

ninexnine_unit ninexnine_unit_7842(
				.clk(clk),
				.rstn(rstn),
				.a0(P4002),
				.a1(P4012),
				.a2(P4022),
				.a3(P4102),
				.a4(P4112),
				.a5(P4122),
				.a6(P4202),
				.a7(P4212),
				.a8(P4222),
				.b0(W41002),
				.b1(W41012),
				.b2(W41022),
				.b3(W41102),
				.b4(W41112),
				.b5(W41122),
				.b6(W41202),
				.b7(W41212),
				.b8(W41222),
				.c(c42001)
);

ninexnine_unit ninexnine_unit_7843(
				.clk(clk),
				.rstn(rstn),
				.a0(P4003),
				.a1(P4013),
				.a2(P4023),
				.a3(P4103),
				.a4(P4113),
				.a5(P4123),
				.a6(P4203),
				.a7(P4213),
				.a8(P4223),
				.b0(W41003),
				.b1(W41013),
				.b2(W41023),
				.b3(W41103),
				.b4(W41113),
				.b5(W41123),
				.b6(W41203),
				.b7(W41213),
				.b8(W41223),
				.c(c43001)
);

ninexnine_unit ninexnine_unit_7844(
				.clk(clk),
				.rstn(rstn),
				.a0(P4004),
				.a1(P4014),
				.a2(P4024),
				.a3(P4104),
				.a4(P4114),
				.a5(P4124),
				.a6(P4204),
				.a7(P4214),
				.a8(P4224),
				.b0(W41004),
				.b1(W41014),
				.b2(W41024),
				.b3(W41104),
				.b4(W41114),
				.b5(W41124),
				.b6(W41204),
				.b7(W41214),
				.b8(W41224),
				.c(c44001)
);

ninexnine_unit ninexnine_unit_7845(
				.clk(clk),
				.rstn(rstn),
				.a0(P4005),
				.a1(P4015),
				.a2(P4025),
				.a3(P4105),
				.a4(P4115),
				.a5(P4125),
				.a6(P4205),
				.a7(P4215),
				.a8(P4225),
				.b0(W41005),
				.b1(W41015),
				.b2(W41025),
				.b3(W41105),
				.b4(W41115),
				.b5(W41125),
				.b6(W41205),
				.b7(W41215),
				.b8(W41225),
				.c(c45001)
);

ninexnine_unit ninexnine_unit_7846(
				.clk(clk),
				.rstn(rstn),
				.a0(P4006),
				.a1(P4016),
				.a2(P4026),
				.a3(P4106),
				.a4(P4116),
				.a5(P4126),
				.a6(P4206),
				.a7(P4216),
				.a8(P4226),
				.b0(W41006),
				.b1(W41016),
				.b2(W41026),
				.b3(W41106),
				.b4(W41116),
				.b5(W41126),
				.b6(W41206),
				.b7(W41216),
				.b8(W41226),
				.c(c46001)
);

ninexnine_unit ninexnine_unit_7847(
				.clk(clk),
				.rstn(rstn),
				.a0(P4007),
				.a1(P4017),
				.a2(P4027),
				.a3(P4107),
				.a4(P4117),
				.a5(P4127),
				.a6(P4207),
				.a7(P4217),
				.a8(P4227),
				.b0(W41007),
				.b1(W41017),
				.b2(W41027),
				.b3(W41107),
				.b4(W41117),
				.b5(W41127),
				.b6(W41207),
				.b7(W41217),
				.b8(W41227),
				.c(c47001)
);

ninexnine_unit ninexnine_unit_7848(
				.clk(clk),
				.rstn(rstn),
				.a0(P4008),
				.a1(P4018),
				.a2(P4028),
				.a3(P4108),
				.a4(P4118),
				.a5(P4128),
				.a6(P4208),
				.a7(P4218),
				.a8(P4228),
				.b0(W41008),
				.b1(W41018),
				.b2(W41028),
				.b3(W41108),
				.b4(W41118),
				.b5(W41128),
				.b6(W41208),
				.b7(W41218),
				.b8(W41228),
				.c(c48001)
);

ninexnine_unit ninexnine_unit_7849(
				.clk(clk),
				.rstn(rstn),
				.a0(P4009),
				.a1(P4019),
				.a2(P4029),
				.a3(P4109),
				.a4(P4119),
				.a5(P4129),
				.a6(P4209),
				.a7(P4219),
				.a8(P4229),
				.b0(W41009),
				.b1(W41019),
				.b2(W41029),
				.b3(W41109),
				.b4(W41119),
				.b5(W41129),
				.b6(W41209),
				.b7(W41219),
				.b8(W41229),
				.c(c49001)
);

ninexnine_unit ninexnine_unit_7850(
				.clk(clk),
				.rstn(rstn),
				.a0(P400A),
				.a1(P401A),
				.a2(P402A),
				.a3(P410A),
				.a4(P411A),
				.a5(P412A),
				.a6(P420A),
				.a7(P421A),
				.a8(P422A),
				.b0(W4100A),
				.b1(W4101A),
				.b2(W4102A),
				.b3(W4110A),
				.b4(W4111A),
				.b5(W4112A),
				.b6(W4120A),
				.b7(W4121A),
				.b8(W4122A),
				.c(c4A001)
);

ninexnine_unit ninexnine_unit_7851(
				.clk(clk),
				.rstn(rstn),
				.a0(P400B),
				.a1(P401B),
				.a2(P402B),
				.a3(P410B),
				.a4(P411B),
				.a5(P412B),
				.a6(P420B),
				.a7(P421B),
				.a8(P422B),
				.b0(W4100B),
				.b1(W4101B),
				.b2(W4102B),
				.b3(W4110B),
				.b4(W4111B),
				.b5(W4112B),
				.b6(W4120B),
				.b7(W4121B),
				.b8(W4122B),
				.c(c4B001)
);

ninexnine_unit ninexnine_unit_7852(
				.clk(clk),
				.rstn(rstn),
				.a0(P400C),
				.a1(P401C),
				.a2(P402C),
				.a3(P410C),
				.a4(P411C),
				.a5(P412C),
				.a6(P420C),
				.a7(P421C),
				.a8(P422C),
				.b0(W4100C),
				.b1(W4101C),
				.b2(W4102C),
				.b3(W4110C),
				.b4(W4111C),
				.b5(W4112C),
				.b6(W4120C),
				.b7(W4121C),
				.b8(W4122C),
				.c(c4C001)
);

ninexnine_unit ninexnine_unit_7853(
				.clk(clk),
				.rstn(rstn),
				.a0(P400D),
				.a1(P401D),
				.a2(P402D),
				.a3(P410D),
				.a4(P411D),
				.a5(P412D),
				.a6(P420D),
				.a7(P421D),
				.a8(P422D),
				.b0(W4100D),
				.b1(W4101D),
				.b2(W4102D),
				.b3(W4110D),
				.b4(W4111D),
				.b5(W4112D),
				.b6(W4120D),
				.b7(W4121D),
				.b8(W4122D),
				.c(c4D001)
);

ninexnine_unit ninexnine_unit_7854(
				.clk(clk),
				.rstn(rstn),
				.a0(P400E),
				.a1(P401E),
				.a2(P402E),
				.a3(P410E),
				.a4(P411E),
				.a5(P412E),
				.a6(P420E),
				.a7(P421E),
				.a8(P422E),
				.b0(W4100E),
				.b1(W4101E),
				.b2(W4102E),
				.b3(W4110E),
				.b4(W4111E),
				.b5(W4112E),
				.b6(W4120E),
				.b7(W4121E),
				.b8(W4122E),
				.c(c4E001)
);

ninexnine_unit ninexnine_unit_7855(
				.clk(clk),
				.rstn(rstn),
				.a0(P400F),
				.a1(P401F),
				.a2(P402F),
				.a3(P410F),
				.a4(P411F),
				.a5(P412F),
				.a6(P420F),
				.a7(P421F),
				.a8(P422F),
				.b0(W4100F),
				.b1(W4101F),
				.b2(W4102F),
				.b3(W4110F),
				.b4(W4111F),
				.b5(W4112F),
				.b6(W4120F),
				.b7(W4121F),
				.b8(W4122F),
				.c(c4F001)
);

ninexnine_unit ninexnine_unit_7856(
				.clk(clk),
				.rstn(rstn),
				.a0(P400G),
				.a1(P401G),
				.a2(P402G),
				.a3(P410G),
				.a4(P411G),
				.a5(P412G),
				.a6(P420G),
				.a7(P421G),
				.a8(P422G),
				.b0(W4100G),
				.b1(W4101G),
				.b2(W4102G),
				.b3(W4110G),
				.b4(W4111G),
				.b5(W4112G),
				.b6(W4120G),
				.b7(W4121G),
				.b8(W4122G),
				.c(c4G001)
);

ninexnine_unit ninexnine_unit_7857(
				.clk(clk),
				.rstn(rstn),
				.a0(P400H),
				.a1(P401H),
				.a2(P402H),
				.a3(P410H),
				.a4(P411H),
				.a5(P412H),
				.a6(P420H),
				.a7(P421H),
				.a8(P422H),
				.b0(W4100H),
				.b1(W4101H),
				.b2(W4102H),
				.b3(W4110H),
				.b4(W4111H),
				.b5(W4112H),
				.b6(W4120H),
				.b7(W4121H),
				.b8(W4122H),
				.c(c4H001)
);

ninexnine_unit ninexnine_unit_7858(
				.clk(clk),
				.rstn(rstn),
				.a0(P400I),
				.a1(P401I),
				.a2(P402I),
				.a3(P410I),
				.a4(P411I),
				.a5(P412I),
				.a6(P420I),
				.a7(P421I),
				.a8(P422I),
				.b0(W4100I),
				.b1(W4101I),
				.b2(W4102I),
				.b3(W4110I),
				.b4(W4111I),
				.b5(W4112I),
				.b6(W4120I),
				.b7(W4121I),
				.b8(W4122I),
				.c(c4I001)
);

ninexnine_unit ninexnine_unit_7859(
				.clk(clk),
				.rstn(rstn),
				.a0(P400J),
				.a1(P401J),
				.a2(P402J),
				.a3(P410J),
				.a4(P411J),
				.a5(P412J),
				.a6(P420J),
				.a7(P421J),
				.a8(P422J),
				.b0(W4100J),
				.b1(W4101J),
				.b2(W4102J),
				.b3(W4110J),
				.b4(W4111J),
				.b5(W4112J),
				.b6(W4120J),
				.b7(W4121J),
				.b8(W4122J),
				.c(c4J001)
);

ninexnine_unit ninexnine_unit_7860(
				.clk(clk),
				.rstn(rstn),
				.a0(P400K),
				.a1(P401K),
				.a2(P402K),
				.a3(P410K),
				.a4(P411K),
				.a5(P412K),
				.a6(P420K),
				.a7(P421K),
				.a8(P422K),
				.b0(W4100K),
				.b1(W4101K),
				.b2(W4102K),
				.b3(W4110K),
				.b4(W4111K),
				.b5(W4112K),
				.b6(W4120K),
				.b7(W4121K),
				.b8(W4122K),
				.c(c4K001)
);

ninexnine_unit ninexnine_unit_7861(
				.clk(clk),
				.rstn(rstn),
				.a0(P400L),
				.a1(P401L),
				.a2(P402L),
				.a3(P410L),
				.a4(P411L),
				.a5(P412L),
				.a6(P420L),
				.a7(P421L),
				.a8(P422L),
				.b0(W4100L),
				.b1(W4101L),
				.b2(W4102L),
				.b3(W4110L),
				.b4(W4111L),
				.b5(W4112L),
				.b6(W4120L),
				.b7(W4121L),
				.b8(W4122L),
				.c(c4L001)
);

ninexnine_unit ninexnine_unit_7862(
				.clk(clk),
				.rstn(rstn),
				.a0(P400M),
				.a1(P401M),
				.a2(P402M),
				.a3(P410M),
				.a4(P411M),
				.a5(P412M),
				.a6(P420M),
				.a7(P421M),
				.a8(P422M),
				.b0(W4100M),
				.b1(W4101M),
				.b2(W4102M),
				.b3(W4110M),
				.b4(W4111M),
				.b5(W4112M),
				.b6(W4120M),
				.b7(W4121M),
				.b8(W4122M),
				.c(c4M001)
);

ninexnine_unit ninexnine_unit_7863(
				.clk(clk),
				.rstn(rstn),
				.a0(P400N),
				.a1(P401N),
				.a2(P402N),
				.a3(P410N),
				.a4(P411N),
				.a5(P412N),
				.a6(P420N),
				.a7(P421N),
				.a8(P422N),
				.b0(W4100N),
				.b1(W4101N),
				.b2(W4102N),
				.b3(W4110N),
				.b4(W4111N),
				.b5(W4112N),
				.b6(W4120N),
				.b7(W4121N),
				.b8(W4122N),
				.c(c4N001)
);

ninexnine_unit ninexnine_unit_7864(
				.clk(clk),
				.rstn(rstn),
				.a0(P400O),
				.a1(P401O),
				.a2(P402O),
				.a3(P410O),
				.a4(P411O),
				.a5(P412O),
				.a6(P420O),
				.a7(P421O),
				.a8(P422O),
				.b0(W4100O),
				.b1(W4101O),
				.b2(W4102O),
				.b3(W4110O),
				.b4(W4111O),
				.b5(W4112O),
				.b6(W4120O),
				.b7(W4121O),
				.b8(W4122O),
				.c(c4O001)
);

ninexnine_unit ninexnine_unit_7865(
				.clk(clk),
				.rstn(rstn),
				.a0(P400P),
				.a1(P401P),
				.a2(P402P),
				.a3(P410P),
				.a4(P411P),
				.a5(P412P),
				.a6(P420P),
				.a7(P421P),
				.a8(P422P),
				.b0(W4100P),
				.b1(W4101P),
				.b2(W4102P),
				.b3(W4110P),
				.b4(W4111P),
				.b5(W4112P),
				.b6(W4120P),
				.b7(W4121P),
				.b8(W4122P),
				.c(c4P001)
);

ninexnine_unit ninexnine_unit_7866(
				.clk(clk),
				.rstn(rstn),
				.a0(P400Q),
				.a1(P401Q),
				.a2(P402Q),
				.a3(P410Q),
				.a4(P411Q),
				.a5(P412Q),
				.a6(P420Q),
				.a7(P421Q),
				.a8(P422Q),
				.b0(W4100Q),
				.b1(W4101Q),
				.b2(W4102Q),
				.b3(W4110Q),
				.b4(W4111Q),
				.b5(W4112Q),
				.b6(W4120Q),
				.b7(W4121Q),
				.b8(W4122Q),
				.c(c4Q001)
);

ninexnine_unit ninexnine_unit_7867(
				.clk(clk),
				.rstn(rstn),
				.a0(P400R),
				.a1(P401R),
				.a2(P402R),
				.a3(P410R),
				.a4(P411R),
				.a5(P412R),
				.a6(P420R),
				.a7(P421R),
				.a8(P422R),
				.b0(W4100R),
				.b1(W4101R),
				.b2(W4102R),
				.b3(W4110R),
				.b4(W4111R),
				.b5(W4112R),
				.b6(W4120R),
				.b7(W4121R),
				.b8(W4122R),
				.c(c4R001)
);

ninexnine_unit ninexnine_unit_7868(
				.clk(clk),
				.rstn(rstn),
				.a0(P400S),
				.a1(P401S),
				.a2(P402S),
				.a3(P410S),
				.a4(P411S),
				.a5(P412S),
				.a6(P420S),
				.a7(P421S),
				.a8(P422S),
				.b0(W4100S),
				.b1(W4101S),
				.b2(W4102S),
				.b3(W4110S),
				.b4(W4111S),
				.b5(W4112S),
				.b6(W4120S),
				.b7(W4121S),
				.b8(W4122S),
				.c(c4S001)
);

ninexnine_unit ninexnine_unit_7869(
				.clk(clk),
				.rstn(rstn),
				.a0(P400T),
				.a1(P401T),
				.a2(P402T),
				.a3(P410T),
				.a4(P411T),
				.a5(P412T),
				.a6(P420T),
				.a7(P421T),
				.a8(P422T),
				.b0(W4100T),
				.b1(W4101T),
				.b2(W4102T),
				.b3(W4110T),
				.b4(W4111T),
				.b5(W4112T),
				.b6(W4120T),
				.b7(W4121T),
				.b8(W4122T),
				.c(c4T001)
);

ninexnine_unit ninexnine_unit_7870(
				.clk(clk),
				.rstn(rstn),
				.a0(P400U),
				.a1(P401U),
				.a2(P402U),
				.a3(P410U),
				.a4(P411U),
				.a5(P412U),
				.a6(P420U),
				.a7(P421U),
				.a8(P422U),
				.b0(W4100U),
				.b1(W4101U),
				.b2(W4102U),
				.b3(W4110U),
				.b4(W4111U),
				.b5(W4112U),
				.b6(W4120U),
				.b7(W4121U),
				.b8(W4122U),
				.c(c4U001)
);

ninexnine_unit ninexnine_unit_7871(
				.clk(clk),
				.rstn(rstn),
				.a0(P400V),
				.a1(P401V),
				.a2(P402V),
				.a3(P410V),
				.a4(P411V),
				.a5(P412V),
				.a6(P420V),
				.a7(P421V),
				.a8(P422V),
				.b0(W4100V),
				.b1(W4101V),
				.b2(W4102V),
				.b3(W4110V),
				.b4(W4111V),
				.b5(W4112V),
				.b6(W4120V),
				.b7(W4121V),
				.b8(W4122V),
				.c(c4V001)
);

assign C4001=c40001+c41001+c42001+c43001+c44001+c45001+c46001+c47001+c48001+c49001+c4A001+c4B001+c4C001+c4D001+c4E001+c4F001+c4G001+c4H001+c4I001+c4J001+c4K001+c4L001+c4M001+c4N001+c4O001+c4P001+c4Q001+c4R001+c4S001+c4T001+c4U001+c4V001;
assign A4001=(C4001>=0)?1:0;

assign P5001=A4001;

endmodule
//layer4 done, begain next layer
