module test_layer4(
clk, 
rstn
);
input clk;
input rstn;

wire P4000;
wire P4010;
wire P4020;
wire P4100;
wire P4110;
wire P4120;
wire P4200;
wire P4210;
wire P4220;
wire P4001;
wire P4011;
wire P4021;
wire P4101;
wire P4111;
wire P4121;
wire P4201;
wire P4211;
wire P4221;
wire P4002;
wire P4012;
wire P4022;
wire P4102;
wire P4112;
wire P4122;
wire P4202;
wire P4212;
wire P4222;
wire P4003;
wire P4013;
wire P4023;
wire P4103;
wire P4113;
wire P4123;
wire P4203;
wire P4213;
wire P4223;
wire P4004;
wire P4014;
wire P4024;
wire P4104;
wire P4114;
wire P4124;
wire P4204;
wire P4214;
wire P4224;
wire P4005;
wire P4015;
wire P4025;
wire P4105;
wire P4115;
wire P4125;
wire P4205;
wire P4215;
wire P4225;
wire P4006;
wire P4016;
wire P4026;
wire P4106;
wire P4116;
wire P4126;
wire P4206;
wire P4216;
wire P4226;
wire P4007;
wire P4017;
wire P4027;
wire P4107;
wire P4117;
wire P4127;
wire P4207;
wire P4217;
wire P4227;
wire P4008;
wire P4018;
wire P4028;
wire P4108;
wire P4118;
wire P4128;
wire P4208;
wire P4218;
wire P4228;
wire P4009;
wire P4019;
wire P4029;
wire P4109;
wire P4119;
wire P4129;
wire P4209;
wire P4219;
wire P4229;
wire P400A;
wire P401A;
wire P402A;
wire P410A;
wire P411A;
wire P412A;
wire P420A;
wire P421A;
wire P422A;
wire P400B;
wire P401B;
wire P402B;
wire P410B;
wire P411B;
wire P412B;
wire P420B;
wire P421B;
wire P422B;
wire P400C;
wire P401C;
wire P402C;
wire P410C;
wire P411C;
wire P412C;
wire P420C;
wire P421C;
wire P422C;
wire P400D;
wire P401D;
wire P402D;
wire P410D;
wire P411D;
wire P412D;
wire P420D;
wire P421D;
wire P422D;
wire P400E;
wire P401E;
wire P402E;
wire P410E;
wire P411E;
wire P412E;
wire P420E;
wire P421E;
wire P422E;
wire P400F;
wire P401F;
wire P402F;
wire P410F;
wire P411F;
wire P412F;
wire P420F;
wire P421F;
wire P422F;
wire P400G;
wire P401G;
wire P402G;
wire P410G;
wire P411G;
wire P412G;
wire P420G;
wire P421G;
wire P422G;
wire P400H;
wire P401H;
wire P402H;
wire P410H;
wire P411H;
wire P412H;
wire P420H;
wire P421H;
wire P422H;
wire P400I;
wire P401I;
wire P402I;
wire P410I;
wire P411I;
wire P412I;
wire P420I;
wire P421I;
wire P422I;
wire P400J;
wire P401J;
wire P402J;
wire P410J;
wire P411J;
wire P412J;
wire P420J;
wire P421J;
wire P422J;
wire P400K;
wire P401K;
wire P402K;
wire P410K;
wire P411K;
wire P412K;
wire P420K;
wire P421K;
wire P422K;
wire P400L;
wire P401L;
wire P402L;
wire P410L;
wire P411L;
wire P412L;
wire P420L;
wire P421L;
wire P422L;
wire P400M;
wire P401M;
wire P402M;
wire P410M;
wire P411M;
wire P412M;
wire P420M;
wire P421M;
wire P422M;
wire P400N;
wire P401N;
wire P402N;
wire P410N;
wire P411N;
wire P412N;
wire P420N;
wire P421N;
wire P422N;
wire P400O;
wire P401O;
wire P402O;
wire P410O;
wire P411O;
wire P412O;
wire P420O;
wire P421O;
wire P422O;
wire P400P;
wire P401P;
wire P402P;
wire P410P;
wire P411P;
wire P412P;
wire P420P;
wire P421P;
wire P422P;
wire P400Q;
wire P401Q;
wire P402Q;
wire P410Q;
wire P411Q;
wire P412Q;
wire P420Q;
wire P421Q;
wire P422Q;
wire P400R;
wire P401R;
wire P402R;
wire P410R;
wire P411R;
wire P412R;
wire P420R;
wire P421R;
wire P422R;
wire P400S;
wire P401S;
wire P402S;
wire P410S;
wire P411S;
wire P412S;
wire P420S;
wire P421S;
wire P422S;
wire P400T;
wire P401T;
wire P402T;
wire P410T;
wire P411T;
wire P412T;
wire P420T;
wire P421T;
wire P422T;
wire P400U;
wire P401U;
wire P402U;
wire P410U;
wire P411U;
wire P412U;
wire P420U;
wire P421U;
wire P422U;
wire P400V;
wire P401V;
wire P402V;
wire P410V;
wire P411V;
wire P412V;
wire P420V;
wire P421V;
wire P422V;
wire P5000;
wire P5001;
wire W40000,W40010,W40020,W40100,W40110,W40120,W40200,W40210,W40220;
wire W40001,W40011,W40021,W40101,W40111,W40121,W40201,W40211,W40221;
wire W40002,W40012,W40022,W40102,W40112,W40122,W40202,W40212,W40222;
wire W40003,W40013,W40023,W40103,W40113,W40123,W40203,W40213,W40223;
wire W40004,W40014,W40024,W40104,W40114,W40124,W40204,W40214,W40224;
wire W40005,W40015,W40025,W40105,W40115,W40125,W40205,W40215,W40225;
wire W40006,W40016,W40026,W40106,W40116,W40126,W40206,W40216,W40226;
wire W40007,W40017,W40027,W40107,W40117,W40127,W40207,W40217,W40227;
wire W40008,W40018,W40028,W40108,W40118,W40128,W40208,W40218,W40228;
wire W40009,W40019,W40029,W40109,W40119,W40129,W40209,W40219,W40229;
wire W4000A,W4001A,W4002A,W4010A,W4011A,W4012A,W4020A,W4021A,W4022A;
wire W4000B,W4001B,W4002B,W4010B,W4011B,W4012B,W4020B,W4021B,W4022B;
wire W4000C,W4001C,W4002C,W4010C,W4011C,W4012C,W4020C,W4021C,W4022C;
wire W4000D,W4001D,W4002D,W4010D,W4011D,W4012D,W4020D,W4021D,W4022D;
wire W4000E,W4001E,W4002E,W4010E,W4011E,W4012E,W4020E,W4021E,W4022E;
wire W4000F,W4001F,W4002F,W4010F,W4011F,W4012F,W4020F,W4021F,W4022F;
wire W4000G,W4001G,W4002G,W4010G,W4011G,W4012G,W4020G,W4021G,W4022G;
wire W4000H,W4001H,W4002H,W4010H,W4011H,W4012H,W4020H,W4021H,W4022H;
wire W4000I,W4001I,W4002I,W4010I,W4011I,W4012I,W4020I,W4021I,W4022I;
wire W4000J,W4001J,W4002J,W4010J,W4011J,W4012J,W4020J,W4021J,W4022J;
wire W4000K,W4001K,W4002K,W4010K,W4011K,W4012K,W4020K,W4021K,W4022K;
wire W4000L,W4001L,W4002L,W4010L,W4011L,W4012L,W4020L,W4021L,W4022L;
wire W4000M,W4001M,W4002M,W4010M,W4011M,W4012M,W4020M,W4021M,W4022M;
wire W4000N,W4001N,W4002N,W4010N,W4011N,W4012N,W4020N,W4021N,W4022N;
wire W4000O,W4001O,W4002O,W4010O,W4011O,W4012O,W4020O,W4021O,W4022O;
wire W4000P,W4001P,W4002P,W4010P,W4011P,W4012P,W4020P,W4021P,W4022P;
wire W4000Q,W4001Q,W4002Q,W4010Q,W4011Q,W4012Q,W4020Q,W4021Q,W4022Q;
wire W4000R,W4001R,W4002R,W4010R,W4011R,W4012R,W4020R,W4021R,W4022R;
wire W4000S,W4001S,W4002S,W4010S,W4011S,W4012S,W4020S,W4021S,W4022S;
wire W4000T,W4001T,W4002T,W4010T,W4011T,W4012T,W4020T,W4021T,W4022T;
wire W4000U,W4001U,W4002U,W4010U,W4011U,W4012U,W4020U,W4021U,W4022U;
wire W4000V,W4001V,W4002V,W4010V,W4011V,W4012V,W4020V,W4021V,W4022V;
wire W41000,W41010,W41020,W41100,W41110,W41120,W41200,W41210,W41220;
wire W41001,W41011,W41021,W41101,W41111,W41121,W41201,W41211,W41221;
wire W41002,W41012,W41022,W41102,W41112,W41122,W41202,W41212,W41222;
wire W41003,W41013,W41023,W41103,W41113,W41123,W41203,W41213,W41223;
wire W41004,W41014,W41024,W41104,W41114,W41124,W41204,W41214,W41224;
wire W41005,W41015,W41025,W41105,W41115,W41125,W41205,W41215,W41225;
wire W41006,W41016,W41026,W41106,W41116,W41126,W41206,W41216,W41226;
wire W41007,W41017,W41027,W41107,W41117,W41127,W41207,W41217,W41227;
wire W41008,W41018,W41028,W41108,W41118,W41128,W41208,W41218,W41228;
wire W41009,W41019,W41029,W41109,W41119,W41129,W41209,W41219,W41229;
wire W4100A,W4101A,W4102A,W4110A,W4111A,W4112A,W4120A,W4121A,W4122A;
wire W4100B,W4101B,W4102B,W4110B,W4111B,W4112B,W4120B,W4121B,W4122B;
wire W4100C,W4101C,W4102C,W4110C,W4111C,W4112C,W4120C,W4121C,W4122C;
wire W4100D,W4101D,W4102D,W4110D,W4111D,W4112D,W4120D,W4121D,W4122D;
wire W4100E,W4101E,W4102E,W4110E,W4111E,W4112E,W4120E,W4121E,W4122E;
wire W4100F,W4101F,W4102F,W4110F,W4111F,W4112F,W4120F,W4121F,W4122F;
wire W4100G,W4101G,W4102G,W4110G,W4111G,W4112G,W4120G,W4121G,W4122G;
wire W4100H,W4101H,W4102H,W4110H,W4111H,W4112H,W4120H,W4121H,W4122H;
wire W4100I,W4101I,W4102I,W4110I,W4111I,W4112I,W4120I,W4121I,W4122I;
wire W4100J,W4101J,W4102J,W4110J,W4111J,W4112J,W4120J,W4121J,W4122J;
wire W4100K,W4101K,W4102K,W4110K,W4111K,W4112K,W4120K,W4121K,W4122K;
wire W4100L,W4101L,W4102L,W4110L,W4111L,W4112L,W4120L,W4121L,W4122L;
wire W4100M,W4101M,W4102M,W4110M,W4111M,W4112M,W4120M,W4121M,W4122M;
wire W4100N,W4101N,W4102N,W4110N,W4111N,W4112N,W4120N,W4121N,W4122N;
wire W4100O,W4101O,W4102O,W4110O,W4111O,W4112O,W4120O,W4121O,W4122O;
wire W4100P,W4101P,W4102P,W4110P,W4111P,W4112P,W4120P,W4121P,W4122P;
wire W4100Q,W4101Q,W4102Q,W4110Q,W4111Q,W4112Q,W4120Q,W4121Q,W4122Q;
wire W4100R,W4101R,W4102R,W4110R,W4111R,W4112R,W4120R,W4121R,W4122R;
wire W4100S,W4101S,W4102S,W4110S,W4111S,W4112S,W4120S,W4121S,W4122S;
wire W4100T,W4101T,W4102T,W4110T,W4111T,W4112T,W4120T,W4121T,W4122T;
wire W4100U,W4101U,W4102U,W4110U,W4111U,W4112U,W4120U,W4121U,W4122U;
wire W4100V,W4101V,W4102V,W4110V,W4111V,W4112V,W4120V,W4121V,W4122V;
wire signed [4:0] c40000,c41000,c42000,c43000,c44000,c45000,c46000,c47000,c48000,c49000,c4A000,c4B000,c4C000,c4D000,c4E000,c4F000,c4G000,c4H000,c4I000,c4J000,c4K000,c4L000,c4M000,c4N000,c4O000,c4P000,c4Q000,c4R000,c4S000,c4T000,c4U000,c4V000;
wire signed [4:0] c40001,c41001,c42001,c43001,c44001,c45001,c46001,c47001,c48001,c49001,c4A001,c4B001,c4C001,c4D001,c4E001,c4F001,c4G001,c4H001,c4I001,c4J001,c4K001,c4L001,c4M001,c4N001,c4O001,c4P001,c4Q001,c4R001,c4S001,c4T001,c4U001,c4V001;
wire signed [9:0] C4000;
wire A4000;
wire signed [9:0] C4001;
wire A4001;
DFF_save_fm DFF_P0(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4000));
DFF_save_fm DFF_P1(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4010));
DFF_save_fm DFF_P2(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4020));
DFF_save_fm DFF_P3(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4100));
DFF_save_fm DFF_P4(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4110));
DFF_save_fm DFF_P5(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4120));
DFF_save_fm DFF_P6(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4200));
DFF_save_fm DFF_P7(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4210));
DFF_save_fm DFF_P8(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4220));
DFF_save_fm DFF_P9(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4001));
DFF_save_fm DFF_P10(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4011));
DFF_save_fm DFF_P11(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4021));
DFF_save_fm DFF_P12(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4101));
DFF_save_fm DFF_P13(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4111));
DFF_save_fm DFF_P14(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4121));
DFF_save_fm DFF_P15(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4201));
DFF_save_fm DFF_P16(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4211));
DFF_save_fm DFF_P17(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4221));
DFF_save_fm DFF_P18(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4002));
DFF_save_fm DFF_P19(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4012));
DFF_save_fm DFF_P20(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4022));
DFF_save_fm DFF_P21(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4102));
DFF_save_fm DFF_P22(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4112));
DFF_save_fm DFF_P23(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4122));
DFF_save_fm DFF_P24(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4202));
DFF_save_fm DFF_P25(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4212));
DFF_save_fm DFF_P26(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4222));
DFF_save_fm DFF_P27(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4003));
DFF_save_fm DFF_P28(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4013));
DFF_save_fm DFF_P29(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4023));
DFF_save_fm DFF_P30(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4103));
DFF_save_fm DFF_P31(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4113));
DFF_save_fm DFF_P32(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4123));
DFF_save_fm DFF_P33(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4203));
DFF_save_fm DFF_P34(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4213));
DFF_save_fm DFF_P35(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4223));
DFF_save_fm DFF_P36(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4004));
DFF_save_fm DFF_P37(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4014));
DFF_save_fm DFF_P38(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4024));
DFF_save_fm DFF_P39(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4104));
DFF_save_fm DFF_P40(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4114));
DFF_save_fm DFF_P41(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4124));
DFF_save_fm DFF_P42(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4204));
DFF_save_fm DFF_P43(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4214));
DFF_save_fm DFF_P44(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4224));
DFF_save_fm DFF_P45(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4005));
DFF_save_fm DFF_P46(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4015));
DFF_save_fm DFF_P47(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4025));
DFF_save_fm DFF_P48(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4105));
DFF_save_fm DFF_P49(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4115));
DFF_save_fm DFF_P50(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4125));
DFF_save_fm DFF_P51(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4205));
DFF_save_fm DFF_P52(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4215));
DFF_save_fm DFF_P53(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4225));
DFF_save_fm DFF_P54(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4006));
DFF_save_fm DFF_P55(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4016));
DFF_save_fm DFF_P56(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4026));
DFF_save_fm DFF_P57(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4106));
DFF_save_fm DFF_P58(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4116));
DFF_save_fm DFF_P59(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4126));
DFF_save_fm DFF_P60(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4206));
DFF_save_fm DFF_P61(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4216));
DFF_save_fm DFF_P62(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4226));
DFF_save_fm DFF_P63(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4007));
DFF_save_fm DFF_P64(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4017));
DFF_save_fm DFF_P65(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4027));
DFF_save_fm DFF_P66(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4107));
DFF_save_fm DFF_P67(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4117));
DFF_save_fm DFF_P68(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4127));
DFF_save_fm DFF_P69(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4207));
DFF_save_fm DFF_P70(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4217));
DFF_save_fm DFF_P71(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4227));
DFF_save_fm DFF_P72(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4008));
DFF_save_fm DFF_P73(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4018));
DFF_save_fm DFF_P74(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4028));
DFF_save_fm DFF_P75(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4108));
DFF_save_fm DFF_P76(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4118));
DFF_save_fm DFF_P77(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4128));
DFF_save_fm DFF_P78(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4208));
DFF_save_fm DFF_P79(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4218));
DFF_save_fm DFF_P80(.clk(clk),.rstn(rstn),.reset_value(0),.q(P4228));
DFF_save_fm DFF_P81(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4009));
DFF_save_fm DFF_P82(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4019));
DFF_save_fm DFF_P83(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4029));
DFF_save_fm DFF_P84(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4109));
DFF_save_fm DFF_P85(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4119));
DFF_save_fm DFF_P86(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4129));
DFF_save_fm DFF_P87(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4209));
DFF_save_fm DFF_P88(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4219));
DFF_save_fm DFF_P89(.clk(clk),.rstn(rstn),.reset_value(1),.q(P4229));
DFF_save_fm DFF_P90(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400A));
DFF_save_fm DFF_P91(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401A));
DFF_save_fm DFF_P92(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402A));
DFF_save_fm DFF_P93(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410A));
DFF_save_fm DFF_P94(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411A));
DFF_save_fm DFF_P95(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412A));
DFF_save_fm DFF_P96(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420A));
DFF_save_fm DFF_P97(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421A));
DFF_save_fm DFF_P98(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422A));
DFF_save_fm DFF_P99(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400B));
DFF_save_fm DFF_P100(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401B));
DFF_save_fm DFF_P101(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402B));
DFF_save_fm DFF_P102(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410B));
DFF_save_fm DFF_P103(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411B));
DFF_save_fm DFF_P104(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412B));
DFF_save_fm DFF_P105(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420B));
DFF_save_fm DFF_P106(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421B));
DFF_save_fm DFF_P107(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422B));
DFF_save_fm DFF_P108(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400C));
DFF_save_fm DFF_P109(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401C));
DFF_save_fm DFF_P110(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402C));
DFF_save_fm DFF_P111(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410C));
DFF_save_fm DFF_P112(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411C));
DFF_save_fm DFF_P113(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412C));
DFF_save_fm DFF_P114(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420C));
DFF_save_fm DFF_P115(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421C));
DFF_save_fm DFF_P116(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422C));
DFF_save_fm DFF_P117(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400D));
DFF_save_fm DFF_P118(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401D));
DFF_save_fm DFF_P119(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402D));
DFF_save_fm DFF_P120(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410D));
DFF_save_fm DFF_P121(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411D));
DFF_save_fm DFF_P122(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412D));
DFF_save_fm DFF_P123(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420D));
DFF_save_fm DFF_P124(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421D));
DFF_save_fm DFF_P125(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422D));
DFF_save_fm DFF_P126(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400E));
DFF_save_fm DFF_P127(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401E));
DFF_save_fm DFF_P128(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402E));
DFF_save_fm DFF_P129(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410E));
DFF_save_fm DFF_P130(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411E));
DFF_save_fm DFF_P131(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412E));
DFF_save_fm DFF_P132(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420E));
DFF_save_fm DFF_P133(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421E));
DFF_save_fm DFF_P134(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422E));
DFF_save_fm DFF_P135(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400F));
DFF_save_fm DFF_P136(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401F));
DFF_save_fm DFF_P137(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402F));
DFF_save_fm DFF_P138(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410F));
DFF_save_fm DFF_P139(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411F));
DFF_save_fm DFF_P140(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412F));
DFF_save_fm DFF_P141(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420F));
DFF_save_fm DFF_P142(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421F));
DFF_save_fm DFF_P143(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422F));
DFF_save_fm DFF_P144(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400G));
DFF_save_fm DFF_P145(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401G));
DFF_save_fm DFF_P146(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402G));
DFF_save_fm DFF_P147(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410G));
DFF_save_fm DFF_P148(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411G));
DFF_save_fm DFF_P149(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412G));
DFF_save_fm DFF_P150(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420G));
DFF_save_fm DFF_P151(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421G));
DFF_save_fm DFF_P152(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422G));
DFF_save_fm DFF_P153(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400H));
DFF_save_fm DFF_P154(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401H));
DFF_save_fm DFF_P155(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402H));
DFF_save_fm DFF_P156(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410H));
DFF_save_fm DFF_P157(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411H));
DFF_save_fm DFF_P158(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412H));
DFF_save_fm DFF_P159(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420H));
DFF_save_fm DFF_P160(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421H));
DFF_save_fm DFF_P161(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422H));
DFF_save_fm DFF_P162(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400I));
DFF_save_fm DFF_P163(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401I));
DFF_save_fm DFF_P164(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402I));
DFF_save_fm DFF_P165(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410I));
DFF_save_fm DFF_P166(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411I));
DFF_save_fm DFF_P167(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412I));
DFF_save_fm DFF_P168(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420I));
DFF_save_fm DFF_P169(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421I));
DFF_save_fm DFF_P170(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422I));
DFF_save_fm DFF_P171(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400J));
DFF_save_fm DFF_P172(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401J));
DFF_save_fm DFF_P173(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402J));
DFF_save_fm DFF_P174(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410J));
DFF_save_fm DFF_P175(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411J));
DFF_save_fm DFF_P176(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412J));
DFF_save_fm DFF_P177(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420J));
DFF_save_fm DFF_P178(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421J));
DFF_save_fm DFF_P179(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422J));
DFF_save_fm DFF_P180(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400K));
DFF_save_fm DFF_P181(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401K));
DFF_save_fm DFF_P182(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402K));
DFF_save_fm DFF_P183(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410K));
DFF_save_fm DFF_P184(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411K));
DFF_save_fm DFF_P185(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412K));
DFF_save_fm DFF_P186(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420K));
DFF_save_fm DFF_P187(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421K));
DFF_save_fm DFF_P188(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422K));
DFF_save_fm DFF_P189(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400L));
DFF_save_fm DFF_P190(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401L));
DFF_save_fm DFF_P191(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402L));
DFF_save_fm DFF_P192(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410L));
DFF_save_fm DFF_P193(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411L));
DFF_save_fm DFF_P194(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412L));
DFF_save_fm DFF_P195(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420L));
DFF_save_fm DFF_P196(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421L));
DFF_save_fm DFF_P197(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422L));
DFF_save_fm DFF_P198(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400M));
DFF_save_fm DFF_P199(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401M));
DFF_save_fm DFF_P200(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402M));
DFF_save_fm DFF_P201(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410M));
DFF_save_fm DFF_P202(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411M));
DFF_save_fm DFF_P203(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412M));
DFF_save_fm DFF_P204(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420M));
DFF_save_fm DFF_P205(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421M));
DFF_save_fm DFF_P206(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422M));
DFF_save_fm DFF_P207(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400N));
DFF_save_fm DFF_P208(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401N));
DFF_save_fm DFF_P209(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402N));
DFF_save_fm DFF_P210(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410N));
DFF_save_fm DFF_P211(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411N));
DFF_save_fm DFF_P212(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412N));
DFF_save_fm DFF_P213(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420N));
DFF_save_fm DFF_P214(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421N));
DFF_save_fm DFF_P215(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422N));
DFF_save_fm DFF_P216(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400O));
DFF_save_fm DFF_P217(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401O));
DFF_save_fm DFF_P218(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402O));
DFF_save_fm DFF_P219(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410O));
DFF_save_fm DFF_P220(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411O));
DFF_save_fm DFF_P221(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412O));
DFF_save_fm DFF_P222(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420O));
DFF_save_fm DFF_P223(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421O));
DFF_save_fm DFF_P224(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422O));
DFF_save_fm DFF_P225(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400P));
DFF_save_fm DFF_P226(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401P));
DFF_save_fm DFF_P227(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402P));
DFF_save_fm DFF_P228(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410P));
DFF_save_fm DFF_P229(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411P));
DFF_save_fm DFF_P230(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412P));
DFF_save_fm DFF_P231(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420P));
DFF_save_fm DFF_P232(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421P));
DFF_save_fm DFF_P233(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422P));
DFF_save_fm DFF_P234(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400Q));
DFF_save_fm DFF_P235(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401Q));
DFF_save_fm DFF_P236(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402Q));
DFF_save_fm DFF_P237(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410Q));
DFF_save_fm DFF_P238(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411Q));
DFF_save_fm DFF_P239(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412Q));
DFF_save_fm DFF_P240(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420Q));
DFF_save_fm DFF_P241(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421Q));
DFF_save_fm DFF_P242(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422Q));
DFF_save_fm DFF_P243(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400R));
DFF_save_fm DFF_P244(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401R));
DFF_save_fm DFF_P245(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402R));
DFF_save_fm DFF_P246(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410R));
DFF_save_fm DFF_P247(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411R));
DFF_save_fm DFF_P248(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412R));
DFF_save_fm DFF_P249(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420R));
DFF_save_fm DFF_P250(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421R));
DFF_save_fm DFF_P251(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422R));
DFF_save_fm DFF_P252(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400S));
DFF_save_fm DFF_P253(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401S));
DFF_save_fm DFF_P254(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402S));
DFF_save_fm DFF_P255(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410S));
DFF_save_fm DFF_P256(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411S));
DFF_save_fm DFF_P257(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412S));
DFF_save_fm DFF_P258(.clk(clk),.rstn(rstn),.reset_value(1),.q(P420S));
DFF_save_fm DFF_P259(.clk(clk),.rstn(rstn),.reset_value(0),.q(P421S));
DFF_save_fm DFF_P260(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422S));
DFF_save_fm DFF_P261(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400T));
DFF_save_fm DFF_P262(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401T));
DFF_save_fm DFF_P263(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402T));
DFF_save_fm DFF_P264(.clk(clk),.rstn(rstn),.reset_value(0),.q(P410T));
DFF_save_fm DFF_P265(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411T));
DFF_save_fm DFF_P266(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412T));
DFF_save_fm DFF_P267(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420T));
DFF_save_fm DFF_P268(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421T));
DFF_save_fm DFF_P269(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422T));
DFF_save_fm DFF_P270(.clk(clk),.rstn(rstn),.reset_value(0),.q(P400U));
DFF_save_fm DFF_P271(.clk(clk),.rstn(rstn),.reset_value(1),.q(P401U));
DFF_save_fm DFF_P272(.clk(clk),.rstn(rstn),.reset_value(0),.q(P402U));
DFF_save_fm DFF_P273(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410U));
DFF_save_fm DFF_P274(.clk(clk),.rstn(rstn),.reset_value(0),.q(P411U));
DFF_save_fm DFF_P275(.clk(clk),.rstn(rstn),.reset_value(0),.q(P412U));
DFF_save_fm DFF_P276(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420U));
DFF_save_fm DFF_P277(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421U));
DFF_save_fm DFF_P278(.clk(clk),.rstn(rstn),.reset_value(1),.q(P422U));
DFF_save_fm DFF_P279(.clk(clk),.rstn(rstn),.reset_value(1),.q(P400V));
DFF_save_fm DFF_P280(.clk(clk),.rstn(rstn),.reset_value(0),.q(P401V));
DFF_save_fm DFF_P281(.clk(clk),.rstn(rstn),.reset_value(1),.q(P402V));
DFF_save_fm DFF_P282(.clk(clk),.rstn(rstn),.reset_value(1),.q(P410V));
DFF_save_fm DFF_P283(.clk(clk),.rstn(rstn),.reset_value(1),.q(P411V));
DFF_save_fm DFF_P284(.clk(clk),.rstn(rstn),.reset_value(1),.q(P412V));
DFF_save_fm DFF_P285(.clk(clk),.rstn(rstn),.reset_value(0),.q(P420V));
DFF_save_fm DFF_P286(.clk(clk),.rstn(rstn),.reset_value(1),.q(P421V));
DFF_save_fm DFF_P287(.clk(clk),.rstn(rstn),.reset_value(0),.q(P422V));
DFF_save_fm DFF_W0(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40000));
DFF_save_fm DFF_W1(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40010));
DFF_save_fm DFF_W2(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40020));
DFF_save_fm DFF_W3(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40100));
DFF_save_fm DFF_W4(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40110));
DFF_save_fm DFF_W5(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40120));
DFF_save_fm DFF_W6(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40200));
DFF_save_fm DFF_W7(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40210));
DFF_save_fm DFF_W8(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40220));
DFF_save_fm DFF_W9(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40001));
DFF_save_fm DFF_W10(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40011));
DFF_save_fm DFF_W11(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40021));
DFF_save_fm DFF_W12(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40101));
DFF_save_fm DFF_W13(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40111));
DFF_save_fm DFF_W14(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40121));
DFF_save_fm DFF_W15(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40201));
DFF_save_fm DFF_W16(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40211));
DFF_save_fm DFF_W17(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40221));
DFF_save_fm DFF_W18(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40002));
DFF_save_fm DFF_W19(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40012));
DFF_save_fm DFF_W20(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40022));
DFF_save_fm DFF_W21(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40102));
DFF_save_fm DFF_W22(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40112));
DFF_save_fm DFF_W23(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40122));
DFF_save_fm DFF_W24(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40202));
DFF_save_fm DFF_W25(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40212));
DFF_save_fm DFF_W26(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40222));
DFF_save_fm DFF_W27(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40003));
DFF_save_fm DFF_W28(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40013));
DFF_save_fm DFF_W29(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40023));
DFF_save_fm DFF_W30(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40103));
DFF_save_fm DFF_W31(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40113));
DFF_save_fm DFF_W32(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40123));
DFF_save_fm DFF_W33(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40203));
DFF_save_fm DFF_W34(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40213));
DFF_save_fm DFF_W35(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40223));
DFF_save_fm DFF_W36(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40004));
DFF_save_fm DFF_W37(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40014));
DFF_save_fm DFF_W38(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40024));
DFF_save_fm DFF_W39(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40104));
DFF_save_fm DFF_W40(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40114));
DFF_save_fm DFF_W41(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40124));
DFF_save_fm DFF_W42(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40204));
DFF_save_fm DFF_W43(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40214));
DFF_save_fm DFF_W44(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40224));
DFF_save_fm DFF_W45(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40005));
DFF_save_fm DFF_W46(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40015));
DFF_save_fm DFF_W47(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40025));
DFF_save_fm DFF_W48(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40105));
DFF_save_fm DFF_W49(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40115));
DFF_save_fm DFF_W50(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40125));
DFF_save_fm DFF_W51(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40205));
DFF_save_fm DFF_W52(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40215));
DFF_save_fm DFF_W53(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40225));
DFF_save_fm DFF_W54(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40006));
DFF_save_fm DFF_W55(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40016));
DFF_save_fm DFF_W56(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40026));
DFF_save_fm DFF_W57(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40106));
DFF_save_fm DFF_W58(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40116));
DFF_save_fm DFF_W59(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40126));
DFF_save_fm DFF_W60(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40206));
DFF_save_fm DFF_W61(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40216));
DFF_save_fm DFF_W62(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40226));
DFF_save_fm DFF_W63(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40007));
DFF_save_fm DFF_W64(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40017));
DFF_save_fm DFF_W65(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40027));
DFF_save_fm DFF_W66(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40107));
DFF_save_fm DFF_W67(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40117));
DFF_save_fm DFF_W68(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40127));
DFF_save_fm DFF_W69(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40207));
DFF_save_fm DFF_W70(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40217));
DFF_save_fm DFF_W71(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40227));
DFF_save_fm DFF_W72(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40008));
DFF_save_fm DFF_W73(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40018));
DFF_save_fm DFF_W74(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40028));
DFF_save_fm DFF_W75(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40108));
DFF_save_fm DFF_W76(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40118));
DFF_save_fm DFF_W77(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40128));
DFF_save_fm DFF_W78(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40208));
DFF_save_fm DFF_W79(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40218));
DFF_save_fm DFF_W80(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40228));
DFF_save_fm DFF_W81(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40009));
DFF_save_fm DFF_W82(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40019));
DFF_save_fm DFF_W83(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40029));
DFF_save_fm DFF_W84(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40109));
DFF_save_fm DFF_W85(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40119));
DFF_save_fm DFF_W86(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40129));
DFF_save_fm DFF_W87(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40209));
DFF_save_fm DFF_W88(.clk(clk),.rstn(rstn),.reset_value(1),.q(W40219));
DFF_save_fm DFF_W89(.clk(clk),.rstn(rstn),.reset_value(0),.q(W40229));
DFF_save_fm DFF_W90(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000A));
DFF_save_fm DFF_W91(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001A));
DFF_save_fm DFF_W92(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002A));
DFF_save_fm DFF_W93(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010A));
DFF_save_fm DFF_W94(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011A));
DFF_save_fm DFF_W95(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012A));
DFF_save_fm DFF_W96(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020A));
DFF_save_fm DFF_W97(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021A));
DFF_save_fm DFF_W98(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022A));
DFF_save_fm DFF_W99(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000B));
DFF_save_fm DFF_W100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001B));
DFF_save_fm DFF_W101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002B));
DFF_save_fm DFF_W102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010B));
DFF_save_fm DFF_W103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011B));
DFF_save_fm DFF_W104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012B));
DFF_save_fm DFF_W105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020B));
DFF_save_fm DFF_W106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021B));
DFF_save_fm DFF_W107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022B));
DFF_save_fm DFF_W108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000C));
DFF_save_fm DFF_W109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001C));
DFF_save_fm DFF_W110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002C));
DFF_save_fm DFF_W111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010C));
DFF_save_fm DFF_W112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011C));
DFF_save_fm DFF_W113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012C));
DFF_save_fm DFF_W114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020C));
DFF_save_fm DFF_W115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021C));
DFF_save_fm DFF_W116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022C));
DFF_save_fm DFF_W117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000D));
DFF_save_fm DFF_W118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001D));
DFF_save_fm DFF_W119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002D));
DFF_save_fm DFF_W120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010D));
DFF_save_fm DFF_W121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011D));
DFF_save_fm DFF_W122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012D));
DFF_save_fm DFF_W123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020D));
DFF_save_fm DFF_W124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021D));
DFF_save_fm DFF_W125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022D));
DFF_save_fm DFF_W126(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000E));
DFF_save_fm DFF_W127(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001E));
DFF_save_fm DFF_W128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002E));
DFF_save_fm DFF_W129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010E));
DFF_save_fm DFF_W130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011E));
DFF_save_fm DFF_W131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012E));
DFF_save_fm DFF_W132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020E));
DFF_save_fm DFF_W133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021E));
DFF_save_fm DFF_W134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022E));
DFF_save_fm DFF_W135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000F));
DFF_save_fm DFF_W136(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001F));
DFF_save_fm DFF_W137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002F));
DFF_save_fm DFF_W138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010F));
DFF_save_fm DFF_W139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011F));
DFF_save_fm DFF_W140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012F));
DFF_save_fm DFF_W141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020F));
DFF_save_fm DFF_W142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021F));
DFF_save_fm DFF_W143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022F));
DFF_save_fm DFF_W144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000G));
DFF_save_fm DFF_W145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001G));
DFF_save_fm DFF_W146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002G));
DFF_save_fm DFF_W147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010G));
DFF_save_fm DFF_W148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011G));
DFF_save_fm DFF_W149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012G));
DFF_save_fm DFF_W150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020G));
DFF_save_fm DFF_W151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021G));
DFF_save_fm DFF_W152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022G));
DFF_save_fm DFF_W153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000H));
DFF_save_fm DFF_W154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001H));
DFF_save_fm DFF_W155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002H));
DFF_save_fm DFF_W156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010H));
DFF_save_fm DFF_W157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011H));
DFF_save_fm DFF_W158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012H));
DFF_save_fm DFF_W159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020H));
DFF_save_fm DFF_W160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021H));
DFF_save_fm DFF_W161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022H));
DFF_save_fm DFF_W162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000I));
DFF_save_fm DFF_W163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001I));
DFF_save_fm DFF_W164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002I));
DFF_save_fm DFF_W165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010I));
DFF_save_fm DFF_W166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011I));
DFF_save_fm DFF_W167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012I));
DFF_save_fm DFF_W168(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020I));
DFF_save_fm DFF_W169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021I));
DFF_save_fm DFF_W170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022I));
DFF_save_fm DFF_W171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000J));
DFF_save_fm DFF_W172(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001J));
DFF_save_fm DFF_W173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002J));
DFF_save_fm DFF_W174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010J));
DFF_save_fm DFF_W175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011J));
DFF_save_fm DFF_W176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012J));
DFF_save_fm DFF_W177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020J));
DFF_save_fm DFF_W178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021J));
DFF_save_fm DFF_W179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022J));
DFF_save_fm DFF_W180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000K));
DFF_save_fm DFF_W181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001K));
DFF_save_fm DFF_W182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002K));
DFF_save_fm DFF_W183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010K));
DFF_save_fm DFF_W184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011K));
DFF_save_fm DFF_W185(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012K));
DFF_save_fm DFF_W186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020K));
DFF_save_fm DFF_W187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021K));
DFF_save_fm DFF_W188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022K));
DFF_save_fm DFF_W189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000L));
DFF_save_fm DFF_W190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001L));
DFF_save_fm DFF_W191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002L));
DFF_save_fm DFF_W192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010L));
DFF_save_fm DFF_W193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011L));
DFF_save_fm DFF_W194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012L));
DFF_save_fm DFF_W195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020L));
DFF_save_fm DFF_W196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021L));
DFF_save_fm DFF_W197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022L));
DFF_save_fm DFF_W198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000M));
DFF_save_fm DFF_W199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001M));
DFF_save_fm DFF_W200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002M));
DFF_save_fm DFF_W201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010M));
DFF_save_fm DFF_W202(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011M));
DFF_save_fm DFF_W203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012M));
DFF_save_fm DFF_W204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020M));
DFF_save_fm DFF_W205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021M));
DFF_save_fm DFF_W206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022M));
DFF_save_fm DFF_W207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000N));
DFF_save_fm DFF_W208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001N));
DFF_save_fm DFF_W209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002N));
DFF_save_fm DFF_W210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010N));
DFF_save_fm DFF_W211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011N));
DFF_save_fm DFF_W212(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012N));
DFF_save_fm DFF_W213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020N));
DFF_save_fm DFF_W214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021N));
DFF_save_fm DFF_W215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022N));
DFF_save_fm DFF_W216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000O));
DFF_save_fm DFF_W217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001O));
DFF_save_fm DFF_W218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002O));
DFF_save_fm DFF_W219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010O));
DFF_save_fm DFF_W220(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011O));
DFF_save_fm DFF_W221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012O));
DFF_save_fm DFF_W222(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020O));
DFF_save_fm DFF_W223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021O));
DFF_save_fm DFF_W224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022O));
DFF_save_fm DFF_W225(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000P));
DFF_save_fm DFF_W226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001P));
DFF_save_fm DFF_W227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002P));
DFF_save_fm DFF_W228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010P));
DFF_save_fm DFF_W229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011P));
DFF_save_fm DFF_W230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4012P));
DFF_save_fm DFF_W231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020P));
DFF_save_fm DFF_W232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021P));
DFF_save_fm DFF_W233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022P));
DFF_save_fm DFF_W234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000Q));
DFF_save_fm DFF_W235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001Q));
DFF_save_fm DFF_W236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002Q));
DFF_save_fm DFF_W237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010Q));
DFF_save_fm DFF_W238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011Q));
DFF_save_fm DFF_W239(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012Q));
DFF_save_fm DFF_W240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4020Q));
DFF_save_fm DFF_W241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021Q));
DFF_save_fm DFF_W242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022Q));
DFF_save_fm DFF_W243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000R));
DFF_save_fm DFF_W244(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001R));
DFF_save_fm DFF_W245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002R));
DFF_save_fm DFF_W246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010R));
DFF_save_fm DFF_W247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011R));
DFF_save_fm DFF_W248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012R));
DFF_save_fm DFF_W249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020R));
DFF_save_fm DFF_W250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021R));
DFF_save_fm DFF_W251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4022R));
DFF_save_fm DFF_W252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000S));
DFF_save_fm DFF_W253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001S));
DFF_save_fm DFF_W254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002S));
DFF_save_fm DFF_W255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010S));
DFF_save_fm DFF_W256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011S));
DFF_save_fm DFF_W257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012S));
DFF_save_fm DFF_W258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020S));
DFF_save_fm DFF_W259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021S));
DFF_save_fm DFF_W260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022S));
DFF_save_fm DFF_W261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4000T));
DFF_save_fm DFF_W262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001T));
DFF_save_fm DFF_W263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002T));
DFF_save_fm DFF_W264(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010T));
DFF_save_fm DFF_W265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4011T));
DFF_save_fm DFF_W266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012T));
DFF_save_fm DFF_W267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020T));
DFF_save_fm DFF_W268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021T));
DFF_save_fm DFF_W269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022T));
DFF_save_fm DFF_W270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000U));
DFF_save_fm DFF_W271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4001U));
DFF_save_fm DFF_W272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4002U));
DFF_save_fm DFF_W273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4010U));
DFF_save_fm DFF_W274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011U));
DFF_save_fm DFF_W275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012U));
DFF_save_fm DFF_W276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020U));
DFF_save_fm DFF_W277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4021U));
DFF_save_fm DFF_W278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022U));
DFF_save_fm DFF_W279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4000V));
DFF_save_fm DFF_W280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4001V));
DFF_save_fm DFF_W281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4002V));
DFF_save_fm DFF_W282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4010V));
DFF_save_fm DFF_W283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4011V));
DFF_save_fm DFF_W284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4012V));
DFF_save_fm DFF_W285(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4020V));
DFF_save_fm DFF_W286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4021V));
DFF_save_fm DFF_W287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4022V));
DFF_save_fm DFF_W288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41000));
DFF_save_fm DFF_W289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41010));
DFF_save_fm DFF_W290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41020));
DFF_save_fm DFF_W291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41100));
DFF_save_fm DFF_W292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41110));
DFF_save_fm DFF_W293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41120));
DFF_save_fm DFF_W294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41200));
DFF_save_fm DFF_W295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41210));
DFF_save_fm DFF_W296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41220));
DFF_save_fm DFF_W297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41001));
DFF_save_fm DFF_W298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41011));
DFF_save_fm DFF_W299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41021));
DFF_save_fm DFF_W300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41101));
DFF_save_fm DFF_W301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41111));
DFF_save_fm DFF_W302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41121));
DFF_save_fm DFF_W303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41201));
DFF_save_fm DFF_W304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41211));
DFF_save_fm DFF_W305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41221));
DFF_save_fm DFF_W306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41002));
DFF_save_fm DFF_W307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41012));
DFF_save_fm DFF_W308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41022));
DFF_save_fm DFF_W309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41102));
DFF_save_fm DFF_W310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41112));
DFF_save_fm DFF_W311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41122));
DFF_save_fm DFF_W312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41202));
DFF_save_fm DFF_W313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41212));
DFF_save_fm DFF_W314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41222));
DFF_save_fm DFF_W315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41003));
DFF_save_fm DFF_W316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41013));
DFF_save_fm DFF_W317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41023));
DFF_save_fm DFF_W318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41103));
DFF_save_fm DFF_W319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41113));
DFF_save_fm DFF_W320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41123));
DFF_save_fm DFF_W321(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41203));
DFF_save_fm DFF_W322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41213));
DFF_save_fm DFF_W323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41223));
DFF_save_fm DFF_W324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41004));
DFF_save_fm DFF_W325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41014));
DFF_save_fm DFF_W326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41024));
DFF_save_fm DFF_W327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41104));
DFF_save_fm DFF_W328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41114));
DFF_save_fm DFF_W329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41124));
DFF_save_fm DFF_W330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41204));
DFF_save_fm DFF_W331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41214));
DFF_save_fm DFF_W332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41224));
DFF_save_fm DFF_W333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41005));
DFF_save_fm DFF_W334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41015));
DFF_save_fm DFF_W335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41025));
DFF_save_fm DFF_W336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41105));
DFF_save_fm DFF_W337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41115));
DFF_save_fm DFF_W338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41125));
DFF_save_fm DFF_W339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41205));
DFF_save_fm DFF_W340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41215));
DFF_save_fm DFF_W341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41225));
DFF_save_fm DFF_W342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41006));
DFF_save_fm DFF_W343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41016));
DFF_save_fm DFF_W344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41026));
DFF_save_fm DFF_W345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41106));
DFF_save_fm DFF_W346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41116));
DFF_save_fm DFF_W347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41126));
DFF_save_fm DFF_W348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41206));
DFF_save_fm DFF_W349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41216));
DFF_save_fm DFF_W350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41226));
DFF_save_fm DFF_W351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41007));
DFF_save_fm DFF_W352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41017));
DFF_save_fm DFF_W353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41027));
DFF_save_fm DFF_W354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41107));
DFF_save_fm DFF_W355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41117));
DFF_save_fm DFF_W356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41127));
DFF_save_fm DFF_W357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41207));
DFF_save_fm DFF_W358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41217));
DFF_save_fm DFF_W359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41227));
DFF_save_fm DFF_W360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41008));
DFF_save_fm DFF_W361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41018));
DFF_save_fm DFF_W362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41028));
DFF_save_fm DFF_W363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41108));
DFF_save_fm DFF_W364(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41118));
DFF_save_fm DFF_W365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41128));
DFF_save_fm DFF_W366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41208));
DFF_save_fm DFF_W367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41218));
DFF_save_fm DFF_W368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41228));
DFF_save_fm DFF_W369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41009));
DFF_save_fm DFF_W370(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41019));
DFF_save_fm DFF_W371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41029));
DFF_save_fm DFF_W372(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41109));
DFF_save_fm DFF_W373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W41119));
DFF_save_fm DFF_W374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41129));
DFF_save_fm DFF_W375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41209));
DFF_save_fm DFF_W376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41219));
DFF_save_fm DFF_W377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W41229));
DFF_save_fm DFF_W378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100A));
DFF_save_fm DFF_W379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101A));
DFF_save_fm DFF_W380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102A));
DFF_save_fm DFF_W381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110A));
DFF_save_fm DFF_W382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111A));
DFF_save_fm DFF_W383(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112A));
DFF_save_fm DFF_W384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120A));
DFF_save_fm DFF_W385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121A));
DFF_save_fm DFF_W386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122A));
DFF_save_fm DFF_W387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100B));
DFF_save_fm DFF_W388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101B));
DFF_save_fm DFF_W389(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102B));
DFF_save_fm DFF_W390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110B));
DFF_save_fm DFF_W391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111B));
DFF_save_fm DFF_W392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112B));
DFF_save_fm DFF_W393(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120B));
DFF_save_fm DFF_W394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121B));
DFF_save_fm DFF_W395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122B));
DFF_save_fm DFF_W396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100C));
DFF_save_fm DFF_W397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101C));
DFF_save_fm DFF_W398(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102C));
DFF_save_fm DFF_W399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110C));
DFF_save_fm DFF_W400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111C));
DFF_save_fm DFF_W401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112C));
DFF_save_fm DFF_W402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120C));
DFF_save_fm DFF_W403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121C));
DFF_save_fm DFF_W404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122C));
DFF_save_fm DFF_W405(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100D));
DFF_save_fm DFF_W406(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101D));
DFF_save_fm DFF_W407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102D));
DFF_save_fm DFF_W408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110D));
DFF_save_fm DFF_W409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111D));
DFF_save_fm DFF_W410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112D));
DFF_save_fm DFF_W411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120D));
DFF_save_fm DFF_W412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121D));
DFF_save_fm DFF_W413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122D));
DFF_save_fm DFF_W414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100E));
DFF_save_fm DFF_W415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101E));
DFF_save_fm DFF_W416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102E));
DFF_save_fm DFF_W417(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110E));
DFF_save_fm DFF_W418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111E));
DFF_save_fm DFF_W419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112E));
DFF_save_fm DFF_W420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120E));
DFF_save_fm DFF_W421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121E));
DFF_save_fm DFF_W422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122E));
DFF_save_fm DFF_W423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100F));
DFF_save_fm DFF_W424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101F));
DFF_save_fm DFF_W425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102F));
DFF_save_fm DFF_W426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110F));
DFF_save_fm DFF_W427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111F));
DFF_save_fm DFF_W428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112F));
DFF_save_fm DFF_W429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120F));
DFF_save_fm DFF_W430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121F));
DFF_save_fm DFF_W431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122F));
DFF_save_fm DFF_W432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100G));
DFF_save_fm DFF_W433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101G));
DFF_save_fm DFF_W434(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102G));
DFF_save_fm DFF_W435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110G));
DFF_save_fm DFF_W436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111G));
DFF_save_fm DFF_W437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112G));
DFF_save_fm DFF_W438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120G));
DFF_save_fm DFF_W439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121G));
DFF_save_fm DFF_W440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122G));
DFF_save_fm DFF_W441(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100H));
DFF_save_fm DFF_W442(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101H));
DFF_save_fm DFF_W443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102H));
DFF_save_fm DFF_W444(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110H));
DFF_save_fm DFF_W445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111H));
DFF_save_fm DFF_W446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112H));
DFF_save_fm DFF_W447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120H));
DFF_save_fm DFF_W448(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121H));
DFF_save_fm DFF_W449(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122H));
DFF_save_fm DFF_W450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100I));
DFF_save_fm DFF_W451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101I));
DFF_save_fm DFF_W452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102I));
DFF_save_fm DFF_W453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110I));
DFF_save_fm DFF_W454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111I));
DFF_save_fm DFF_W455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112I));
DFF_save_fm DFF_W456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120I));
DFF_save_fm DFF_W457(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121I));
DFF_save_fm DFF_W458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122I));
DFF_save_fm DFF_W459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100J));
DFF_save_fm DFF_W460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101J));
DFF_save_fm DFF_W461(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102J));
DFF_save_fm DFF_W462(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110J));
DFF_save_fm DFF_W463(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111J));
DFF_save_fm DFF_W464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112J));
DFF_save_fm DFF_W465(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120J));
DFF_save_fm DFF_W466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121J));
DFF_save_fm DFF_W467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122J));
DFF_save_fm DFF_W468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100K));
DFF_save_fm DFF_W469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101K));
DFF_save_fm DFF_W470(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102K));
DFF_save_fm DFF_W471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110K));
DFF_save_fm DFF_W472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111K));
DFF_save_fm DFF_W473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112K));
DFF_save_fm DFF_W474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120K));
DFF_save_fm DFF_W475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121K));
DFF_save_fm DFF_W476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122K));
DFF_save_fm DFF_W477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100L));
DFF_save_fm DFF_W478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101L));
DFF_save_fm DFF_W479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102L));
DFF_save_fm DFF_W480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110L));
DFF_save_fm DFF_W481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111L));
DFF_save_fm DFF_W482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112L));
DFF_save_fm DFF_W483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120L));
DFF_save_fm DFF_W484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121L));
DFF_save_fm DFF_W485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122L));
DFF_save_fm DFF_W486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100M));
DFF_save_fm DFF_W487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101M));
DFF_save_fm DFF_W488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102M));
DFF_save_fm DFF_W489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110M));
DFF_save_fm DFF_W490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111M));
DFF_save_fm DFF_W491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112M));
DFF_save_fm DFF_W492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120M));
DFF_save_fm DFF_W493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121M));
DFF_save_fm DFF_W494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122M));
DFF_save_fm DFF_W495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100N));
DFF_save_fm DFF_W496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101N));
DFF_save_fm DFF_W497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102N));
DFF_save_fm DFF_W498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110N));
DFF_save_fm DFF_W499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111N));
DFF_save_fm DFF_W500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112N));
DFF_save_fm DFF_W501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120N));
DFF_save_fm DFF_W502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121N));
DFF_save_fm DFF_W503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122N));
DFF_save_fm DFF_W504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100O));
DFF_save_fm DFF_W505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101O));
DFF_save_fm DFF_W506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102O));
DFF_save_fm DFF_W507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110O));
DFF_save_fm DFF_W508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111O));
DFF_save_fm DFF_W509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112O));
DFF_save_fm DFF_W510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120O));
DFF_save_fm DFF_W511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121O));
DFF_save_fm DFF_W512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122O));
DFF_save_fm DFF_W513(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100P));
DFF_save_fm DFF_W514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101P));
DFF_save_fm DFF_W515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4102P));
DFF_save_fm DFF_W516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110P));
DFF_save_fm DFF_W517(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111P));
DFF_save_fm DFF_W518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112P));
DFF_save_fm DFF_W519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120P));
DFF_save_fm DFF_W520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121P));
DFF_save_fm DFF_W521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122P));
DFF_save_fm DFF_W522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100Q));
DFF_save_fm DFF_W523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101Q));
DFF_save_fm DFF_W524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102Q));
DFF_save_fm DFF_W525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110Q));
DFF_save_fm DFF_W526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111Q));
DFF_save_fm DFF_W527(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112Q));
DFF_save_fm DFF_W528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120Q));
DFF_save_fm DFF_W529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121Q));
DFF_save_fm DFF_W530(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122Q));
DFF_save_fm DFF_W531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100R));
DFF_save_fm DFF_W532(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101R));
DFF_save_fm DFF_W533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102R));
DFF_save_fm DFF_W534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110R));
DFF_save_fm DFF_W535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111R));
DFF_save_fm DFF_W536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112R));
DFF_save_fm DFF_W537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4120R));
DFF_save_fm DFF_W538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4121R));
DFF_save_fm DFF_W539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122R));
DFF_save_fm DFF_W540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100S));
DFF_save_fm DFF_W541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101S));
DFF_save_fm DFF_W542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102S));
DFF_save_fm DFF_W543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110S));
DFF_save_fm DFF_W544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111S));
DFF_save_fm DFF_W545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112S));
DFF_save_fm DFF_W546(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120S));
DFF_save_fm DFF_W547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121S));
DFF_save_fm DFF_W548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122S));
DFF_save_fm DFF_W549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100T));
DFF_save_fm DFF_W550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101T));
DFF_save_fm DFF_W551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102T));
DFF_save_fm DFF_W552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110T));
DFF_save_fm DFF_W553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111T));
DFF_save_fm DFF_W554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4112T));
DFF_save_fm DFF_W555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120T));
DFF_save_fm DFF_W556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121T));
DFF_save_fm DFF_W557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122T));
DFF_save_fm DFF_W558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4100U));
DFF_save_fm DFF_W559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4101U));
DFF_save_fm DFF_W560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102U));
DFF_save_fm DFF_W561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4110U));
DFF_save_fm DFF_W562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4111U));
DFF_save_fm DFF_W563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112U));
DFF_save_fm DFF_W564(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120U));
DFF_save_fm DFF_W565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121U));
DFF_save_fm DFF_W566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4122U));
DFF_save_fm DFF_W567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4100V));
DFF_save_fm DFF_W568(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4101V));
DFF_save_fm DFF_W569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4102V));
DFF_save_fm DFF_W570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W4110V));
DFF_save_fm DFF_W571(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4111V));
DFF_save_fm DFF_W572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4112V));
DFF_save_fm DFF_W573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4120V));
DFF_save_fm DFF_W574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4121V));
DFF_save_fm DFF_W575(.clk(clk),.rstn(rstn),.reset_value(1),.q(W4122V));
ninexnine_unit ninexnine_unit_0(
				.clk(clk),
				.rstn(rstn),
				.a0(P4000),
				.a1(P4010),
				.a2(P4020),
				.a3(P4100),
				.a4(P4110),
				.a5(P4120),
				.a6(P4200),
				.a7(P4210),
				.a8(P4220),
				.b0(W40000),
				.b1(W40010),
				.b2(W40020),
				.b3(W40100),
				.b4(W40110),
				.b5(W40120),
				.b6(W40200),
				.b7(W40210),
				.b8(W40220),
				.c(c40000)
);

ninexnine_unit ninexnine_unit_1(
				.clk(clk),
				.rstn(rstn),
				.a0(P4001),
				.a1(P4011),
				.a2(P4021),
				.a3(P4101),
				.a4(P4111),
				.a5(P4121),
				.a6(P4201),
				.a7(P4211),
				.a8(P4221),
				.b0(W40001),
				.b1(W40011),
				.b2(W40021),
				.b3(W40101),
				.b4(W40111),
				.b5(W40121),
				.b6(W40201),
				.b7(W40211),
				.b8(W40221),
				.c(c41000)
);

ninexnine_unit ninexnine_unit_2(
				.clk(clk),
				.rstn(rstn),
				.a0(P4002),
				.a1(P4012),
				.a2(P4022),
				.a3(P4102),
				.a4(P4112),
				.a5(P4122),
				.a6(P4202),
				.a7(P4212),
				.a8(P4222),
				.b0(W40002),
				.b1(W40012),
				.b2(W40022),
				.b3(W40102),
				.b4(W40112),
				.b5(W40122),
				.b6(W40202),
				.b7(W40212),
				.b8(W40222),
				.c(c42000)
);

ninexnine_unit ninexnine_unit_3(
				.clk(clk),
				.rstn(rstn),
				.a0(P4003),
				.a1(P4013),
				.a2(P4023),
				.a3(P4103),
				.a4(P4113),
				.a5(P4123),
				.a6(P4203),
				.a7(P4213),
				.a8(P4223),
				.b0(W40003),
				.b1(W40013),
				.b2(W40023),
				.b3(W40103),
				.b4(W40113),
				.b5(W40123),
				.b6(W40203),
				.b7(W40213),
				.b8(W40223),
				.c(c43000)
);

ninexnine_unit ninexnine_unit_4(
				.clk(clk),
				.rstn(rstn),
				.a0(P4004),
				.a1(P4014),
				.a2(P4024),
				.a3(P4104),
				.a4(P4114),
				.a5(P4124),
				.a6(P4204),
				.a7(P4214),
				.a8(P4224),
				.b0(W40004),
				.b1(W40014),
				.b2(W40024),
				.b3(W40104),
				.b4(W40114),
				.b5(W40124),
				.b6(W40204),
				.b7(W40214),
				.b8(W40224),
				.c(c44000)
);

ninexnine_unit ninexnine_unit_5(
				.clk(clk),
				.rstn(rstn),
				.a0(P4005),
				.a1(P4015),
				.a2(P4025),
				.a3(P4105),
				.a4(P4115),
				.a5(P4125),
				.a6(P4205),
				.a7(P4215),
				.a8(P4225),
				.b0(W40005),
				.b1(W40015),
				.b2(W40025),
				.b3(W40105),
				.b4(W40115),
				.b5(W40125),
				.b6(W40205),
				.b7(W40215),
				.b8(W40225),
				.c(c45000)
);

ninexnine_unit ninexnine_unit_6(
				.clk(clk),
				.rstn(rstn),
				.a0(P4006),
				.a1(P4016),
				.a2(P4026),
				.a3(P4106),
				.a4(P4116),
				.a5(P4126),
				.a6(P4206),
				.a7(P4216),
				.a8(P4226),
				.b0(W40006),
				.b1(W40016),
				.b2(W40026),
				.b3(W40106),
				.b4(W40116),
				.b5(W40126),
				.b6(W40206),
				.b7(W40216),
				.b8(W40226),
				.c(c46000)
);

ninexnine_unit ninexnine_unit_7(
				.clk(clk),
				.rstn(rstn),
				.a0(P4007),
				.a1(P4017),
				.a2(P4027),
				.a3(P4107),
				.a4(P4117),
				.a5(P4127),
				.a6(P4207),
				.a7(P4217),
				.a8(P4227),
				.b0(W40007),
				.b1(W40017),
				.b2(W40027),
				.b3(W40107),
				.b4(W40117),
				.b5(W40127),
				.b6(W40207),
				.b7(W40217),
				.b8(W40227),
				.c(c47000)
);

ninexnine_unit ninexnine_unit_8(
				.clk(clk),
				.rstn(rstn),
				.a0(P4008),
				.a1(P4018),
				.a2(P4028),
				.a3(P4108),
				.a4(P4118),
				.a5(P4128),
				.a6(P4208),
				.a7(P4218),
				.a8(P4228),
				.b0(W40008),
				.b1(W40018),
				.b2(W40028),
				.b3(W40108),
				.b4(W40118),
				.b5(W40128),
				.b6(W40208),
				.b7(W40218),
				.b8(W40228),
				.c(c48000)
);

ninexnine_unit ninexnine_unit_9(
				.clk(clk),
				.rstn(rstn),
				.a0(P4009),
				.a1(P4019),
				.a2(P4029),
				.a3(P4109),
				.a4(P4119),
				.a5(P4129),
				.a6(P4209),
				.a7(P4219),
				.a8(P4229),
				.b0(W40009),
				.b1(W40019),
				.b2(W40029),
				.b3(W40109),
				.b4(W40119),
				.b5(W40129),
				.b6(W40209),
				.b7(W40219),
				.b8(W40229),
				.c(c49000)
);

ninexnine_unit ninexnine_unit_10(
				.clk(clk),
				.rstn(rstn),
				.a0(P400A),
				.a1(P401A),
				.a2(P402A),
				.a3(P410A),
				.a4(P411A),
				.a5(P412A),
				.a6(P420A),
				.a7(P421A),
				.a8(P422A),
				.b0(W4000A),
				.b1(W4001A),
				.b2(W4002A),
				.b3(W4010A),
				.b4(W4011A),
				.b5(W4012A),
				.b6(W4020A),
				.b7(W4021A),
				.b8(W4022A),
				.c(c4A000)
);

ninexnine_unit ninexnine_unit_11(
				.clk(clk),
				.rstn(rstn),
				.a0(P400B),
				.a1(P401B),
				.a2(P402B),
				.a3(P410B),
				.a4(P411B),
				.a5(P412B),
				.a6(P420B),
				.a7(P421B),
				.a8(P422B),
				.b0(W4000B),
				.b1(W4001B),
				.b2(W4002B),
				.b3(W4010B),
				.b4(W4011B),
				.b5(W4012B),
				.b6(W4020B),
				.b7(W4021B),
				.b8(W4022B),
				.c(c4B000)
);

ninexnine_unit ninexnine_unit_12(
				.clk(clk),
				.rstn(rstn),
				.a0(P400C),
				.a1(P401C),
				.a2(P402C),
				.a3(P410C),
				.a4(P411C),
				.a5(P412C),
				.a6(P420C),
				.a7(P421C),
				.a8(P422C),
				.b0(W4000C),
				.b1(W4001C),
				.b2(W4002C),
				.b3(W4010C),
				.b4(W4011C),
				.b5(W4012C),
				.b6(W4020C),
				.b7(W4021C),
				.b8(W4022C),
				.c(c4C000)
);

ninexnine_unit ninexnine_unit_13(
				.clk(clk),
				.rstn(rstn),
				.a0(P400D),
				.a1(P401D),
				.a2(P402D),
				.a3(P410D),
				.a4(P411D),
				.a5(P412D),
				.a6(P420D),
				.a7(P421D),
				.a8(P422D),
				.b0(W4000D),
				.b1(W4001D),
				.b2(W4002D),
				.b3(W4010D),
				.b4(W4011D),
				.b5(W4012D),
				.b6(W4020D),
				.b7(W4021D),
				.b8(W4022D),
				.c(c4D000)
);

ninexnine_unit ninexnine_unit_14(
				.clk(clk),
				.rstn(rstn),
				.a0(P400E),
				.a1(P401E),
				.a2(P402E),
				.a3(P410E),
				.a4(P411E),
				.a5(P412E),
				.a6(P420E),
				.a7(P421E),
				.a8(P422E),
				.b0(W4000E),
				.b1(W4001E),
				.b2(W4002E),
				.b3(W4010E),
				.b4(W4011E),
				.b5(W4012E),
				.b6(W4020E),
				.b7(W4021E),
				.b8(W4022E),
				.c(c4E000)
);

ninexnine_unit ninexnine_unit_15(
				.clk(clk),
				.rstn(rstn),
				.a0(P400F),
				.a1(P401F),
				.a2(P402F),
				.a3(P410F),
				.a4(P411F),
				.a5(P412F),
				.a6(P420F),
				.a7(P421F),
				.a8(P422F),
				.b0(W4000F),
				.b1(W4001F),
				.b2(W4002F),
				.b3(W4010F),
				.b4(W4011F),
				.b5(W4012F),
				.b6(W4020F),
				.b7(W4021F),
				.b8(W4022F),
				.c(c4F000)
);

ninexnine_unit ninexnine_unit_16(
				.clk(clk),
				.rstn(rstn),
				.a0(P400G),
				.a1(P401G),
				.a2(P402G),
				.a3(P410G),
				.a4(P411G),
				.a5(P412G),
				.a6(P420G),
				.a7(P421G),
				.a8(P422G),
				.b0(W4000G),
				.b1(W4001G),
				.b2(W4002G),
				.b3(W4010G),
				.b4(W4011G),
				.b5(W4012G),
				.b6(W4020G),
				.b7(W4021G),
				.b8(W4022G),
				.c(c4G000)
);

ninexnine_unit ninexnine_unit_17(
				.clk(clk),
				.rstn(rstn),
				.a0(P400H),
				.a1(P401H),
				.a2(P402H),
				.a3(P410H),
				.a4(P411H),
				.a5(P412H),
				.a6(P420H),
				.a7(P421H),
				.a8(P422H),
				.b0(W4000H),
				.b1(W4001H),
				.b2(W4002H),
				.b3(W4010H),
				.b4(W4011H),
				.b5(W4012H),
				.b6(W4020H),
				.b7(W4021H),
				.b8(W4022H),
				.c(c4H000)
);

ninexnine_unit ninexnine_unit_18(
				.clk(clk),
				.rstn(rstn),
				.a0(P400I),
				.a1(P401I),
				.a2(P402I),
				.a3(P410I),
				.a4(P411I),
				.a5(P412I),
				.a6(P420I),
				.a7(P421I),
				.a8(P422I),
				.b0(W4000I),
				.b1(W4001I),
				.b2(W4002I),
				.b3(W4010I),
				.b4(W4011I),
				.b5(W4012I),
				.b6(W4020I),
				.b7(W4021I),
				.b8(W4022I),
				.c(c4I000)
);

ninexnine_unit ninexnine_unit_19(
				.clk(clk),
				.rstn(rstn),
				.a0(P400J),
				.a1(P401J),
				.a2(P402J),
				.a3(P410J),
				.a4(P411J),
				.a5(P412J),
				.a6(P420J),
				.a7(P421J),
				.a8(P422J),
				.b0(W4000J),
				.b1(W4001J),
				.b2(W4002J),
				.b3(W4010J),
				.b4(W4011J),
				.b5(W4012J),
				.b6(W4020J),
				.b7(W4021J),
				.b8(W4022J),
				.c(c4J000)
);

ninexnine_unit ninexnine_unit_20(
				.clk(clk),
				.rstn(rstn),
				.a0(P400K),
				.a1(P401K),
				.a2(P402K),
				.a3(P410K),
				.a4(P411K),
				.a5(P412K),
				.a6(P420K),
				.a7(P421K),
				.a8(P422K),
				.b0(W4000K),
				.b1(W4001K),
				.b2(W4002K),
				.b3(W4010K),
				.b4(W4011K),
				.b5(W4012K),
				.b6(W4020K),
				.b7(W4021K),
				.b8(W4022K),
				.c(c4K000)
);

ninexnine_unit ninexnine_unit_21(
				.clk(clk),
				.rstn(rstn),
				.a0(P400L),
				.a1(P401L),
				.a2(P402L),
				.a3(P410L),
				.a4(P411L),
				.a5(P412L),
				.a6(P420L),
				.a7(P421L),
				.a8(P422L),
				.b0(W4000L),
				.b1(W4001L),
				.b2(W4002L),
				.b3(W4010L),
				.b4(W4011L),
				.b5(W4012L),
				.b6(W4020L),
				.b7(W4021L),
				.b8(W4022L),
				.c(c4L000)
);

ninexnine_unit ninexnine_unit_22(
				.clk(clk),
				.rstn(rstn),
				.a0(P400M),
				.a1(P401M),
				.a2(P402M),
				.a3(P410M),
				.a4(P411M),
				.a5(P412M),
				.a6(P420M),
				.a7(P421M),
				.a8(P422M),
				.b0(W4000M),
				.b1(W4001M),
				.b2(W4002M),
				.b3(W4010M),
				.b4(W4011M),
				.b5(W4012M),
				.b6(W4020M),
				.b7(W4021M),
				.b8(W4022M),
				.c(c4M000)
);

ninexnine_unit ninexnine_unit_23(
				.clk(clk),
				.rstn(rstn),
				.a0(P400N),
				.a1(P401N),
				.a2(P402N),
				.a3(P410N),
				.a4(P411N),
				.a5(P412N),
				.a6(P420N),
				.a7(P421N),
				.a8(P422N),
				.b0(W4000N),
				.b1(W4001N),
				.b2(W4002N),
				.b3(W4010N),
				.b4(W4011N),
				.b5(W4012N),
				.b6(W4020N),
				.b7(W4021N),
				.b8(W4022N),
				.c(c4N000)
);

ninexnine_unit ninexnine_unit_24(
				.clk(clk),
				.rstn(rstn),
				.a0(P400O),
				.a1(P401O),
				.a2(P402O),
				.a3(P410O),
				.a4(P411O),
				.a5(P412O),
				.a6(P420O),
				.a7(P421O),
				.a8(P422O),
				.b0(W4000O),
				.b1(W4001O),
				.b2(W4002O),
				.b3(W4010O),
				.b4(W4011O),
				.b5(W4012O),
				.b6(W4020O),
				.b7(W4021O),
				.b8(W4022O),
				.c(c4O000)
);

ninexnine_unit ninexnine_unit_25(
				.clk(clk),
				.rstn(rstn),
				.a0(P400P),
				.a1(P401P),
				.a2(P402P),
				.a3(P410P),
				.a4(P411P),
				.a5(P412P),
				.a6(P420P),
				.a7(P421P),
				.a8(P422P),
				.b0(W4000P),
				.b1(W4001P),
				.b2(W4002P),
				.b3(W4010P),
				.b4(W4011P),
				.b5(W4012P),
				.b6(W4020P),
				.b7(W4021P),
				.b8(W4022P),
				.c(c4P000)
);

ninexnine_unit ninexnine_unit_26(
				.clk(clk),
				.rstn(rstn),
				.a0(P400Q),
				.a1(P401Q),
				.a2(P402Q),
				.a3(P410Q),
				.a4(P411Q),
				.a5(P412Q),
				.a6(P420Q),
				.a7(P421Q),
				.a8(P422Q),
				.b0(W4000Q),
				.b1(W4001Q),
				.b2(W4002Q),
				.b3(W4010Q),
				.b4(W4011Q),
				.b5(W4012Q),
				.b6(W4020Q),
				.b7(W4021Q),
				.b8(W4022Q),
				.c(c4Q000)
);

ninexnine_unit ninexnine_unit_27(
				.clk(clk),
				.rstn(rstn),
				.a0(P400R),
				.a1(P401R),
				.a2(P402R),
				.a3(P410R),
				.a4(P411R),
				.a5(P412R),
				.a6(P420R),
				.a7(P421R),
				.a8(P422R),
				.b0(W4000R),
				.b1(W4001R),
				.b2(W4002R),
				.b3(W4010R),
				.b4(W4011R),
				.b5(W4012R),
				.b6(W4020R),
				.b7(W4021R),
				.b8(W4022R),
				.c(c4R000)
);

ninexnine_unit ninexnine_unit_28(
				.clk(clk),
				.rstn(rstn),
				.a0(P400S),
				.a1(P401S),
				.a2(P402S),
				.a3(P410S),
				.a4(P411S),
				.a5(P412S),
				.a6(P420S),
				.a7(P421S),
				.a8(P422S),
				.b0(W4000S),
				.b1(W4001S),
				.b2(W4002S),
				.b3(W4010S),
				.b4(W4011S),
				.b5(W4012S),
				.b6(W4020S),
				.b7(W4021S),
				.b8(W4022S),
				.c(c4S000)
);

ninexnine_unit ninexnine_unit_29(
				.clk(clk),
				.rstn(rstn),
				.a0(P400T),
				.a1(P401T),
				.a2(P402T),
				.a3(P410T),
				.a4(P411T),
				.a5(P412T),
				.a6(P420T),
				.a7(P421T),
				.a8(P422T),
				.b0(W4000T),
				.b1(W4001T),
				.b2(W4002T),
				.b3(W4010T),
				.b4(W4011T),
				.b5(W4012T),
				.b6(W4020T),
				.b7(W4021T),
				.b8(W4022T),
				.c(c4T000)
);

ninexnine_unit ninexnine_unit_30(
				.clk(clk),
				.rstn(rstn),
				.a0(P400U),
				.a1(P401U),
				.a2(P402U),
				.a3(P410U),
				.a4(P411U),
				.a5(P412U),
				.a6(P420U),
				.a7(P421U),
				.a8(P422U),
				.b0(W4000U),
				.b1(W4001U),
				.b2(W4002U),
				.b3(W4010U),
				.b4(W4011U),
				.b5(W4012U),
				.b6(W4020U),
				.b7(W4021U),
				.b8(W4022U),
				.c(c4U000)
);

ninexnine_unit ninexnine_unit_31(
				.clk(clk),
				.rstn(rstn),
				.a0(P400V),
				.a1(P401V),
				.a2(P402V),
				.a3(P410V),
				.a4(P411V),
				.a5(P412V),
				.a6(P420V),
				.a7(P421V),
				.a8(P422V),
				.b0(W4000V),
				.b1(W4001V),
				.b2(W4002V),
				.b3(W4010V),
				.b4(W4011V),
				.b5(W4012V),
				.b6(W4020V),
				.b7(W4021V),
				.b8(W4022V),
				.c(c4V000)
);

assign C4000=c40000+c41000+c42000+c43000+c44000+c45000+c46000+c47000+c48000+c49000+c4A000+c4B000+c4C000+c4D000+c4E000+c4F000+c4G000+c4H000+c4I000+c4J000+c4K000+c4L000+c4M000+c4N000+c4O000+c4P000+c4Q000+c4R000+c4S000+c4T000+c4U000+c4V000;
assign A4000=(C4000>=0)?1:0;

assign P5000=A4000;

ninexnine_unit ninexnine_unit_32(
				.clk(clk),
				.rstn(rstn),
				.a0(P4000),
				.a1(P4010),
				.a2(P4020),
				.a3(P4100),
				.a4(P4110),
				.a5(P4120),
				.a6(P4200),
				.a7(P4210),
				.a8(P4220),
				.b0(W41000),
				.b1(W41010),
				.b2(W41020),
				.b3(W41100),
				.b4(W41110),
				.b5(W41120),
				.b6(W41200),
				.b7(W41210),
				.b8(W41220),
				.c(c40001)
);

ninexnine_unit ninexnine_unit_33(
				.clk(clk),
				.rstn(rstn),
				.a0(P4001),
				.a1(P4011),
				.a2(P4021),
				.a3(P4101),
				.a4(P4111),
				.a5(P4121),
				.a6(P4201),
				.a7(P4211),
				.a8(P4221),
				.b0(W41001),
				.b1(W41011),
				.b2(W41021),
				.b3(W41101),
				.b4(W41111),
				.b5(W41121),
				.b6(W41201),
				.b7(W41211),
				.b8(W41221),
				.c(c41001)
);

ninexnine_unit ninexnine_unit_34(
				.clk(clk),
				.rstn(rstn),
				.a0(P4002),
				.a1(P4012),
				.a2(P4022),
				.a3(P4102),
				.a4(P4112),
				.a5(P4122),
				.a6(P4202),
				.a7(P4212),
				.a8(P4222),
				.b0(W41002),
				.b1(W41012),
				.b2(W41022),
				.b3(W41102),
				.b4(W41112),
				.b5(W41122),
				.b6(W41202),
				.b7(W41212),
				.b8(W41222),
				.c(c42001)
);

ninexnine_unit ninexnine_unit_35(
				.clk(clk),
				.rstn(rstn),
				.a0(P4003),
				.a1(P4013),
				.a2(P4023),
				.a3(P4103),
				.a4(P4113),
				.a5(P4123),
				.a6(P4203),
				.a7(P4213),
				.a8(P4223),
				.b0(W41003),
				.b1(W41013),
				.b2(W41023),
				.b3(W41103),
				.b4(W41113),
				.b5(W41123),
				.b6(W41203),
				.b7(W41213),
				.b8(W41223),
				.c(c43001)
);

ninexnine_unit ninexnine_unit_36(
				.clk(clk),
				.rstn(rstn),
				.a0(P4004),
				.a1(P4014),
				.a2(P4024),
				.a3(P4104),
				.a4(P4114),
				.a5(P4124),
				.a6(P4204),
				.a7(P4214),
				.a8(P4224),
				.b0(W41004),
				.b1(W41014),
				.b2(W41024),
				.b3(W41104),
				.b4(W41114),
				.b5(W41124),
				.b6(W41204),
				.b7(W41214),
				.b8(W41224),
				.c(c44001)
);

ninexnine_unit ninexnine_unit_37(
				.clk(clk),
				.rstn(rstn),
				.a0(P4005),
				.a1(P4015),
				.a2(P4025),
				.a3(P4105),
				.a4(P4115),
				.a5(P4125),
				.a6(P4205),
				.a7(P4215),
				.a8(P4225),
				.b0(W41005),
				.b1(W41015),
				.b2(W41025),
				.b3(W41105),
				.b4(W41115),
				.b5(W41125),
				.b6(W41205),
				.b7(W41215),
				.b8(W41225),
				.c(c45001)
);

ninexnine_unit ninexnine_unit_38(
				.clk(clk),
				.rstn(rstn),
				.a0(P4006),
				.a1(P4016),
				.a2(P4026),
				.a3(P4106),
				.a4(P4116),
				.a5(P4126),
				.a6(P4206),
				.a7(P4216),
				.a8(P4226),
				.b0(W41006),
				.b1(W41016),
				.b2(W41026),
				.b3(W41106),
				.b4(W41116),
				.b5(W41126),
				.b6(W41206),
				.b7(W41216),
				.b8(W41226),
				.c(c46001)
);

ninexnine_unit ninexnine_unit_39(
				.clk(clk),
				.rstn(rstn),
				.a0(P4007),
				.a1(P4017),
				.a2(P4027),
				.a3(P4107),
				.a4(P4117),
				.a5(P4127),
				.a6(P4207),
				.a7(P4217),
				.a8(P4227),
				.b0(W41007),
				.b1(W41017),
				.b2(W41027),
				.b3(W41107),
				.b4(W41117),
				.b5(W41127),
				.b6(W41207),
				.b7(W41217),
				.b8(W41227),
				.c(c47001)
);

ninexnine_unit ninexnine_unit_40(
				.clk(clk),
				.rstn(rstn),
				.a0(P4008),
				.a1(P4018),
				.a2(P4028),
				.a3(P4108),
				.a4(P4118),
				.a5(P4128),
				.a6(P4208),
				.a7(P4218),
				.a8(P4228),
				.b0(W41008),
				.b1(W41018),
				.b2(W41028),
				.b3(W41108),
				.b4(W41118),
				.b5(W41128),
				.b6(W41208),
				.b7(W41218),
				.b8(W41228),
				.c(c48001)
);

ninexnine_unit ninexnine_unit_41(
				.clk(clk),
				.rstn(rstn),
				.a0(P4009),
				.a1(P4019),
				.a2(P4029),
				.a3(P4109),
				.a4(P4119),
				.a5(P4129),
				.a6(P4209),
				.a7(P4219),
				.a8(P4229),
				.b0(W41009),
				.b1(W41019),
				.b2(W41029),
				.b3(W41109),
				.b4(W41119),
				.b5(W41129),
				.b6(W41209),
				.b7(W41219),
				.b8(W41229),
				.c(c49001)
);

ninexnine_unit ninexnine_unit_42(
				.clk(clk),
				.rstn(rstn),
				.a0(P400A),
				.a1(P401A),
				.a2(P402A),
				.a3(P410A),
				.a4(P411A),
				.a5(P412A),
				.a6(P420A),
				.a7(P421A),
				.a8(P422A),
				.b0(W4100A),
				.b1(W4101A),
				.b2(W4102A),
				.b3(W4110A),
				.b4(W4111A),
				.b5(W4112A),
				.b6(W4120A),
				.b7(W4121A),
				.b8(W4122A),
				.c(c4A001)
);

ninexnine_unit ninexnine_unit_43(
				.clk(clk),
				.rstn(rstn),
				.a0(P400B),
				.a1(P401B),
				.a2(P402B),
				.a3(P410B),
				.a4(P411B),
				.a5(P412B),
				.a6(P420B),
				.a7(P421B),
				.a8(P422B),
				.b0(W4100B),
				.b1(W4101B),
				.b2(W4102B),
				.b3(W4110B),
				.b4(W4111B),
				.b5(W4112B),
				.b6(W4120B),
				.b7(W4121B),
				.b8(W4122B),
				.c(c4B001)
);

ninexnine_unit ninexnine_unit_44(
				.clk(clk),
				.rstn(rstn),
				.a0(P400C),
				.a1(P401C),
				.a2(P402C),
				.a3(P410C),
				.a4(P411C),
				.a5(P412C),
				.a6(P420C),
				.a7(P421C),
				.a8(P422C),
				.b0(W4100C),
				.b1(W4101C),
				.b2(W4102C),
				.b3(W4110C),
				.b4(W4111C),
				.b5(W4112C),
				.b6(W4120C),
				.b7(W4121C),
				.b8(W4122C),
				.c(c4C001)
);

ninexnine_unit ninexnine_unit_45(
				.clk(clk),
				.rstn(rstn),
				.a0(P400D),
				.a1(P401D),
				.a2(P402D),
				.a3(P410D),
				.a4(P411D),
				.a5(P412D),
				.a6(P420D),
				.a7(P421D),
				.a8(P422D),
				.b0(W4100D),
				.b1(W4101D),
				.b2(W4102D),
				.b3(W4110D),
				.b4(W4111D),
				.b5(W4112D),
				.b6(W4120D),
				.b7(W4121D),
				.b8(W4122D),
				.c(c4D001)
);

ninexnine_unit ninexnine_unit_46(
				.clk(clk),
				.rstn(rstn),
				.a0(P400E),
				.a1(P401E),
				.a2(P402E),
				.a3(P410E),
				.a4(P411E),
				.a5(P412E),
				.a6(P420E),
				.a7(P421E),
				.a8(P422E),
				.b0(W4100E),
				.b1(W4101E),
				.b2(W4102E),
				.b3(W4110E),
				.b4(W4111E),
				.b5(W4112E),
				.b6(W4120E),
				.b7(W4121E),
				.b8(W4122E),
				.c(c4E001)
);

ninexnine_unit ninexnine_unit_47(
				.clk(clk),
				.rstn(rstn),
				.a0(P400F),
				.a1(P401F),
				.a2(P402F),
				.a3(P410F),
				.a4(P411F),
				.a5(P412F),
				.a6(P420F),
				.a7(P421F),
				.a8(P422F),
				.b0(W4100F),
				.b1(W4101F),
				.b2(W4102F),
				.b3(W4110F),
				.b4(W4111F),
				.b5(W4112F),
				.b6(W4120F),
				.b7(W4121F),
				.b8(W4122F),
				.c(c4F001)
);

ninexnine_unit ninexnine_unit_48(
				.clk(clk),
				.rstn(rstn),
				.a0(P400G),
				.a1(P401G),
				.a2(P402G),
				.a3(P410G),
				.a4(P411G),
				.a5(P412G),
				.a6(P420G),
				.a7(P421G),
				.a8(P422G),
				.b0(W4100G),
				.b1(W4101G),
				.b2(W4102G),
				.b3(W4110G),
				.b4(W4111G),
				.b5(W4112G),
				.b6(W4120G),
				.b7(W4121G),
				.b8(W4122G),
				.c(c4G001)
);

ninexnine_unit ninexnine_unit_49(
				.clk(clk),
				.rstn(rstn),
				.a0(P400H),
				.a1(P401H),
				.a2(P402H),
				.a3(P410H),
				.a4(P411H),
				.a5(P412H),
				.a6(P420H),
				.a7(P421H),
				.a8(P422H),
				.b0(W4100H),
				.b1(W4101H),
				.b2(W4102H),
				.b3(W4110H),
				.b4(W4111H),
				.b5(W4112H),
				.b6(W4120H),
				.b7(W4121H),
				.b8(W4122H),
				.c(c4H001)
);

ninexnine_unit ninexnine_unit_50(
				.clk(clk),
				.rstn(rstn),
				.a0(P400I),
				.a1(P401I),
				.a2(P402I),
				.a3(P410I),
				.a4(P411I),
				.a5(P412I),
				.a6(P420I),
				.a7(P421I),
				.a8(P422I),
				.b0(W4100I),
				.b1(W4101I),
				.b2(W4102I),
				.b3(W4110I),
				.b4(W4111I),
				.b5(W4112I),
				.b6(W4120I),
				.b7(W4121I),
				.b8(W4122I),
				.c(c4I001)
);

ninexnine_unit ninexnine_unit_51(
				.clk(clk),
				.rstn(rstn),
				.a0(P400J),
				.a1(P401J),
				.a2(P402J),
				.a3(P410J),
				.a4(P411J),
				.a5(P412J),
				.a6(P420J),
				.a7(P421J),
				.a8(P422J),
				.b0(W4100J),
				.b1(W4101J),
				.b2(W4102J),
				.b3(W4110J),
				.b4(W4111J),
				.b5(W4112J),
				.b6(W4120J),
				.b7(W4121J),
				.b8(W4122J),
				.c(c4J001)
);

ninexnine_unit ninexnine_unit_52(
				.clk(clk),
				.rstn(rstn),
				.a0(P400K),
				.a1(P401K),
				.a2(P402K),
				.a3(P410K),
				.a4(P411K),
				.a5(P412K),
				.a6(P420K),
				.a7(P421K),
				.a8(P422K),
				.b0(W4100K),
				.b1(W4101K),
				.b2(W4102K),
				.b3(W4110K),
				.b4(W4111K),
				.b5(W4112K),
				.b6(W4120K),
				.b7(W4121K),
				.b8(W4122K),
				.c(c4K001)
);

ninexnine_unit ninexnine_unit_53(
				.clk(clk),
				.rstn(rstn),
				.a0(P400L),
				.a1(P401L),
				.a2(P402L),
				.a3(P410L),
				.a4(P411L),
				.a5(P412L),
				.a6(P420L),
				.a7(P421L),
				.a8(P422L),
				.b0(W4100L),
				.b1(W4101L),
				.b2(W4102L),
				.b3(W4110L),
				.b4(W4111L),
				.b5(W4112L),
				.b6(W4120L),
				.b7(W4121L),
				.b8(W4122L),
				.c(c4L001)
);

ninexnine_unit ninexnine_unit_54(
				.clk(clk),
				.rstn(rstn),
				.a0(P400M),
				.a1(P401M),
				.a2(P402M),
				.a3(P410M),
				.a4(P411M),
				.a5(P412M),
				.a6(P420M),
				.a7(P421M),
				.a8(P422M),
				.b0(W4100M),
				.b1(W4101M),
				.b2(W4102M),
				.b3(W4110M),
				.b4(W4111M),
				.b5(W4112M),
				.b6(W4120M),
				.b7(W4121M),
				.b8(W4122M),
				.c(c4M001)
);

ninexnine_unit ninexnine_unit_55(
				.clk(clk),
				.rstn(rstn),
				.a0(P400N),
				.a1(P401N),
				.a2(P402N),
				.a3(P410N),
				.a4(P411N),
				.a5(P412N),
				.a6(P420N),
				.a7(P421N),
				.a8(P422N),
				.b0(W4100N),
				.b1(W4101N),
				.b2(W4102N),
				.b3(W4110N),
				.b4(W4111N),
				.b5(W4112N),
				.b6(W4120N),
				.b7(W4121N),
				.b8(W4122N),
				.c(c4N001)
);

ninexnine_unit ninexnine_unit_56(
				.clk(clk),
				.rstn(rstn),
				.a0(P400O),
				.a1(P401O),
				.a2(P402O),
				.a3(P410O),
				.a4(P411O),
				.a5(P412O),
				.a6(P420O),
				.a7(P421O),
				.a8(P422O),
				.b0(W4100O),
				.b1(W4101O),
				.b2(W4102O),
				.b3(W4110O),
				.b4(W4111O),
				.b5(W4112O),
				.b6(W4120O),
				.b7(W4121O),
				.b8(W4122O),
				.c(c4O001)
);

ninexnine_unit ninexnine_unit_57(
				.clk(clk),
				.rstn(rstn),
				.a0(P400P),
				.a1(P401P),
				.a2(P402P),
				.a3(P410P),
				.a4(P411P),
				.a5(P412P),
				.a6(P420P),
				.a7(P421P),
				.a8(P422P),
				.b0(W4100P),
				.b1(W4101P),
				.b2(W4102P),
				.b3(W4110P),
				.b4(W4111P),
				.b5(W4112P),
				.b6(W4120P),
				.b7(W4121P),
				.b8(W4122P),
				.c(c4P001)
);

ninexnine_unit ninexnine_unit_58(
				.clk(clk),
				.rstn(rstn),
				.a0(P400Q),
				.a1(P401Q),
				.a2(P402Q),
				.a3(P410Q),
				.a4(P411Q),
				.a5(P412Q),
				.a6(P420Q),
				.a7(P421Q),
				.a8(P422Q),
				.b0(W4100Q),
				.b1(W4101Q),
				.b2(W4102Q),
				.b3(W4110Q),
				.b4(W4111Q),
				.b5(W4112Q),
				.b6(W4120Q),
				.b7(W4121Q),
				.b8(W4122Q),
				.c(c4Q001)
);

ninexnine_unit ninexnine_unit_59(
				.clk(clk),
				.rstn(rstn),
				.a0(P400R),
				.a1(P401R),
				.a2(P402R),
				.a3(P410R),
				.a4(P411R),
				.a5(P412R),
				.a6(P420R),
				.a7(P421R),
				.a8(P422R),
				.b0(W4100R),
				.b1(W4101R),
				.b2(W4102R),
				.b3(W4110R),
				.b4(W4111R),
				.b5(W4112R),
				.b6(W4120R),
				.b7(W4121R),
				.b8(W4122R),
				.c(c4R001)
);

ninexnine_unit ninexnine_unit_60(
				.clk(clk),
				.rstn(rstn),
				.a0(P400S),
				.a1(P401S),
				.a2(P402S),
				.a3(P410S),
				.a4(P411S),
				.a5(P412S),
				.a6(P420S),
				.a7(P421S),
				.a8(P422S),
				.b0(W4100S),
				.b1(W4101S),
				.b2(W4102S),
				.b3(W4110S),
				.b4(W4111S),
				.b5(W4112S),
				.b6(W4120S),
				.b7(W4121S),
				.b8(W4122S),
				.c(c4S001)
);

ninexnine_unit ninexnine_unit_61(
				.clk(clk),
				.rstn(rstn),
				.a0(P400T),
				.a1(P401T),
				.a2(P402T),
				.a3(P410T),
				.a4(P411T),
				.a5(P412T),
				.a6(P420T),
				.a7(P421T),
				.a8(P422T),
				.b0(W4100T),
				.b1(W4101T),
				.b2(W4102T),
				.b3(W4110T),
				.b4(W4111T),
				.b5(W4112T),
				.b6(W4120T),
				.b7(W4121T),
				.b8(W4122T),
				.c(c4T001)
);

ninexnine_unit ninexnine_unit_62(
				.clk(clk),
				.rstn(rstn),
				.a0(P400U),
				.a1(P401U),
				.a2(P402U),
				.a3(P410U),
				.a4(P411U),
				.a5(P412U),
				.a6(P420U),
				.a7(P421U),
				.a8(P422U),
				.b0(W4100U),
				.b1(W4101U),
				.b2(W4102U),
				.b3(W4110U),
				.b4(W4111U),
				.b5(W4112U),
				.b6(W4120U),
				.b7(W4121U),
				.b8(W4122U),
				.c(c4U001)
);

ninexnine_unit ninexnine_unit_63(
				.clk(clk),
				.rstn(rstn),
				.a0(P400V),
				.a1(P401V),
				.a2(P402V),
				.a3(P410V),
				.a4(P411V),
				.a5(P412V),
				.a6(P420V),
				.a7(P421V),
				.a8(P422V),
				.b0(W4100V),
				.b1(W4101V),
				.b2(W4102V),
				.b3(W4110V),
				.b4(W4111V),
				.b5(W4112V),
				.b6(W4120V),
				.b7(W4121V),
				.b8(W4122V),
				.c(c4V001)
);

assign C4001=c40001+c41001+c42001+c43001+c44001+c45001+c46001+c47001+c48001+c49001+c4A001+c4B001+c4C001+c4D001+c4E001+c4F001+c4G001+c4H001+c4I001+c4J001+c4K001+c4L001+c4M001+c4N001+c4O001+c4P001+c4Q001+c4R001+c4S001+c4T001+c4U001+c4V001;
assign A4001=(C4001>=0)?1:0;

assign P5001=A4001;

endmodule