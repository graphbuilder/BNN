module test_layer_all(
clk, 
rstn
);
input clk;
input rstn;

wire P0000;
wire P0010;
wire P0020;
wire P0030;
wire P0040;
wire P0050;
wire P0060;
wire P0100;
wire P0110;
wire P0120;
wire P0130;
wire P0140;
wire P0150;
wire P0160;
wire P0200;
wire P0210;
wire P0220;
wire P0230;
wire P0240;
wire P0250;
wire P0260;
wire P0300;
wire P0310;
wire P0320;
wire P0330;
wire P0340;
wire P0350;
wire P0360;
wire P0400;
wire P0410;
wire P0420;
wire P0430;
wire P0440;
wire P0450;
wire P0460;
wire P0500;
wire P0510;
wire P0520;
wire P0530;
wire P0540;
wire P0550;
wire P0560;
wire P0600;
wire P0610;
wire P0620;
wire P0630;
wire P0640;
wire P0650;
wire P0660;
wire P0001;
wire P0011;
wire P0021;
wire P0031;
wire P0041;
wire P0051;
wire P0061;
wire P0101;
wire P0111;
wire P0121;
wire P0131;
wire P0141;
wire P0151;
wire P0161;
wire P0201;
wire P0211;
wire P0221;
wire P0231;
wire P0241;
wire P0251;
wire P0261;
wire P0301;
wire P0311;
wire P0321;
wire P0331;
wire P0341;
wire P0351;
wire P0361;
wire P0401;
wire P0411;
wire P0421;
wire P0431;
wire P0441;
wire P0451;
wire P0461;
wire P0501;
wire P0511;
wire P0521;
wire P0531;
wire P0541;
wire P0551;
wire P0561;
wire P0601;
wire P0611;
wire P0621;
wire P0631;
wire P0641;
wire P0651;
wire P0661;
wire P0002;
wire P0012;
wire P0022;
wire P0032;
wire P0042;
wire P0052;
wire P0062;
wire P0102;
wire P0112;
wire P0122;
wire P0132;
wire P0142;
wire P0152;
wire P0162;
wire P0202;
wire P0212;
wire P0222;
wire P0232;
wire P0242;
wire P0252;
wire P0262;
wire P0302;
wire P0312;
wire P0322;
wire P0332;
wire P0342;
wire P0352;
wire P0362;
wire P0402;
wire P0412;
wire P0422;
wire P0432;
wire P0442;
wire P0452;
wire P0462;
wire P0502;
wire P0512;
wire P0522;
wire P0532;
wire P0542;
wire P0552;
wire P0562;
wire P0602;
wire P0612;
wire P0622;
wire P0632;
wire P0642;
wire P0652;
wire P0662;
wire P1000;
wire P1010;
wire P1020;
wire P1030;
wire P1040;
wire P1100;
wire P1110;
wire P1120;
wire P1130;
wire P1140;
wire P1200;
wire P1210;
wire P1220;
wire P1230;
wire P1240;
wire P1300;
wire P1310;
wire P1320;
wire P1330;
wire P1340;
wire P1400;
wire P1410;
wire P1420;
wire P1430;
wire P1440;
wire P1001;
wire P1011;
wire P1021;
wire P1031;
wire P1041;
wire P1101;
wire P1111;
wire P1121;
wire P1131;
wire P1141;
wire P1201;
wire P1211;
wire P1221;
wire P1231;
wire P1241;
wire P1301;
wire P1311;
wire P1321;
wire P1331;
wire P1341;
wire P1401;
wire P1411;
wire P1421;
wire P1431;
wire P1441;
wire P1002;
wire P1012;
wire P1022;
wire P1032;
wire P1042;
wire P1102;
wire P1112;
wire P1122;
wire P1132;
wire P1142;
wire P1202;
wire P1212;
wire P1222;
wire P1232;
wire P1242;
wire P1302;
wire P1312;
wire P1322;
wire P1332;
wire P1342;
wire P1402;
wire P1412;
wire P1422;
wire P1432;
wire P1442;
wire P1003;
wire P1013;
wire P1023;
wire P1033;
wire P1043;
wire P1103;
wire P1113;
wire P1123;
wire P1133;
wire P1143;
wire P1203;
wire P1213;
wire P1223;
wire P1233;
wire P1243;
wire P1303;
wire P1313;
wire P1323;
wire P1333;
wire P1343;
wire P1403;
wire P1413;
wire P1423;
wire P1433;
wire P1443;
wire P1004;
wire P1014;
wire P1024;
wire P1034;
wire P1044;
wire P1104;
wire P1114;
wire P1124;
wire P1134;
wire P1144;
wire P1204;
wire P1214;
wire P1224;
wire P1234;
wire P1244;
wire P1304;
wire P1314;
wire P1324;
wire P1334;
wire P1344;
wire P1404;
wire P1414;
wire P1424;
wire P1434;
wire P1444;
wire P1005;
wire P1015;
wire P1025;
wire P1035;
wire P1045;
wire P1105;
wire P1115;
wire P1125;
wire P1135;
wire P1145;
wire P1205;
wire P1215;
wire P1225;
wire P1235;
wire P1245;
wire P1305;
wire P1315;
wire P1325;
wire P1335;
wire P1345;
wire P1405;
wire P1415;
wire P1425;
wire P1435;
wire P1445;
wire P1006;
wire P1016;
wire P1026;
wire P1036;
wire P1046;
wire P1106;
wire P1116;
wire P1126;
wire P1136;
wire P1146;
wire P1206;
wire P1216;
wire P1226;
wire P1236;
wire P1246;
wire P1306;
wire P1316;
wire P1326;
wire P1336;
wire P1346;
wire P1406;
wire P1416;
wire P1426;
wire P1436;
wire P1446;
wire P1007;
wire P1017;
wire P1027;
wire P1037;
wire P1047;
wire P1107;
wire P1117;
wire P1127;
wire P1137;
wire P1147;
wire P1207;
wire P1217;
wire P1227;
wire P1237;
wire P1247;
wire P1307;
wire P1317;
wire P1327;
wire P1337;
wire P1347;
wire P1407;
wire P1417;
wire P1427;
wire P1437;
wire P1447;
wire P1008;
wire P1018;
wire P1028;
wire P1038;
wire P1048;
wire P1108;
wire P1118;
wire P1128;
wire P1138;
wire P1148;
wire P1208;
wire P1218;
wire P1228;
wire P1238;
wire P1248;
wire P1308;
wire P1318;
wire P1328;
wire P1338;
wire P1348;
wire P1408;
wire P1418;
wire P1428;
wire P1438;
wire P1448;
wire P1009;
wire P1019;
wire P1029;
wire P1039;
wire P1049;
wire P1109;
wire P1119;
wire P1129;
wire P1139;
wire P1149;
wire P1209;
wire P1219;
wire P1229;
wire P1239;
wire P1249;
wire P1309;
wire P1319;
wire P1329;
wire P1339;
wire P1349;
wire P1409;
wire P1419;
wire P1429;
wire P1439;
wire P1449;
wire P100A;
wire P101A;
wire P102A;
wire P103A;
wire P104A;
wire P110A;
wire P111A;
wire P112A;
wire P113A;
wire P114A;
wire P120A;
wire P121A;
wire P122A;
wire P123A;
wire P124A;
wire P130A;
wire P131A;
wire P132A;
wire P133A;
wire P134A;
wire P140A;
wire P141A;
wire P142A;
wire P143A;
wire P144A;
wire P100B;
wire P101B;
wire P102B;
wire P103B;
wire P104B;
wire P110B;
wire P111B;
wire P112B;
wire P113B;
wire P114B;
wire P120B;
wire P121B;
wire P122B;
wire P123B;
wire P124B;
wire P130B;
wire P131B;
wire P132B;
wire P133B;
wire P134B;
wire P140B;
wire P141B;
wire P142B;
wire P143B;
wire P144B;
wire P100C;
wire P101C;
wire P102C;
wire P103C;
wire P104C;
wire P110C;
wire P111C;
wire P112C;
wire P113C;
wire P114C;
wire P120C;
wire P121C;
wire P122C;
wire P123C;
wire P124C;
wire P130C;
wire P131C;
wire P132C;
wire P133C;
wire P134C;
wire P140C;
wire P141C;
wire P142C;
wire P143C;
wire P144C;
wire P100D;
wire P101D;
wire P102D;
wire P103D;
wire P104D;
wire P110D;
wire P111D;
wire P112D;
wire P113D;
wire P114D;
wire P120D;
wire P121D;
wire P122D;
wire P123D;
wire P124D;
wire P130D;
wire P131D;
wire P132D;
wire P133D;
wire P134D;
wire P140D;
wire P141D;
wire P142D;
wire P143D;
wire P144D;
wire P100E;
wire P101E;
wire P102E;
wire P103E;
wire P104E;
wire P110E;
wire P111E;
wire P112E;
wire P113E;
wire P114E;
wire P120E;
wire P121E;
wire P122E;
wire P123E;
wire P124E;
wire P130E;
wire P131E;
wire P132E;
wire P133E;
wire P134E;
wire P140E;
wire P141E;
wire P142E;
wire P143E;
wire P144E;
wire P100F;
wire P101F;
wire P102F;
wire P103F;
wire P104F;
wire P110F;
wire P111F;
wire P112F;
wire P113F;
wire P114F;
wire P120F;
wire P121F;
wire P122F;
wire P123F;
wire P124F;
wire P130F;
wire P131F;
wire P132F;
wire P133F;
wire P134F;
wire P140F;
wire P141F;
wire P142F;
wire P143F;
wire P144F;
wire W00000,W00010,W00020,W00100,W00110,W00120,W00200,W00210,W00220;
wire W00001,W00011,W00021,W00101,W00111,W00121,W00201,W00211,W00221;
wire W00002,W00012,W00022,W00102,W00112,W00122,W00202,W00212,W00222;
wire W01000,W01010,W01020,W01100,W01110,W01120,W01200,W01210,W01220;
wire W01001,W01011,W01021,W01101,W01111,W01121,W01201,W01211,W01221;
wire W01002,W01012,W01022,W01102,W01112,W01122,W01202,W01212,W01222;
wire W02000,W02010,W02020,W02100,W02110,W02120,W02200,W02210,W02220;
wire W02001,W02011,W02021,W02101,W02111,W02121,W02201,W02211,W02221;
wire W02002,W02012,W02022,W02102,W02112,W02122,W02202,W02212,W02222;
wire W03000,W03010,W03020,W03100,W03110,W03120,W03200,W03210,W03220;
wire W03001,W03011,W03021,W03101,W03111,W03121,W03201,W03211,W03221;
wire W03002,W03012,W03022,W03102,W03112,W03122,W03202,W03212,W03222;
wire W04000,W04010,W04020,W04100,W04110,W04120,W04200,W04210,W04220;
wire W04001,W04011,W04021,W04101,W04111,W04121,W04201,W04211,W04221;
wire W04002,W04012,W04022,W04102,W04112,W04122,W04202,W04212,W04222;
wire W05000,W05010,W05020,W05100,W05110,W05120,W05200,W05210,W05220;
wire W05001,W05011,W05021,W05101,W05111,W05121,W05201,W05211,W05221;
wire W05002,W05012,W05022,W05102,W05112,W05122,W05202,W05212,W05222;
wire W06000,W06010,W06020,W06100,W06110,W06120,W06200,W06210,W06220;
wire W06001,W06011,W06021,W06101,W06111,W06121,W06201,W06211,W06221;
wire W06002,W06012,W06022,W06102,W06112,W06122,W06202,W06212,W06222;
wire W07000,W07010,W07020,W07100,W07110,W07120,W07200,W07210,W07220;
wire W07001,W07011,W07021,W07101,W07111,W07121,W07201,W07211,W07221;
wire W07002,W07012,W07022,W07102,W07112,W07122,W07202,W07212,W07222;
wire W08000,W08010,W08020,W08100,W08110,W08120,W08200,W08210,W08220;
wire W08001,W08011,W08021,W08101,W08111,W08121,W08201,W08211,W08221;
wire W08002,W08012,W08022,W08102,W08112,W08122,W08202,W08212,W08222;
wire W09000,W09010,W09020,W09100,W09110,W09120,W09200,W09210,W09220;
wire W09001,W09011,W09021,W09101,W09111,W09121,W09201,W09211,W09221;
wire W09002,W09012,W09022,W09102,W09112,W09122,W09202,W09212,W09222;
wire W0A000,W0A010,W0A020,W0A100,W0A110,W0A120,W0A200,W0A210,W0A220;
wire W0A001,W0A011,W0A021,W0A101,W0A111,W0A121,W0A201,W0A211,W0A221;
wire W0A002,W0A012,W0A022,W0A102,W0A112,W0A122,W0A202,W0A212,W0A222;
wire W0B000,W0B010,W0B020,W0B100,W0B110,W0B120,W0B200,W0B210,W0B220;
wire W0B001,W0B011,W0B021,W0B101,W0B111,W0B121,W0B201,W0B211,W0B221;
wire W0B002,W0B012,W0B022,W0B102,W0B112,W0B122,W0B202,W0B212,W0B222;
wire W0C000,W0C010,W0C020,W0C100,W0C110,W0C120,W0C200,W0C210,W0C220;
wire W0C001,W0C011,W0C021,W0C101,W0C111,W0C121,W0C201,W0C211,W0C221;
wire W0C002,W0C012,W0C022,W0C102,W0C112,W0C122,W0C202,W0C212,W0C222;
wire W0D000,W0D010,W0D020,W0D100,W0D110,W0D120,W0D200,W0D210,W0D220;
wire W0D001,W0D011,W0D021,W0D101,W0D111,W0D121,W0D201,W0D211,W0D221;
wire W0D002,W0D012,W0D022,W0D102,W0D112,W0D122,W0D202,W0D212,W0D222;
wire W0E000,W0E010,W0E020,W0E100,W0E110,W0E120,W0E200,W0E210,W0E220;
wire W0E001,W0E011,W0E021,W0E101,W0E111,W0E121,W0E201,W0E211,W0E221;
wire W0E002,W0E012,W0E022,W0E102,W0E112,W0E122,W0E202,W0E212,W0E222;
wire W0F000,W0F010,W0F020,W0F100,W0F110,W0F120,W0F200,W0F210,W0F220;
wire W0F001,W0F011,W0F021,W0F101,W0F111,W0F121,W0F201,W0F211,W0F221;
wire W0F002,W0F012,W0F022,W0F102,W0F112,W0F122,W0F202,W0F212,W0F222;
wire signed [4:0] c00000,c01000,c02000;
wire signed [4:0] c00010,c01010,c02010;
wire signed [4:0] c00020,c01020,c02020;
wire signed [4:0] c00030,c01030,c02030;
wire signed [4:0] c00040,c01040,c02040;
wire signed [4:0] c00100,c01100,c02100;
wire signed [4:0] c00110,c01110,c02110;
wire signed [4:0] c00120,c01120,c02120;
wire signed [4:0] c00130,c01130,c02130;
wire signed [4:0] c00140,c01140,c02140;
wire signed [4:0] c00200,c01200,c02200;
wire signed [4:0] c00210,c01210,c02210;
wire signed [4:0] c00220,c01220,c02220;
wire signed [4:0] c00230,c01230,c02230;
wire signed [4:0] c00240,c01240,c02240;
wire signed [4:0] c00300,c01300,c02300;
wire signed [4:0] c00310,c01310,c02310;
wire signed [4:0] c00320,c01320,c02320;
wire signed [4:0] c00330,c01330,c02330;
wire signed [4:0] c00340,c01340,c02340;
wire signed [4:0] c00400,c01400,c02400;
wire signed [4:0] c00410,c01410,c02410;
wire signed [4:0] c00420,c01420,c02420;
wire signed [4:0] c00430,c01430,c02430;
wire signed [4:0] c00440,c01440,c02440;
wire signed [4:0] c00001,c01001,c02001;
wire signed [4:0] c00011,c01011,c02011;
wire signed [4:0] c00021,c01021,c02021;
wire signed [4:0] c00031,c01031,c02031;
wire signed [4:0] c00041,c01041,c02041;
wire signed [4:0] c00101,c01101,c02101;
wire signed [4:0] c00111,c01111,c02111;
wire signed [4:0] c00121,c01121,c02121;
wire signed [4:0] c00131,c01131,c02131;
wire signed [4:0] c00141,c01141,c02141;
wire signed [4:0] c00201,c01201,c02201;
wire signed [4:0] c00211,c01211,c02211;
wire signed [4:0] c00221,c01221,c02221;
wire signed [4:0] c00231,c01231,c02231;
wire signed [4:0] c00241,c01241,c02241;
wire signed [4:0] c00301,c01301,c02301;
wire signed [4:0] c00311,c01311,c02311;
wire signed [4:0] c00321,c01321,c02321;
wire signed [4:0] c00331,c01331,c02331;
wire signed [4:0] c00341,c01341,c02341;
wire signed [4:0] c00401,c01401,c02401;
wire signed [4:0] c00411,c01411,c02411;
wire signed [4:0] c00421,c01421,c02421;
wire signed [4:0] c00431,c01431,c02431;
wire signed [4:0] c00441,c01441,c02441;
wire signed [4:0] c00002,c01002,c02002;
wire signed [4:0] c00012,c01012,c02012;
wire signed [4:0] c00022,c01022,c02022;
wire signed [4:0] c00032,c01032,c02032;
wire signed [4:0] c00042,c01042,c02042;
wire signed [4:0] c00102,c01102,c02102;
wire signed [4:0] c00112,c01112,c02112;
wire signed [4:0] c00122,c01122,c02122;
wire signed [4:0] c00132,c01132,c02132;
wire signed [4:0] c00142,c01142,c02142;
wire signed [4:0] c00202,c01202,c02202;
wire signed [4:0] c00212,c01212,c02212;
wire signed [4:0] c00222,c01222,c02222;
wire signed [4:0] c00232,c01232,c02232;
wire signed [4:0] c00242,c01242,c02242;
wire signed [4:0] c00302,c01302,c02302;
wire signed [4:0] c00312,c01312,c02312;
wire signed [4:0] c00322,c01322,c02322;
wire signed [4:0] c00332,c01332,c02332;
wire signed [4:0] c00342,c01342,c02342;
wire signed [4:0] c00402,c01402,c02402;
wire signed [4:0] c00412,c01412,c02412;
wire signed [4:0] c00422,c01422,c02422;
wire signed [4:0] c00432,c01432,c02432;
wire signed [4:0] c00442,c01442,c02442;
wire signed [4:0] c00003,c01003,c02003;
wire signed [4:0] c00013,c01013,c02013;
wire signed [4:0] c00023,c01023,c02023;
wire signed [4:0] c00033,c01033,c02033;
wire signed [4:0] c00043,c01043,c02043;
wire signed [4:0] c00103,c01103,c02103;
wire signed [4:0] c00113,c01113,c02113;
wire signed [4:0] c00123,c01123,c02123;
wire signed [4:0] c00133,c01133,c02133;
wire signed [4:0] c00143,c01143,c02143;
wire signed [4:0] c00203,c01203,c02203;
wire signed [4:0] c00213,c01213,c02213;
wire signed [4:0] c00223,c01223,c02223;
wire signed [4:0] c00233,c01233,c02233;
wire signed [4:0] c00243,c01243,c02243;
wire signed [4:0] c00303,c01303,c02303;
wire signed [4:0] c00313,c01313,c02313;
wire signed [4:0] c00323,c01323,c02323;
wire signed [4:0] c00333,c01333,c02333;
wire signed [4:0] c00343,c01343,c02343;
wire signed [4:0] c00403,c01403,c02403;
wire signed [4:0] c00413,c01413,c02413;
wire signed [4:0] c00423,c01423,c02423;
wire signed [4:0] c00433,c01433,c02433;
wire signed [4:0] c00443,c01443,c02443;
wire signed [4:0] c00004,c01004,c02004;
wire signed [4:0] c00014,c01014,c02014;
wire signed [4:0] c00024,c01024,c02024;
wire signed [4:0] c00034,c01034,c02034;
wire signed [4:0] c00044,c01044,c02044;
wire signed [4:0] c00104,c01104,c02104;
wire signed [4:0] c00114,c01114,c02114;
wire signed [4:0] c00124,c01124,c02124;
wire signed [4:0] c00134,c01134,c02134;
wire signed [4:0] c00144,c01144,c02144;
wire signed [4:0] c00204,c01204,c02204;
wire signed [4:0] c00214,c01214,c02214;
wire signed [4:0] c00224,c01224,c02224;
wire signed [4:0] c00234,c01234,c02234;
wire signed [4:0] c00244,c01244,c02244;
wire signed [4:0] c00304,c01304,c02304;
wire signed [4:0] c00314,c01314,c02314;
wire signed [4:0] c00324,c01324,c02324;
wire signed [4:0] c00334,c01334,c02334;
wire signed [4:0] c00344,c01344,c02344;
wire signed [4:0] c00404,c01404,c02404;
wire signed [4:0] c00414,c01414,c02414;
wire signed [4:0] c00424,c01424,c02424;
wire signed [4:0] c00434,c01434,c02434;
wire signed [4:0] c00444,c01444,c02444;
wire signed [4:0] c00005,c01005,c02005;
wire signed [4:0] c00015,c01015,c02015;
wire signed [4:0] c00025,c01025,c02025;
wire signed [4:0] c00035,c01035,c02035;
wire signed [4:0] c00045,c01045,c02045;
wire signed [4:0] c00105,c01105,c02105;
wire signed [4:0] c00115,c01115,c02115;
wire signed [4:0] c00125,c01125,c02125;
wire signed [4:0] c00135,c01135,c02135;
wire signed [4:0] c00145,c01145,c02145;
wire signed [4:0] c00205,c01205,c02205;
wire signed [4:0] c00215,c01215,c02215;
wire signed [4:0] c00225,c01225,c02225;
wire signed [4:0] c00235,c01235,c02235;
wire signed [4:0] c00245,c01245,c02245;
wire signed [4:0] c00305,c01305,c02305;
wire signed [4:0] c00315,c01315,c02315;
wire signed [4:0] c00325,c01325,c02325;
wire signed [4:0] c00335,c01335,c02335;
wire signed [4:0] c00345,c01345,c02345;
wire signed [4:0] c00405,c01405,c02405;
wire signed [4:0] c00415,c01415,c02415;
wire signed [4:0] c00425,c01425,c02425;
wire signed [4:0] c00435,c01435,c02435;
wire signed [4:0] c00445,c01445,c02445;
wire signed [4:0] c00006,c01006,c02006;
wire signed [4:0] c00016,c01016,c02016;
wire signed [4:0] c00026,c01026,c02026;
wire signed [4:0] c00036,c01036,c02036;
wire signed [4:0] c00046,c01046,c02046;
wire signed [4:0] c00106,c01106,c02106;
wire signed [4:0] c00116,c01116,c02116;
wire signed [4:0] c00126,c01126,c02126;
wire signed [4:0] c00136,c01136,c02136;
wire signed [4:0] c00146,c01146,c02146;
wire signed [4:0] c00206,c01206,c02206;
wire signed [4:0] c00216,c01216,c02216;
wire signed [4:0] c00226,c01226,c02226;
wire signed [4:0] c00236,c01236,c02236;
wire signed [4:0] c00246,c01246,c02246;
wire signed [4:0] c00306,c01306,c02306;
wire signed [4:0] c00316,c01316,c02316;
wire signed [4:0] c00326,c01326,c02326;
wire signed [4:0] c00336,c01336,c02336;
wire signed [4:0] c00346,c01346,c02346;
wire signed [4:0] c00406,c01406,c02406;
wire signed [4:0] c00416,c01416,c02416;
wire signed [4:0] c00426,c01426,c02426;
wire signed [4:0] c00436,c01436,c02436;
wire signed [4:0] c00446,c01446,c02446;
wire signed [4:0] c00007,c01007,c02007;
wire signed [4:0] c00017,c01017,c02017;
wire signed [4:0] c00027,c01027,c02027;
wire signed [4:0] c00037,c01037,c02037;
wire signed [4:0] c00047,c01047,c02047;
wire signed [4:0] c00107,c01107,c02107;
wire signed [4:0] c00117,c01117,c02117;
wire signed [4:0] c00127,c01127,c02127;
wire signed [4:0] c00137,c01137,c02137;
wire signed [4:0] c00147,c01147,c02147;
wire signed [4:0] c00207,c01207,c02207;
wire signed [4:0] c00217,c01217,c02217;
wire signed [4:0] c00227,c01227,c02227;
wire signed [4:0] c00237,c01237,c02237;
wire signed [4:0] c00247,c01247,c02247;
wire signed [4:0] c00307,c01307,c02307;
wire signed [4:0] c00317,c01317,c02317;
wire signed [4:0] c00327,c01327,c02327;
wire signed [4:0] c00337,c01337,c02337;
wire signed [4:0] c00347,c01347,c02347;
wire signed [4:0] c00407,c01407,c02407;
wire signed [4:0] c00417,c01417,c02417;
wire signed [4:0] c00427,c01427,c02427;
wire signed [4:0] c00437,c01437,c02437;
wire signed [4:0] c00447,c01447,c02447;
wire signed [4:0] c00008,c01008,c02008;
wire signed [4:0] c00018,c01018,c02018;
wire signed [4:0] c00028,c01028,c02028;
wire signed [4:0] c00038,c01038,c02038;
wire signed [4:0] c00048,c01048,c02048;
wire signed [4:0] c00108,c01108,c02108;
wire signed [4:0] c00118,c01118,c02118;
wire signed [4:0] c00128,c01128,c02128;
wire signed [4:0] c00138,c01138,c02138;
wire signed [4:0] c00148,c01148,c02148;
wire signed [4:0] c00208,c01208,c02208;
wire signed [4:0] c00218,c01218,c02218;
wire signed [4:0] c00228,c01228,c02228;
wire signed [4:0] c00238,c01238,c02238;
wire signed [4:0] c00248,c01248,c02248;
wire signed [4:0] c00308,c01308,c02308;
wire signed [4:0] c00318,c01318,c02318;
wire signed [4:0] c00328,c01328,c02328;
wire signed [4:0] c00338,c01338,c02338;
wire signed [4:0] c00348,c01348,c02348;
wire signed [4:0] c00408,c01408,c02408;
wire signed [4:0] c00418,c01418,c02418;
wire signed [4:0] c00428,c01428,c02428;
wire signed [4:0] c00438,c01438,c02438;
wire signed [4:0] c00448,c01448,c02448;
wire signed [4:0] c00009,c01009,c02009;
wire signed [4:0] c00019,c01019,c02019;
wire signed [4:0] c00029,c01029,c02029;
wire signed [4:0] c00039,c01039,c02039;
wire signed [4:0] c00049,c01049,c02049;
wire signed [4:0] c00109,c01109,c02109;
wire signed [4:0] c00119,c01119,c02119;
wire signed [4:0] c00129,c01129,c02129;
wire signed [4:0] c00139,c01139,c02139;
wire signed [4:0] c00149,c01149,c02149;
wire signed [4:0] c00209,c01209,c02209;
wire signed [4:0] c00219,c01219,c02219;
wire signed [4:0] c00229,c01229,c02229;
wire signed [4:0] c00239,c01239,c02239;
wire signed [4:0] c00249,c01249,c02249;
wire signed [4:0] c00309,c01309,c02309;
wire signed [4:0] c00319,c01319,c02319;
wire signed [4:0] c00329,c01329,c02329;
wire signed [4:0] c00339,c01339,c02339;
wire signed [4:0] c00349,c01349,c02349;
wire signed [4:0] c00409,c01409,c02409;
wire signed [4:0] c00419,c01419,c02419;
wire signed [4:0] c00429,c01429,c02429;
wire signed [4:0] c00439,c01439,c02439;
wire signed [4:0] c00449,c01449,c02449;
wire signed [4:0] c0000A,c0100A,c0200A;
wire signed [4:0] c0001A,c0101A,c0201A;
wire signed [4:0] c0002A,c0102A,c0202A;
wire signed [4:0] c0003A,c0103A,c0203A;
wire signed [4:0] c0004A,c0104A,c0204A;
wire signed [4:0] c0010A,c0110A,c0210A;
wire signed [4:0] c0011A,c0111A,c0211A;
wire signed [4:0] c0012A,c0112A,c0212A;
wire signed [4:0] c0013A,c0113A,c0213A;
wire signed [4:0] c0014A,c0114A,c0214A;
wire signed [4:0] c0020A,c0120A,c0220A;
wire signed [4:0] c0021A,c0121A,c0221A;
wire signed [4:0] c0022A,c0122A,c0222A;
wire signed [4:0] c0023A,c0123A,c0223A;
wire signed [4:0] c0024A,c0124A,c0224A;
wire signed [4:0] c0030A,c0130A,c0230A;
wire signed [4:0] c0031A,c0131A,c0231A;
wire signed [4:0] c0032A,c0132A,c0232A;
wire signed [4:0] c0033A,c0133A,c0233A;
wire signed [4:0] c0034A,c0134A,c0234A;
wire signed [4:0] c0040A,c0140A,c0240A;
wire signed [4:0] c0041A,c0141A,c0241A;
wire signed [4:0] c0042A,c0142A,c0242A;
wire signed [4:0] c0043A,c0143A,c0243A;
wire signed [4:0] c0044A,c0144A,c0244A;
wire signed [4:0] c0000B,c0100B,c0200B;
wire signed [4:0] c0001B,c0101B,c0201B;
wire signed [4:0] c0002B,c0102B,c0202B;
wire signed [4:0] c0003B,c0103B,c0203B;
wire signed [4:0] c0004B,c0104B,c0204B;
wire signed [4:0] c0010B,c0110B,c0210B;
wire signed [4:0] c0011B,c0111B,c0211B;
wire signed [4:0] c0012B,c0112B,c0212B;
wire signed [4:0] c0013B,c0113B,c0213B;
wire signed [4:0] c0014B,c0114B,c0214B;
wire signed [4:0] c0020B,c0120B,c0220B;
wire signed [4:0] c0021B,c0121B,c0221B;
wire signed [4:0] c0022B,c0122B,c0222B;
wire signed [4:0] c0023B,c0123B,c0223B;
wire signed [4:0] c0024B,c0124B,c0224B;
wire signed [4:0] c0030B,c0130B,c0230B;
wire signed [4:0] c0031B,c0131B,c0231B;
wire signed [4:0] c0032B,c0132B,c0232B;
wire signed [4:0] c0033B,c0133B,c0233B;
wire signed [4:0] c0034B,c0134B,c0234B;
wire signed [4:0] c0040B,c0140B,c0240B;
wire signed [4:0] c0041B,c0141B,c0241B;
wire signed [4:0] c0042B,c0142B,c0242B;
wire signed [4:0] c0043B,c0143B,c0243B;
wire signed [4:0] c0044B,c0144B,c0244B;
wire signed [4:0] c0000C,c0100C,c0200C;
wire signed [4:0] c0001C,c0101C,c0201C;
wire signed [4:0] c0002C,c0102C,c0202C;
wire signed [4:0] c0003C,c0103C,c0203C;
wire signed [4:0] c0004C,c0104C,c0204C;
wire signed [4:0] c0010C,c0110C,c0210C;
wire signed [4:0] c0011C,c0111C,c0211C;
wire signed [4:0] c0012C,c0112C,c0212C;
wire signed [4:0] c0013C,c0113C,c0213C;
wire signed [4:0] c0014C,c0114C,c0214C;
wire signed [4:0] c0020C,c0120C,c0220C;
wire signed [4:0] c0021C,c0121C,c0221C;
wire signed [4:0] c0022C,c0122C,c0222C;
wire signed [4:0] c0023C,c0123C,c0223C;
wire signed [4:0] c0024C,c0124C,c0224C;
wire signed [4:0] c0030C,c0130C,c0230C;
wire signed [4:0] c0031C,c0131C,c0231C;
wire signed [4:0] c0032C,c0132C,c0232C;
wire signed [4:0] c0033C,c0133C,c0233C;
wire signed [4:0] c0034C,c0134C,c0234C;
wire signed [4:0] c0040C,c0140C,c0240C;
wire signed [4:0] c0041C,c0141C,c0241C;
wire signed [4:0] c0042C,c0142C,c0242C;
wire signed [4:0] c0043C,c0143C,c0243C;
wire signed [4:0] c0044C,c0144C,c0244C;
wire signed [4:0] c0000D,c0100D,c0200D;
wire signed [4:0] c0001D,c0101D,c0201D;
wire signed [4:0] c0002D,c0102D,c0202D;
wire signed [4:0] c0003D,c0103D,c0203D;
wire signed [4:0] c0004D,c0104D,c0204D;
wire signed [4:0] c0010D,c0110D,c0210D;
wire signed [4:0] c0011D,c0111D,c0211D;
wire signed [4:0] c0012D,c0112D,c0212D;
wire signed [4:0] c0013D,c0113D,c0213D;
wire signed [4:0] c0014D,c0114D,c0214D;
wire signed [4:0] c0020D,c0120D,c0220D;
wire signed [4:0] c0021D,c0121D,c0221D;
wire signed [4:0] c0022D,c0122D,c0222D;
wire signed [4:0] c0023D,c0123D,c0223D;
wire signed [4:0] c0024D,c0124D,c0224D;
wire signed [4:0] c0030D,c0130D,c0230D;
wire signed [4:0] c0031D,c0131D,c0231D;
wire signed [4:0] c0032D,c0132D,c0232D;
wire signed [4:0] c0033D,c0133D,c0233D;
wire signed [4:0] c0034D,c0134D,c0234D;
wire signed [4:0] c0040D,c0140D,c0240D;
wire signed [4:0] c0041D,c0141D,c0241D;
wire signed [4:0] c0042D,c0142D,c0242D;
wire signed [4:0] c0043D,c0143D,c0243D;
wire signed [4:0] c0044D,c0144D,c0244D;
wire signed [4:0] c0000E,c0100E,c0200E;
wire signed [4:0] c0001E,c0101E,c0201E;
wire signed [4:0] c0002E,c0102E,c0202E;
wire signed [4:0] c0003E,c0103E,c0203E;
wire signed [4:0] c0004E,c0104E,c0204E;
wire signed [4:0] c0010E,c0110E,c0210E;
wire signed [4:0] c0011E,c0111E,c0211E;
wire signed [4:0] c0012E,c0112E,c0212E;
wire signed [4:0] c0013E,c0113E,c0213E;
wire signed [4:0] c0014E,c0114E,c0214E;
wire signed [4:0] c0020E,c0120E,c0220E;
wire signed [4:0] c0021E,c0121E,c0221E;
wire signed [4:0] c0022E,c0122E,c0222E;
wire signed [4:0] c0023E,c0123E,c0223E;
wire signed [4:0] c0024E,c0124E,c0224E;
wire signed [4:0] c0030E,c0130E,c0230E;
wire signed [4:0] c0031E,c0131E,c0231E;
wire signed [4:0] c0032E,c0132E,c0232E;
wire signed [4:0] c0033E,c0133E,c0233E;
wire signed [4:0] c0034E,c0134E,c0234E;
wire signed [4:0] c0040E,c0140E,c0240E;
wire signed [4:0] c0041E,c0141E,c0241E;
wire signed [4:0] c0042E,c0142E,c0242E;
wire signed [4:0] c0043E,c0143E,c0243E;
wire signed [4:0] c0044E,c0144E,c0244E;
wire signed [4:0] c0000F,c0100F,c0200F;
wire signed [4:0] c0001F,c0101F,c0201F;
wire signed [4:0] c0002F,c0102F,c0202F;
wire signed [4:0] c0003F,c0103F,c0203F;
wire signed [4:0] c0004F,c0104F,c0204F;
wire signed [4:0] c0010F,c0110F,c0210F;
wire signed [4:0] c0011F,c0111F,c0211F;
wire signed [4:0] c0012F,c0112F,c0212F;
wire signed [4:0] c0013F,c0113F,c0213F;
wire signed [4:0] c0014F,c0114F,c0214F;
wire signed [4:0] c0020F,c0120F,c0220F;
wire signed [4:0] c0021F,c0121F,c0221F;
wire signed [4:0] c0022F,c0122F,c0222F;
wire signed [4:0] c0023F,c0123F,c0223F;
wire signed [4:0] c0024F,c0124F,c0224F;
wire signed [4:0] c0030F,c0130F,c0230F;
wire signed [4:0] c0031F,c0131F,c0231F;
wire signed [4:0] c0032F,c0132F,c0232F;
wire signed [4:0] c0033F,c0133F,c0233F;
wire signed [4:0] c0034F,c0134F,c0234F;
wire signed [4:0] c0040F,c0140F,c0240F;
wire signed [4:0] c0041F,c0141F,c0241F;
wire signed [4:0] c0042F,c0142F,c0242F;
wire signed [4:0] c0043F,c0143F,c0243F;
wire signed [4:0] c0044F,c0144F,c0244F;
wire signed [6:0] C0000;
wire A0000;
wire signed [6:0] C0010;
wire A0010;
wire signed [6:0] C0020;
wire A0020;
wire signed [6:0] C0030;
wire A0030;
wire signed [6:0] C0040;
wire A0040;
wire signed [6:0] C0100;
wire A0100;
wire signed [6:0] C0110;
wire A0110;
wire signed [6:0] C0120;
wire A0120;
wire signed [6:0] C0130;
wire A0130;
wire signed [6:0] C0140;
wire A0140;
wire signed [6:0] C0200;
wire A0200;
wire signed [6:0] C0210;
wire A0210;
wire signed [6:0] C0220;
wire A0220;
wire signed [6:0] C0230;
wire A0230;
wire signed [6:0] C0240;
wire A0240;
wire signed [6:0] C0300;
wire A0300;
wire signed [6:0] C0310;
wire A0310;
wire signed [6:0] C0320;
wire A0320;
wire signed [6:0] C0330;
wire A0330;
wire signed [6:0] C0340;
wire A0340;
wire signed [6:0] C0400;
wire A0400;
wire signed [6:0] C0410;
wire A0410;
wire signed [6:0] C0420;
wire A0420;
wire signed [6:0] C0430;
wire A0430;
wire signed [6:0] C0440;
wire A0440;
wire signed [6:0] C0001;
wire A0001;
wire signed [6:0] C0011;
wire A0011;
wire signed [6:0] C0021;
wire A0021;
wire signed [6:0] C0031;
wire A0031;
wire signed [6:0] C0041;
wire A0041;
wire signed [6:0] C0101;
wire A0101;
wire signed [6:0] C0111;
wire A0111;
wire signed [6:0] C0121;
wire A0121;
wire signed [6:0] C0131;
wire A0131;
wire signed [6:0] C0141;
wire A0141;
wire signed [6:0] C0201;
wire A0201;
wire signed [6:0] C0211;
wire A0211;
wire signed [6:0] C0221;
wire A0221;
wire signed [6:0] C0231;
wire A0231;
wire signed [6:0] C0241;
wire A0241;
wire signed [6:0] C0301;
wire A0301;
wire signed [6:0] C0311;
wire A0311;
wire signed [6:0] C0321;
wire A0321;
wire signed [6:0] C0331;
wire A0331;
wire signed [6:0] C0341;
wire A0341;
wire signed [6:0] C0401;
wire A0401;
wire signed [6:0] C0411;
wire A0411;
wire signed [6:0] C0421;
wire A0421;
wire signed [6:0] C0431;
wire A0431;
wire signed [6:0] C0441;
wire A0441;
wire signed [6:0] C0002;
wire A0002;
wire signed [6:0] C0012;
wire A0012;
wire signed [6:0] C0022;
wire A0022;
wire signed [6:0] C0032;
wire A0032;
wire signed [6:0] C0042;
wire A0042;
wire signed [6:0] C0102;
wire A0102;
wire signed [6:0] C0112;
wire A0112;
wire signed [6:0] C0122;
wire A0122;
wire signed [6:0] C0132;
wire A0132;
wire signed [6:0] C0142;
wire A0142;
wire signed [6:0] C0202;
wire A0202;
wire signed [6:0] C0212;
wire A0212;
wire signed [6:0] C0222;
wire A0222;
wire signed [6:0] C0232;
wire A0232;
wire signed [6:0] C0242;
wire A0242;
wire signed [6:0] C0302;
wire A0302;
wire signed [6:0] C0312;
wire A0312;
wire signed [6:0] C0322;
wire A0322;
wire signed [6:0] C0332;
wire A0332;
wire signed [6:0] C0342;
wire A0342;
wire signed [6:0] C0402;
wire A0402;
wire signed [6:0] C0412;
wire A0412;
wire signed [6:0] C0422;
wire A0422;
wire signed [6:0] C0432;
wire A0432;
wire signed [6:0] C0442;
wire A0442;
wire signed [6:0] C0003;
wire A0003;
wire signed [6:0] C0013;
wire A0013;
wire signed [6:0] C0023;
wire A0023;
wire signed [6:0] C0033;
wire A0033;
wire signed [6:0] C0043;
wire A0043;
wire signed [6:0] C0103;
wire A0103;
wire signed [6:0] C0113;
wire A0113;
wire signed [6:0] C0123;
wire A0123;
wire signed [6:0] C0133;
wire A0133;
wire signed [6:0] C0143;
wire A0143;
wire signed [6:0] C0203;
wire A0203;
wire signed [6:0] C0213;
wire A0213;
wire signed [6:0] C0223;
wire A0223;
wire signed [6:0] C0233;
wire A0233;
wire signed [6:0] C0243;
wire A0243;
wire signed [6:0] C0303;
wire A0303;
wire signed [6:0] C0313;
wire A0313;
wire signed [6:0] C0323;
wire A0323;
wire signed [6:0] C0333;
wire A0333;
wire signed [6:0] C0343;
wire A0343;
wire signed [6:0] C0403;
wire A0403;
wire signed [6:0] C0413;
wire A0413;
wire signed [6:0] C0423;
wire A0423;
wire signed [6:0] C0433;
wire A0433;
wire signed [6:0] C0443;
wire A0443;
wire signed [6:0] C0004;
wire A0004;
wire signed [6:0] C0014;
wire A0014;
wire signed [6:0] C0024;
wire A0024;
wire signed [6:0] C0034;
wire A0034;
wire signed [6:0] C0044;
wire A0044;
wire signed [6:0] C0104;
wire A0104;
wire signed [6:0] C0114;
wire A0114;
wire signed [6:0] C0124;
wire A0124;
wire signed [6:0] C0134;
wire A0134;
wire signed [6:0] C0144;
wire A0144;
wire signed [6:0] C0204;
wire A0204;
wire signed [6:0] C0214;
wire A0214;
wire signed [6:0] C0224;
wire A0224;
wire signed [6:0] C0234;
wire A0234;
wire signed [6:0] C0244;
wire A0244;
wire signed [6:0] C0304;
wire A0304;
wire signed [6:0] C0314;
wire A0314;
wire signed [6:0] C0324;
wire A0324;
wire signed [6:0] C0334;
wire A0334;
wire signed [6:0] C0344;
wire A0344;
wire signed [6:0] C0404;
wire A0404;
wire signed [6:0] C0414;
wire A0414;
wire signed [6:0] C0424;
wire A0424;
wire signed [6:0] C0434;
wire A0434;
wire signed [6:0] C0444;
wire A0444;
wire signed [6:0] C0005;
wire A0005;
wire signed [6:0] C0015;
wire A0015;
wire signed [6:0] C0025;
wire A0025;
wire signed [6:0] C0035;
wire A0035;
wire signed [6:0] C0045;
wire A0045;
wire signed [6:0] C0105;
wire A0105;
wire signed [6:0] C0115;
wire A0115;
wire signed [6:0] C0125;
wire A0125;
wire signed [6:0] C0135;
wire A0135;
wire signed [6:0] C0145;
wire A0145;
wire signed [6:0] C0205;
wire A0205;
wire signed [6:0] C0215;
wire A0215;
wire signed [6:0] C0225;
wire A0225;
wire signed [6:0] C0235;
wire A0235;
wire signed [6:0] C0245;
wire A0245;
wire signed [6:0] C0305;
wire A0305;
wire signed [6:0] C0315;
wire A0315;
wire signed [6:0] C0325;
wire A0325;
wire signed [6:0] C0335;
wire A0335;
wire signed [6:0] C0345;
wire A0345;
wire signed [6:0] C0405;
wire A0405;
wire signed [6:0] C0415;
wire A0415;
wire signed [6:0] C0425;
wire A0425;
wire signed [6:0] C0435;
wire A0435;
wire signed [6:0] C0445;
wire A0445;
wire signed [6:0] C0006;
wire A0006;
wire signed [6:0] C0016;
wire A0016;
wire signed [6:0] C0026;
wire A0026;
wire signed [6:0] C0036;
wire A0036;
wire signed [6:0] C0046;
wire A0046;
wire signed [6:0] C0106;
wire A0106;
wire signed [6:0] C0116;
wire A0116;
wire signed [6:0] C0126;
wire A0126;
wire signed [6:0] C0136;
wire A0136;
wire signed [6:0] C0146;
wire A0146;
wire signed [6:0] C0206;
wire A0206;
wire signed [6:0] C0216;
wire A0216;
wire signed [6:0] C0226;
wire A0226;
wire signed [6:0] C0236;
wire A0236;
wire signed [6:0] C0246;
wire A0246;
wire signed [6:0] C0306;
wire A0306;
wire signed [6:0] C0316;
wire A0316;
wire signed [6:0] C0326;
wire A0326;
wire signed [6:0] C0336;
wire A0336;
wire signed [6:0] C0346;
wire A0346;
wire signed [6:0] C0406;
wire A0406;
wire signed [6:0] C0416;
wire A0416;
wire signed [6:0] C0426;
wire A0426;
wire signed [6:0] C0436;
wire A0436;
wire signed [6:0] C0446;
wire A0446;
wire signed [6:0] C0007;
wire A0007;
wire signed [6:0] C0017;
wire A0017;
wire signed [6:0] C0027;
wire A0027;
wire signed [6:0] C0037;
wire A0037;
wire signed [6:0] C0047;
wire A0047;
wire signed [6:0] C0107;
wire A0107;
wire signed [6:0] C0117;
wire A0117;
wire signed [6:0] C0127;
wire A0127;
wire signed [6:0] C0137;
wire A0137;
wire signed [6:0] C0147;
wire A0147;
wire signed [6:0] C0207;
wire A0207;
wire signed [6:0] C0217;
wire A0217;
wire signed [6:0] C0227;
wire A0227;
wire signed [6:0] C0237;
wire A0237;
wire signed [6:0] C0247;
wire A0247;
wire signed [6:0] C0307;
wire A0307;
wire signed [6:0] C0317;
wire A0317;
wire signed [6:0] C0327;
wire A0327;
wire signed [6:0] C0337;
wire A0337;
wire signed [6:0] C0347;
wire A0347;
wire signed [6:0] C0407;
wire A0407;
wire signed [6:0] C0417;
wire A0417;
wire signed [6:0] C0427;
wire A0427;
wire signed [6:0] C0437;
wire A0437;
wire signed [6:0] C0447;
wire A0447;
wire signed [6:0] C0008;
wire A0008;
wire signed [6:0] C0018;
wire A0018;
wire signed [6:0] C0028;
wire A0028;
wire signed [6:0] C0038;
wire A0038;
wire signed [6:0] C0048;
wire A0048;
wire signed [6:0] C0108;
wire A0108;
wire signed [6:0] C0118;
wire A0118;
wire signed [6:0] C0128;
wire A0128;
wire signed [6:0] C0138;
wire A0138;
wire signed [6:0] C0148;
wire A0148;
wire signed [6:0] C0208;
wire A0208;
wire signed [6:0] C0218;
wire A0218;
wire signed [6:0] C0228;
wire A0228;
wire signed [6:0] C0238;
wire A0238;
wire signed [6:0] C0248;
wire A0248;
wire signed [6:0] C0308;
wire A0308;
wire signed [6:0] C0318;
wire A0318;
wire signed [6:0] C0328;
wire A0328;
wire signed [6:0] C0338;
wire A0338;
wire signed [6:0] C0348;
wire A0348;
wire signed [6:0] C0408;
wire A0408;
wire signed [6:0] C0418;
wire A0418;
wire signed [6:0] C0428;
wire A0428;
wire signed [6:0] C0438;
wire A0438;
wire signed [6:0] C0448;
wire A0448;
wire signed [6:0] C0009;
wire A0009;
wire signed [6:0] C0019;
wire A0019;
wire signed [6:0] C0029;
wire A0029;
wire signed [6:0] C0039;
wire A0039;
wire signed [6:0] C0049;
wire A0049;
wire signed [6:0] C0109;
wire A0109;
wire signed [6:0] C0119;
wire A0119;
wire signed [6:0] C0129;
wire A0129;
wire signed [6:0] C0139;
wire A0139;
wire signed [6:0] C0149;
wire A0149;
wire signed [6:0] C0209;
wire A0209;
wire signed [6:0] C0219;
wire A0219;
wire signed [6:0] C0229;
wire A0229;
wire signed [6:0] C0239;
wire A0239;
wire signed [6:0] C0249;
wire A0249;
wire signed [6:0] C0309;
wire A0309;
wire signed [6:0] C0319;
wire A0319;
wire signed [6:0] C0329;
wire A0329;
wire signed [6:0] C0339;
wire A0339;
wire signed [6:0] C0349;
wire A0349;
wire signed [6:0] C0409;
wire A0409;
wire signed [6:0] C0419;
wire A0419;
wire signed [6:0] C0429;
wire A0429;
wire signed [6:0] C0439;
wire A0439;
wire signed [6:0] C0449;
wire A0449;
wire signed [6:0] C000A;
wire A000A;
wire signed [6:0] C001A;
wire A001A;
wire signed [6:0] C002A;
wire A002A;
wire signed [6:0] C003A;
wire A003A;
wire signed [6:0] C004A;
wire A004A;
wire signed [6:0] C010A;
wire A010A;
wire signed [6:0] C011A;
wire A011A;
wire signed [6:0] C012A;
wire A012A;
wire signed [6:0] C013A;
wire A013A;
wire signed [6:0] C014A;
wire A014A;
wire signed [6:0] C020A;
wire A020A;
wire signed [6:0] C021A;
wire A021A;
wire signed [6:0] C022A;
wire A022A;
wire signed [6:0] C023A;
wire A023A;
wire signed [6:0] C024A;
wire A024A;
wire signed [6:0] C030A;
wire A030A;
wire signed [6:0] C031A;
wire A031A;
wire signed [6:0] C032A;
wire A032A;
wire signed [6:0] C033A;
wire A033A;
wire signed [6:0] C034A;
wire A034A;
wire signed [6:0] C040A;
wire A040A;
wire signed [6:0] C041A;
wire A041A;
wire signed [6:0] C042A;
wire A042A;
wire signed [6:0] C043A;
wire A043A;
wire signed [6:0] C044A;
wire A044A;
wire signed [6:0] C000B;
wire A000B;
wire signed [6:0] C001B;
wire A001B;
wire signed [6:0] C002B;
wire A002B;
wire signed [6:0] C003B;
wire A003B;
wire signed [6:0] C004B;
wire A004B;
wire signed [6:0] C010B;
wire A010B;
wire signed [6:0] C011B;
wire A011B;
wire signed [6:0] C012B;
wire A012B;
wire signed [6:0] C013B;
wire A013B;
wire signed [6:0] C014B;
wire A014B;
wire signed [6:0] C020B;
wire A020B;
wire signed [6:0] C021B;
wire A021B;
wire signed [6:0] C022B;
wire A022B;
wire signed [6:0] C023B;
wire A023B;
wire signed [6:0] C024B;
wire A024B;
wire signed [6:0] C030B;
wire A030B;
wire signed [6:0] C031B;
wire A031B;
wire signed [6:0] C032B;
wire A032B;
wire signed [6:0] C033B;
wire A033B;
wire signed [6:0] C034B;
wire A034B;
wire signed [6:0] C040B;
wire A040B;
wire signed [6:0] C041B;
wire A041B;
wire signed [6:0] C042B;
wire A042B;
wire signed [6:0] C043B;
wire A043B;
wire signed [6:0] C044B;
wire A044B;
wire signed [6:0] C000C;
wire A000C;
wire signed [6:0] C001C;
wire A001C;
wire signed [6:0] C002C;
wire A002C;
wire signed [6:0] C003C;
wire A003C;
wire signed [6:0] C004C;
wire A004C;
wire signed [6:0] C010C;
wire A010C;
wire signed [6:0] C011C;
wire A011C;
wire signed [6:0] C012C;
wire A012C;
wire signed [6:0] C013C;
wire A013C;
wire signed [6:0] C014C;
wire A014C;
wire signed [6:0] C020C;
wire A020C;
wire signed [6:0] C021C;
wire A021C;
wire signed [6:0] C022C;
wire A022C;
wire signed [6:0] C023C;
wire A023C;
wire signed [6:0] C024C;
wire A024C;
wire signed [6:0] C030C;
wire A030C;
wire signed [6:0] C031C;
wire A031C;
wire signed [6:0] C032C;
wire A032C;
wire signed [6:0] C033C;
wire A033C;
wire signed [6:0] C034C;
wire A034C;
wire signed [6:0] C040C;
wire A040C;
wire signed [6:0] C041C;
wire A041C;
wire signed [6:0] C042C;
wire A042C;
wire signed [6:0] C043C;
wire A043C;
wire signed [6:0] C044C;
wire A044C;
wire signed [6:0] C000D;
wire A000D;
wire signed [6:0] C001D;
wire A001D;
wire signed [6:0] C002D;
wire A002D;
wire signed [6:0] C003D;
wire A003D;
wire signed [6:0] C004D;
wire A004D;
wire signed [6:0] C010D;
wire A010D;
wire signed [6:0] C011D;
wire A011D;
wire signed [6:0] C012D;
wire A012D;
wire signed [6:0] C013D;
wire A013D;
wire signed [6:0] C014D;
wire A014D;
wire signed [6:0] C020D;
wire A020D;
wire signed [6:0] C021D;
wire A021D;
wire signed [6:0] C022D;
wire A022D;
wire signed [6:0] C023D;
wire A023D;
wire signed [6:0] C024D;
wire A024D;
wire signed [6:0] C030D;
wire A030D;
wire signed [6:0] C031D;
wire A031D;
wire signed [6:0] C032D;
wire A032D;
wire signed [6:0] C033D;
wire A033D;
wire signed [6:0] C034D;
wire A034D;
wire signed [6:0] C040D;
wire A040D;
wire signed [6:0] C041D;
wire A041D;
wire signed [6:0] C042D;
wire A042D;
wire signed [6:0] C043D;
wire A043D;
wire signed [6:0] C044D;
wire A044D;
wire signed [6:0] C000E;
wire A000E;
wire signed [6:0] C001E;
wire A001E;
wire signed [6:0] C002E;
wire A002E;
wire signed [6:0] C003E;
wire A003E;
wire signed [6:0] C004E;
wire A004E;
wire signed [6:0] C010E;
wire A010E;
wire signed [6:0] C011E;
wire A011E;
wire signed [6:0] C012E;
wire A012E;
wire signed [6:0] C013E;
wire A013E;
wire signed [6:0] C014E;
wire A014E;
wire signed [6:0] C020E;
wire A020E;
wire signed [6:0] C021E;
wire A021E;
wire signed [6:0] C022E;
wire A022E;
wire signed [6:0] C023E;
wire A023E;
wire signed [6:0] C024E;
wire A024E;
wire signed [6:0] C030E;
wire A030E;
wire signed [6:0] C031E;
wire A031E;
wire signed [6:0] C032E;
wire A032E;
wire signed [6:0] C033E;
wire A033E;
wire signed [6:0] C034E;
wire A034E;
wire signed [6:0] C040E;
wire A040E;
wire signed [6:0] C041E;
wire A041E;
wire signed [6:0] C042E;
wire A042E;
wire signed [6:0] C043E;
wire A043E;
wire signed [6:0] C044E;
wire A044E;
wire signed [6:0] C000F;
wire A000F;
wire signed [6:0] C001F;
wire A001F;
wire signed [6:0] C002F;
wire A002F;
wire signed [6:0] C003F;
wire A003F;
wire signed [6:0] C004F;
wire A004F;
wire signed [6:0] C010F;
wire A010F;
wire signed [6:0] C011F;
wire A011F;
wire signed [6:0] C012F;
wire A012F;
wire signed [6:0] C013F;
wire A013F;
wire signed [6:0] C014F;
wire A014F;
wire signed [6:0] C020F;
wire A020F;
wire signed [6:0] C021F;
wire A021F;
wire signed [6:0] C022F;
wire A022F;
wire signed [6:0] C023F;
wire A023F;
wire signed [6:0] C024F;
wire A024F;
wire signed [6:0] C030F;
wire A030F;
wire signed [6:0] C031F;
wire A031F;
wire signed [6:0] C032F;
wire A032F;
wire signed [6:0] C033F;
wire A033F;
wire signed [6:0] C034F;
wire A034F;
wire signed [6:0] C040F;
wire A040F;
wire signed [6:0] C041F;
wire A041F;
wire signed [6:0] C042F;
wire A042F;
wire signed [6:0] C043F;
wire A043F;
wire signed [6:0] C044F;
wire A044F;
DFF_save_fm DFF_P0(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0000));
DFF_save_fm DFF_P1(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0010));
DFF_save_fm DFF_P2(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0020));
DFF_save_fm DFF_P3(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0030));
DFF_save_fm DFF_P4(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0040));
DFF_save_fm DFF_P5(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0050));
DFF_save_fm DFF_P6(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0060));
DFF_save_fm DFF_P7(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0100));
DFF_save_fm DFF_P8(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0110));
DFF_save_fm DFF_P9(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0120));
DFF_save_fm DFF_P10(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0130));
DFF_save_fm DFF_P11(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0140));
DFF_save_fm DFF_P12(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0150));
DFF_save_fm DFF_P13(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0160));
DFF_save_fm DFF_P14(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0200));
DFF_save_fm DFF_P15(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0210));
DFF_save_fm DFF_P16(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0220));
DFF_save_fm DFF_P17(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0230));
DFF_save_fm DFF_P18(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0240));
DFF_save_fm DFF_P19(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0250));
DFF_save_fm DFF_P20(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0260));
DFF_save_fm DFF_P21(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0300));
DFF_save_fm DFF_P22(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0310));
DFF_save_fm DFF_P23(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0320));
DFF_save_fm DFF_P24(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0330));
DFF_save_fm DFF_P25(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0340));
DFF_save_fm DFF_P26(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0350));
DFF_save_fm DFF_P27(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0360));
DFF_save_fm DFF_P28(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0400));
DFF_save_fm DFF_P29(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0410));
DFF_save_fm DFF_P30(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0420));
DFF_save_fm DFF_P31(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0430));
DFF_save_fm DFF_P32(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0440));
DFF_save_fm DFF_P33(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0450));
DFF_save_fm DFF_P34(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0460));
DFF_save_fm DFF_P35(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0500));
DFF_save_fm DFF_P36(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0510));
DFF_save_fm DFF_P37(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0520));
DFF_save_fm DFF_P38(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0530));
DFF_save_fm DFF_P39(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0540));
DFF_save_fm DFF_P40(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0550));
DFF_save_fm DFF_P41(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0560));
DFF_save_fm DFF_P42(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0600));
DFF_save_fm DFF_P43(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0610));
DFF_save_fm DFF_P44(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0620));
DFF_save_fm DFF_P45(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0630));
DFF_save_fm DFF_P46(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0640));
DFF_save_fm DFF_P47(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0650));
DFF_save_fm DFF_P48(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0660));
DFF_save_fm DFF_P49(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0001));
DFF_save_fm DFF_P50(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0011));
DFF_save_fm DFF_P51(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0021));
DFF_save_fm DFF_P52(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0031));
DFF_save_fm DFF_P53(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0041));
DFF_save_fm DFF_P54(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0051));
DFF_save_fm DFF_P55(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0061));
DFF_save_fm DFF_P56(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0101));
DFF_save_fm DFF_P57(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0111));
DFF_save_fm DFF_P58(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0121));
DFF_save_fm DFF_P59(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0131));
DFF_save_fm DFF_P60(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0141));
DFF_save_fm DFF_P61(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0151));
DFF_save_fm DFF_P62(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0161));
DFF_save_fm DFF_P63(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0201));
DFF_save_fm DFF_P64(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0211));
DFF_save_fm DFF_P65(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0221));
DFF_save_fm DFF_P66(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0231));
DFF_save_fm DFF_P67(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0241));
DFF_save_fm DFF_P68(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0251));
DFF_save_fm DFF_P69(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0261));
DFF_save_fm DFF_P70(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0301));
DFF_save_fm DFF_P71(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0311));
DFF_save_fm DFF_P72(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0321));
DFF_save_fm DFF_P73(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0331));
DFF_save_fm DFF_P74(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0341));
DFF_save_fm DFF_P75(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0351));
DFF_save_fm DFF_P76(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0361));
DFF_save_fm DFF_P77(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0401));
DFF_save_fm DFF_P78(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0411));
DFF_save_fm DFF_P79(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0421));
DFF_save_fm DFF_P80(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0431));
DFF_save_fm DFF_P81(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0441));
DFF_save_fm DFF_P82(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0451));
DFF_save_fm DFF_P83(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0461));
DFF_save_fm DFF_P84(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0501));
DFF_save_fm DFF_P85(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0511));
DFF_save_fm DFF_P86(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0521));
DFF_save_fm DFF_P87(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0531));
DFF_save_fm DFF_P88(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0541));
DFF_save_fm DFF_P89(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0551));
DFF_save_fm DFF_P90(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0561));
DFF_save_fm DFF_P91(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0601));
DFF_save_fm DFF_P92(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0611));
DFF_save_fm DFF_P93(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0621));
DFF_save_fm DFF_P94(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0631));
DFF_save_fm DFF_P95(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0641));
DFF_save_fm DFF_P96(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0651));
DFF_save_fm DFF_P97(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0661));
DFF_save_fm DFF_P98(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0002));
DFF_save_fm DFF_P99(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0012));
DFF_save_fm DFF_P100(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0022));
DFF_save_fm DFF_P101(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0032));
DFF_save_fm DFF_P102(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0042));
DFF_save_fm DFF_P103(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0052));
DFF_save_fm DFF_P104(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0062));
DFF_save_fm DFF_P105(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0102));
DFF_save_fm DFF_P106(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0112));
DFF_save_fm DFF_P107(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0122));
DFF_save_fm DFF_P108(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0132));
DFF_save_fm DFF_P109(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0142));
DFF_save_fm DFF_P110(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0152));
DFF_save_fm DFF_P111(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0162));
DFF_save_fm DFF_P112(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0202));
DFF_save_fm DFF_P113(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0212));
DFF_save_fm DFF_P114(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0222));
DFF_save_fm DFF_P115(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0232));
DFF_save_fm DFF_P116(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0242));
DFF_save_fm DFF_P117(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0252));
DFF_save_fm DFF_P118(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0262));
DFF_save_fm DFF_P119(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0302));
DFF_save_fm DFF_P120(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0312));
DFF_save_fm DFF_P121(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0322));
DFF_save_fm DFF_P122(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0332));
DFF_save_fm DFF_P123(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0342));
DFF_save_fm DFF_P124(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0352));
DFF_save_fm DFF_P125(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0362));
DFF_save_fm DFF_P126(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0402));
DFF_save_fm DFF_P127(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0412));
DFF_save_fm DFF_P128(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0422));
DFF_save_fm DFF_P129(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0432));
DFF_save_fm DFF_P130(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0442));
DFF_save_fm DFF_P131(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0452));
DFF_save_fm DFF_P132(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0462));
DFF_save_fm DFF_P133(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0502));
DFF_save_fm DFF_P134(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0512));
DFF_save_fm DFF_P135(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0522));
DFF_save_fm DFF_P136(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0532));
DFF_save_fm DFF_P137(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0542));
DFF_save_fm DFF_P138(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0552));
DFF_save_fm DFF_P139(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0562));
DFF_save_fm DFF_P140(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0602));
DFF_save_fm DFF_P141(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0612));
DFF_save_fm DFF_P142(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0622));
DFF_save_fm DFF_P143(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0632));
DFF_save_fm DFF_P144(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0642));
DFF_save_fm DFF_P145(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0652));
DFF_save_fm DFF_P146(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0662));
DFF_save_fm DFF_W0(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00000));
DFF_save_fm DFF_W1(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00010));
DFF_save_fm DFF_W2(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00020));
DFF_save_fm DFF_W3(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00100));
DFF_save_fm DFF_W4(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00110));
DFF_save_fm DFF_W5(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00120));
DFF_save_fm DFF_W6(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00200));
DFF_save_fm DFF_W7(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00210));
DFF_save_fm DFF_W8(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00220));
DFF_save_fm DFF_W9(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00001));
DFF_save_fm DFF_W10(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00011));
DFF_save_fm DFF_W11(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00021));
DFF_save_fm DFF_W12(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00101));
DFF_save_fm DFF_W13(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00111));
DFF_save_fm DFF_W14(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00121));
DFF_save_fm DFF_W15(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00201));
DFF_save_fm DFF_W16(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00211));
DFF_save_fm DFF_W17(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00221));
DFF_save_fm DFF_W18(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00002));
DFF_save_fm DFF_W19(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00012));
DFF_save_fm DFF_W20(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00022));
DFF_save_fm DFF_W21(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00102));
DFF_save_fm DFF_W22(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00112));
DFF_save_fm DFF_W23(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00122));
DFF_save_fm DFF_W24(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00202));
DFF_save_fm DFF_W25(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00212));
DFF_save_fm DFF_W26(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00222));
DFF_save_fm DFF_W27(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01000));
DFF_save_fm DFF_W28(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01010));
DFF_save_fm DFF_W29(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01020));
DFF_save_fm DFF_W30(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01100));
DFF_save_fm DFF_W31(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01110));
DFF_save_fm DFF_W32(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01120));
DFF_save_fm DFF_W33(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01200));
DFF_save_fm DFF_W34(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01210));
DFF_save_fm DFF_W35(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01220));
DFF_save_fm DFF_W36(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01001));
DFF_save_fm DFF_W37(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01011));
DFF_save_fm DFF_W38(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01021));
DFF_save_fm DFF_W39(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01101));
DFF_save_fm DFF_W40(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01111));
DFF_save_fm DFF_W41(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01121));
DFF_save_fm DFF_W42(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01201));
DFF_save_fm DFF_W43(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01211));
DFF_save_fm DFF_W44(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01221));
DFF_save_fm DFF_W45(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01002));
DFF_save_fm DFF_W46(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01012));
DFF_save_fm DFF_W47(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01022));
DFF_save_fm DFF_W48(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01102));
DFF_save_fm DFF_W49(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01112));
DFF_save_fm DFF_W50(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01122));
DFF_save_fm DFF_W51(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01202));
DFF_save_fm DFF_W52(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01212));
DFF_save_fm DFF_W53(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01222));
DFF_save_fm DFF_W54(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02000));
DFF_save_fm DFF_W55(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02010));
DFF_save_fm DFF_W56(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02020));
DFF_save_fm DFF_W57(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02100));
DFF_save_fm DFF_W58(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02110));
DFF_save_fm DFF_W59(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02120));
DFF_save_fm DFF_W60(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02200));
DFF_save_fm DFF_W61(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02210));
DFF_save_fm DFF_W62(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02220));
DFF_save_fm DFF_W63(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02001));
DFF_save_fm DFF_W64(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02011));
DFF_save_fm DFF_W65(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02021));
DFF_save_fm DFF_W66(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02101));
DFF_save_fm DFF_W67(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02111));
DFF_save_fm DFF_W68(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02121));
DFF_save_fm DFF_W69(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02201));
DFF_save_fm DFF_W70(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02211));
DFF_save_fm DFF_W71(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02221));
DFF_save_fm DFF_W72(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02002));
DFF_save_fm DFF_W73(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02012));
DFF_save_fm DFF_W74(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02022));
DFF_save_fm DFF_W75(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02102));
DFF_save_fm DFF_W76(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02112));
DFF_save_fm DFF_W77(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02122));
DFF_save_fm DFF_W78(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02202));
DFF_save_fm DFF_W79(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02212));
DFF_save_fm DFF_W80(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02222));
DFF_save_fm DFF_W81(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03000));
DFF_save_fm DFF_W82(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03010));
DFF_save_fm DFF_W83(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03020));
DFF_save_fm DFF_W84(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03100));
DFF_save_fm DFF_W85(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03110));
DFF_save_fm DFF_W86(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03120));
DFF_save_fm DFF_W87(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03200));
DFF_save_fm DFF_W88(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03210));
DFF_save_fm DFF_W89(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03220));
DFF_save_fm DFF_W90(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03001));
DFF_save_fm DFF_W91(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03011));
DFF_save_fm DFF_W92(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03021));
DFF_save_fm DFF_W93(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03101));
DFF_save_fm DFF_W94(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03111));
DFF_save_fm DFF_W95(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03121));
DFF_save_fm DFF_W96(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03201));
DFF_save_fm DFF_W97(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03211));
DFF_save_fm DFF_W98(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03221));
DFF_save_fm DFF_W99(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03002));
DFF_save_fm DFF_W100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03012));
DFF_save_fm DFF_W101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03022));
DFF_save_fm DFF_W102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03102));
DFF_save_fm DFF_W103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03112));
DFF_save_fm DFF_W104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03122));
DFF_save_fm DFF_W105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03202));
DFF_save_fm DFF_W106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03212));
DFF_save_fm DFF_W107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03222));
DFF_save_fm DFF_W108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04000));
DFF_save_fm DFF_W109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04010));
DFF_save_fm DFF_W110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04020));
DFF_save_fm DFF_W111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04100));
DFF_save_fm DFF_W112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04110));
DFF_save_fm DFF_W113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04120));
DFF_save_fm DFF_W114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04200));
DFF_save_fm DFF_W115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04210));
DFF_save_fm DFF_W116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04220));
DFF_save_fm DFF_W117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04001));
DFF_save_fm DFF_W118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04011));
DFF_save_fm DFF_W119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04021));
DFF_save_fm DFF_W120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04101));
DFF_save_fm DFF_W121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04111));
DFF_save_fm DFF_W122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04121));
DFF_save_fm DFF_W123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04201));
DFF_save_fm DFF_W124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04211));
DFF_save_fm DFF_W125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04221));
DFF_save_fm DFF_W126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04002));
DFF_save_fm DFF_W127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04012));
DFF_save_fm DFF_W128(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04022));
DFF_save_fm DFF_W129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04102));
DFF_save_fm DFF_W130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W04112));
DFF_save_fm DFF_W131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04122));
DFF_save_fm DFF_W132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04202));
DFF_save_fm DFF_W133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04212));
DFF_save_fm DFF_W134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W04222));
DFF_save_fm DFF_W135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05000));
DFF_save_fm DFF_W136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05010));
DFF_save_fm DFF_W137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05020));
DFF_save_fm DFF_W138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05100));
DFF_save_fm DFF_W139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05110));
DFF_save_fm DFF_W140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05120));
DFF_save_fm DFF_W141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05200));
DFF_save_fm DFF_W142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05210));
DFF_save_fm DFF_W143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05220));
DFF_save_fm DFF_W144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05001));
DFF_save_fm DFF_W145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05011));
DFF_save_fm DFF_W146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05021));
DFF_save_fm DFF_W147(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05101));
DFF_save_fm DFF_W148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05111));
DFF_save_fm DFF_W149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05121));
DFF_save_fm DFF_W150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05201));
DFF_save_fm DFF_W151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05211));
DFF_save_fm DFF_W152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05221));
DFF_save_fm DFF_W153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05002));
DFF_save_fm DFF_W154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05012));
DFF_save_fm DFF_W155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05022));
DFF_save_fm DFF_W156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05102));
DFF_save_fm DFF_W157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05112));
DFF_save_fm DFF_W158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05122));
DFF_save_fm DFF_W159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05202));
DFF_save_fm DFF_W160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W05212));
DFF_save_fm DFF_W161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W05222));
DFF_save_fm DFF_W162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06000));
DFF_save_fm DFF_W163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06010));
DFF_save_fm DFF_W164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06020));
DFF_save_fm DFF_W165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06100));
DFF_save_fm DFF_W166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06110));
DFF_save_fm DFF_W167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06120));
DFF_save_fm DFF_W168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06200));
DFF_save_fm DFF_W169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06210));
DFF_save_fm DFF_W170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06220));
DFF_save_fm DFF_W171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06001));
DFF_save_fm DFF_W172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06011));
DFF_save_fm DFF_W173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06021));
DFF_save_fm DFF_W174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06101));
DFF_save_fm DFF_W175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06111));
DFF_save_fm DFF_W176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06121));
DFF_save_fm DFF_W177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06201));
DFF_save_fm DFF_W178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06211));
DFF_save_fm DFF_W179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06221));
DFF_save_fm DFF_W180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06002));
DFF_save_fm DFF_W181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06012));
DFF_save_fm DFF_W182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06022));
DFF_save_fm DFF_W183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06102));
DFF_save_fm DFF_W184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06112));
DFF_save_fm DFF_W185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W06122));
DFF_save_fm DFF_W186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06202));
DFF_save_fm DFF_W187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06212));
DFF_save_fm DFF_W188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W06222));
DFF_save_fm DFF_W189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07000));
DFF_save_fm DFF_W190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07010));
DFF_save_fm DFF_W191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07020));
DFF_save_fm DFF_W192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07100));
DFF_save_fm DFF_W193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07110));
DFF_save_fm DFF_W194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07120));
DFF_save_fm DFF_W195(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07200));
DFF_save_fm DFF_W196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07210));
DFF_save_fm DFF_W197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07220));
DFF_save_fm DFF_W198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07001));
DFF_save_fm DFF_W199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07011));
DFF_save_fm DFF_W200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07021));
DFF_save_fm DFF_W201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07101));
DFF_save_fm DFF_W202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07111));
DFF_save_fm DFF_W203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07121));
DFF_save_fm DFF_W204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07201));
DFF_save_fm DFF_W205(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07211));
DFF_save_fm DFF_W206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07221));
DFF_save_fm DFF_W207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07002));
DFF_save_fm DFF_W208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07012));
DFF_save_fm DFF_W209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07022));
DFF_save_fm DFF_W210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07102));
DFF_save_fm DFF_W211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07112));
DFF_save_fm DFF_W212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W07122));
DFF_save_fm DFF_W213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07202));
DFF_save_fm DFF_W214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07212));
DFF_save_fm DFF_W215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W07222));
DFF_save_fm DFF_W216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08000));
DFF_save_fm DFF_W217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08010));
DFF_save_fm DFF_W218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08020));
DFF_save_fm DFF_W219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08100));
DFF_save_fm DFF_W220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08110));
DFF_save_fm DFF_W221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08120));
DFF_save_fm DFF_W222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08200));
DFF_save_fm DFF_W223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08210));
DFF_save_fm DFF_W224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08220));
DFF_save_fm DFF_W225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08001));
DFF_save_fm DFF_W226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08011));
DFF_save_fm DFF_W227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08021));
DFF_save_fm DFF_W228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08101));
DFF_save_fm DFF_W229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08111));
DFF_save_fm DFF_W230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08121));
DFF_save_fm DFF_W231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08201));
DFF_save_fm DFF_W232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08211));
DFF_save_fm DFF_W233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08221));
DFF_save_fm DFF_W234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08002));
DFF_save_fm DFF_W235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08012));
DFF_save_fm DFF_W236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08022));
DFF_save_fm DFF_W237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08102));
DFF_save_fm DFF_W238(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08112));
DFF_save_fm DFF_W239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08122));
DFF_save_fm DFF_W240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08202));
DFF_save_fm DFF_W241(.clk(clk),.rstn(rstn),.reset_value(0),.q(W08212));
DFF_save_fm DFF_W242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W08222));
DFF_save_fm DFF_W243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09000));
DFF_save_fm DFF_W244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09010));
DFF_save_fm DFF_W245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09020));
DFF_save_fm DFF_W246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09100));
DFF_save_fm DFF_W247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09110));
DFF_save_fm DFF_W248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09120));
DFF_save_fm DFF_W249(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09200));
DFF_save_fm DFF_W250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09210));
DFF_save_fm DFF_W251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09220));
DFF_save_fm DFF_W252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09001));
DFF_save_fm DFF_W253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09011));
DFF_save_fm DFF_W254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09021));
DFF_save_fm DFF_W255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09101));
DFF_save_fm DFF_W256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09111));
DFF_save_fm DFF_W257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09121));
DFF_save_fm DFF_W258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09201));
DFF_save_fm DFF_W259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09211));
DFF_save_fm DFF_W260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09221));
DFF_save_fm DFF_W261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09002));
DFF_save_fm DFF_W262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09012));
DFF_save_fm DFF_W263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09022));
DFF_save_fm DFF_W264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09102));
DFF_save_fm DFF_W265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09112));
DFF_save_fm DFF_W266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09122));
DFF_save_fm DFF_W267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09202));
DFF_save_fm DFF_W268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W09212));
DFF_save_fm DFF_W269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W09222));
DFF_save_fm DFF_W270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A000));
DFF_save_fm DFF_W271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A010));
DFF_save_fm DFF_W272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A020));
DFF_save_fm DFF_W273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A100));
DFF_save_fm DFF_W274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A110));
DFF_save_fm DFF_W275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A120));
DFF_save_fm DFF_W276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A200));
DFF_save_fm DFF_W277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A210));
DFF_save_fm DFF_W278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A220));
DFF_save_fm DFF_W279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A001));
DFF_save_fm DFF_W280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A011));
DFF_save_fm DFF_W281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A021));
DFF_save_fm DFF_W282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A101));
DFF_save_fm DFF_W283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A111));
DFF_save_fm DFF_W284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A121));
DFF_save_fm DFF_W285(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A201));
DFF_save_fm DFF_W286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A211));
DFF_save_fm DFF_W287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A221));
DFF_save_fm DFF_W288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A002));
DFF_save_fm DFF_W289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A012));
DFF_save_fm DFF_W290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A022));
DFF_save_fm DFF_W291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A102));
DFF_save_fm DFF_W292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A112));
DFF_save_fm DFF_W293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A122));
DFF_save_fm DFF_W294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0A202));
DFF_save_fm DFF_W295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A212));
DFF_save_fm DFF_W296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0A222));
DFF_save_fm DFF_W297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B000));
DFF_save_fm DFF_W298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B010));
DFF_save_fm DFF_W299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B020));
DFF_save_fm DFF_W300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B100));
DFF_save_fm DFF_W301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B110));
DFF_save_fm DFF_W302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B120));
DFF_save_fm DFF_W303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B200));
DFF_save_fm DFF_W304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B210));
DFF_save_fm DFF_W305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B220));
DFF_save_fm DFF_W306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B001));
DFF_save_fm DFF_W307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B011));
DFF_save_fm DFF_W308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B021));
DFF_save_fm DFF_W309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B101));
DFF_save_fm DFF_W310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B111));
DFF_save_fm DFF_W311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B121));
DFF_save_fm DFF_W312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B201));
DFF_save_fm DFF_W313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B211));
DFF_save_fm DFF_W314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B221));
DFF_save_fm DFF_W315(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B002));
DFF_save_fm DFF_W316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B012));
DFF_save_fm DFF_W317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B022));
DFF_save_fm DFF_W318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B102));
DFF_save_fm DFF_W319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0B112));
DFF_save_fm DFF_W320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B122));
DFF_save_fm DFF_W321(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B202));
DFF_save_fm DFF_W322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B212));
DFF_save_fm DFF_W323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0B222));
DFF_save_fm DFF_W324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C000));
DFF_save_fm DFF_W325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C010));
DFF_save_fm DFF_W326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C020));
DFF_save_fm DFF_W327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C100));
DFF_save_fm DFF_W328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C110));
DFF_save_fm DFF_W329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C120));
DFF_save_fm DFF_W330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C200));
DFF_save_fm DFF_W331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C210));
DFF_save_fm DFF_W332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C220));
DFF_save_fm DFF_W333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C001));
DFF_save_fm DFF_W334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C011));
DFF_save_fm DFF_W335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C021));
DFF_save_fm DFF_W336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C101));
DFF_save_fm DFF_W337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C111));
DFF_save_fm DFF_W338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C121));
DFF_save_fm DFF_W339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C201));
DFF_save_fm DFF_W340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C211));
DFF_save_fm DFF_W341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C221));
DFF_save_fm DFF_W342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C002));
DFF_save_fm DFF_W343(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C012));
DFF_save_fm DFF_W344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C022));
DFF_save_fm DFF_W345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C102));
DFF_save_fm DFF_W346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C112));
DFF_save_fm DFF_W347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C122));
DFF_save_fm DFF_W348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C202));
DFF_save_fm DFF_W349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0C212));
DFF_save_fm DFF_W350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0C222));
DFF_save_fm DFF_W351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D000));
DFF_save_fm DFF_W352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D010));
DFF_save_fm DFF_W353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D020));
DFF_save_fm DFF_W354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D100));
DFF_save_fm DFF_W355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D110));
DFF_save_fm DFF_W356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D120));
DFF_save_fm DFF_W357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D200));
DFF_save_fm DFF_W358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D210));
DFF_save_fm DFF_W359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D220));
DFF_save_fm DFF_W360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D001));
DFF_save_fm DFF_W361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D011));
DFF_save_fm DFF_W362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D021));
DFF_save_fm DFF_W363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D101));
DFF_save_fm DFF_W364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D111));
DFF_save_fm DFF_W365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D121));
DFF_save_fm DFF_W366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D201));
DFF_save_fm DFF_W367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D211));
DFF_save_fm DFF_W368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D221));
DFF_save_fm DFF_W369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D002));
DFF_save_fm DFF_W370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D012));
DFF_save_fm DFF_W371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D022));
DFF_save_fm DFF_W372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D102));
DFF_save_fm DFF_W373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D112));
DFF_save_fm DFF_W374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D122));
DFF_save_fm DFF_W375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D202));
DFF_save_fm DFF_W376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0D212));
DFF_save_fm DFF_W377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0D222));
DFF_save_fm DFF_W378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E000));
DFF_save_fm DFF_W379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E010));
DFF_save_fm DFF_W380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E020));
DFF_save_fm DFF_W381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E100));
DFF_save_fm DFF_W382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E110));
DFF_save_fm DFF_W383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E120));
DFF_save_fm DFF_W384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E200));
DFF_save_fm DFF_W385(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E210));
DFF_save_fm DFF_W386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E220));
DFF_save_fm DFF_W387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E001));
DFF_save_fm DFF_W388(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E011));
DFF_save_fm DFF_W389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E021));
DFF_save_fm DFF_W390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E101));
DFF_save_fm DFF_W391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E111));
DFF_save_fm DFF_W392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E121));
DFF_save_fm DFF_W393(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E201));
DFF_save_fm DFF_W394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E211));
DFF_save_fm DFF_W395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E221));
DFF_save_fm DFF_W396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E002));
DFF_save_fm DFF_W397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E012));
DFF_save_fm DFF_W398(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E022));
DFF_save_fm DFF_W399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E102));
DFF_save_fm DFF_W400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E112));
DFF_save_fm DFF_W401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E122));
DFF_save_fm DFF_W402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0E202));
DFF_save_fm DFF_W403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E212));
DFF_save_fm DFF_W404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0E222));
DFF_save_fm DFF_W405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F000));
DFF_save_fm DFF_W406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F010));
DFF_save_fm DFF_W407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F020));
DFF_save_fm DFF_W408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F100));
DFF_save_fm DFF_W409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F110));
DFF_save_fm DFF_W410(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F120));
DFF_save_fm DFF_W411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F200));
DFF_save_fm DFF_W412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F210));
DFF_save_fm DFF_W413(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F220));
DFF_save_fm DFF_W414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F001));
DFF_save_fm DFF_W415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F011));
DFF_save_fm DFF_W416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F021));
DFF_save_fm DFF_W417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F101));
DFF_save_fm DFF_W418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F111));
DFF_save_fm DFF_W419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F121));
DFF_save_fm DFF_W420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F201));
DFF_save_fm DFF_W421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F211));
DFF_save_fm DFF_W422(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F221));
DFF_save_fm DFF_W423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F002));
DFF_save_fm DFF_W424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F012));
DFF_save_fm DFF_W425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F022));
DFF_save_fm DFF_W426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F102));
DFF_save_fm DFF_W427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F112));
DFF_save_fm DFF_W428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W0F122));
DFF_save_fm DFF_W429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F202));
DFF_save_fm DFF_W430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F212));
DFF_save_fm DFF_W431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W0F222));
ninexnine_unit ninexnine_unit_0(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00000)
);

ninexnine_unit ninexnine_unit_1(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01000)
);

ninexnine_unit ninexnine_unit_2(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02000)
);

assign C0000=c00000+c01000+c02000;
assign A0000=(C0000>=0)?1:0;

assign P1000=A0000;

ninexnine_unit ninexnine_unit_3(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00010)
);

ninexnine_unit ninexnine_unit_4(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01010)
);

ninexnine_unit ninexnine_unit_5(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02010)
);

assign C0010=c00010+c01010+c02010;
assign A0010=(C0010>=0)?1:0;

assign P1010=A0010;

ninexnine_unit ninexnine_unit_6(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00020)
);

ninexnine_unit ninexnine_unit_7(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01020)
);

ninexnine_unit ninexnine_unit_8(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02020)
);

assign C0020=c00020+c01020+c02020;
assign A0020=(C0020>=0)?1:0;

assign P1020=A0020;

ninexnine_unit ninexnine_unit_9(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00030)
);

ninexnine_unit ninexnine_unit_10(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01030)
);

ninexnine_unit ninexnine_unit_11(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02030)
);

assign C0030=c00030+c01030+c02030;
assign A0030=(C0030>=0)?1:0;

assign P1030=A0030;

ninexnine_unit ninexnine_unit_12(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00040)
);

ninexnine_unit ninexnine_unit_13(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01040)
);

ninexnine_unit ninexnine_unit_14(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02040)
);

assign C0040=c00040+c01040+c02040;
assign A0040=(C0040>=0)?1:0;

assign P1040=A0040;

ninexnine_unit ninexnine_unit_15(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00100)
);

ninexnine_unit ninexnine_unit_16(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01100)
);

ninexnine_unit ninexnine_unit_17(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02100)
);

assign C0100=c00100+c01100+c02100;
assign A0100=(C0100>=0)?1:0;

assign P1100=A0100;

ninexnine_unit ninexnine_unit_18(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00110)
);

ninexnine_unit ninexnine_unit_19(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01110)
);

ninexnine_unit ninexnine_unit_20(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02110)
);

assign C0110=c00110+c01110+c02110;
assign A0110=(C0110>=0)?1:0;

assign P1110=A0110;

ninexnine_unit ninexnine_unit_21(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00120)
);

ninexnine_unit ninexnine_unit_22(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01120)
);

ninexnine_unit ninexnine_unit_23(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02120)
);

assign C0120=c00120+c01120+c02120;
assign A0120=(C0120>=0)?1:0;

assign P1120=A0120;

ninexnine_unit ninexnine_unit_24(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00130)
);

ninexnine_unit ninexnine_unit_25(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01130)
);

ninexnine_unit ninexnine_unit_26(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02130)
);

assign C0130=c00130+c01130+c02130;
assign A0130=(C0130>=0)?1:0;

assign P1130=A0130;

ninexnine_unit ninexnine_unit_27(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00140)
);

ninexnine_unit ninexnine_unit_28(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01140)
);

ninexnine_unit ninexnine_unit_29(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02140)
);

assign C0140=c00140+c01140+c02140;
assign A0140=(C0140>=0)?1:0;

assign P1140=A0140;

ninexnine_unit ninexnine_unit_30(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00200)
);

ninexnine_unit ninexnine_unit_31(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01200)
);

ninexnine_unit ninexnine_unit_32(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02200)
);

assign C0200=c00200+c01200+c02200;
assign A0200=(C0200>=0)?1:0;

assign P1200=A0200;

ninexnine_unit ninexnine_unit_33(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00210)
);

ninexnine_unit ninexnine_unit_34(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01210)
);

ninexnine_unit ninexnine_unit_35(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02210)
);

assign C0210=c00210+c01210+c02210;
assign A0210=(C0210>=0)?1:0;

assign P1210=A0210;

ninexnine_unit ninexnine_unit_36(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00220)
);

ninexnine_unit ninexnine_unit_37(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01220)
);

ninexnine_unit ninexnine_unit_38(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02220)
);

assign C0220=c00220+c01220+c02220;
assign A0220=(C0220>=0)?1:0;

assign P1220=A0220;

ninexnine_unit ninexnine_unit_39(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00230)
);

ninexnine_unit ninexnine_unit_40(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01230)
);

ninexnine_unit ninexnine_unit_41(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02230)
);

assign C0230=c00230+c01230+c02230;
assign A0230=(C0230>=0)?1:0;

assign P1230=A0230;

ninexnine_unit ninexnine_unit_42(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00240)
);

ninexnine_unit ninexnine_unit_43(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01240)
);

ninexnine_unit ninexnine_unit_44(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02240)
);

assign C0240=c00240+c01240+c02240;
assign A0240=(C0240>=0)?1:0;

assign P1240=A0240;

ninexnine_unit ninexnine_unit_45(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00300)
);

ninexnine_unit ninexnine_unit_46(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01300)
);

ninexnine_unit ninexnine_unit_47(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02300)
);

assign C0300=c00300+c01300+c02300;
assign A0300=(C0300>=0)?1:0;

assign P1300=A0300;

ninexnine_unit ninexnine_unit_48(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00310)
);

ninexnine_unit ninexnine_unit_49(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01310)
);

ninexnine_unit ninexnine_unit_50(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02310)
);

assign C0310=c00310+c01310+c02310;
assign A0310=(C0310>=0)?1:0;

assign P1310=A0310;

ninexnine_unit ninexnine_unit_51(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00320)
);

ninexnine_unit ninexnine_unit_52(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01320)
);

ninexnine_unit ninexnine_unit_53(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02320)
);

assign C0320=c00320+c01320+c02320;
assign A0320=(C0320>=0)?1:0;

assign P1320=A0320;

ninexnine_unit ninexnine_unit_54(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00330)
);

ninexnine_unit ninexnine_unit_55(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01330)
);

ninexnine_unit ninexnine_unit_56(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02330)
);

assign C0330=c00330+c01330+c02330;
assign A0330=(C0330>=0)?1:0;

assign P1330=A0330;

ninexnine_unit ninexnine_unit_57(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00340)
);

ninexnine_unit ninexnine_unit_58(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01340)
);

ninexnine_unit ninexnine_unit_59(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02340)
);

assign C0340=c00340+c01340+c02340;
assign A0340=(C0340>=0)?1:0;

assign P1340=A0340;

ninexnine_unit ninexnine_unit_60(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00400)
);

ninexnine_unit ninexnine_unit_61(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01400)
);

ninexnine_unit ninexnine_unit_62(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02400)
);

assign C0400=c00400+c01400+c02400;
assign A0400=(C0400>=0)?1:0;

assign P1400=A0400;

ninexnine_unit ninexnine_unit_63(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00410)
);

ninexnine_unit ninexnine_unit_64(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01410)
);

ninexnine_unit ninexnine_unit_65(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02410)
);

assign C0410=c00410+c01410+c02410;
assign A0410=(C0410>=0)?1:0;

assign P1410=A0410;

ninexnine_unit ninexnine_unit_66(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00420)
);

ninexnine_unit ninexnine_unit_67(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01420)
);

ninexnine_unit ninexnine_unit_68(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02420)
);

assign C0420=c00420+c01420+c02420;
assign A0420=(C0420>=0)?1:0;

assign P1420=A0420;

ninexnine_unit ninexnine_unit_69(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00430)
);

ninexnine_unit ninexnine_unit_70(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01430)
);

ninexnine_unit ninexnine_unit_71(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02430)
);

assign C0430=c00430+c01430+c02430;
assign A0430=(C0430>=0)?1:0;

assign P1430=A0430;

ninexnine_unit ninexnine_unit_72(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00440)
);

ninexnine_unit ninexnine_unit_73(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01440)
);

ninexnine_unit ninexnine_unit_74(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02440)
);

assign C0440=c00440+c01440+c02440;
assign A0440=(C0440>=0)?1:0;

assign P1440=A0440;

ninexnine_unit ninexnine_unit_75(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00001)
);

ninexnine_unit ninexnine_unit_76(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01001)
);

ninexnine_unit ninexnine_unit_77(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02001)
);

assign C0001=c00001+c01001+c02001;
assign A0001=(C0001>=0)?1:0;

assign P1001=A0001;

ninexnine_unit ninexnine_unit_78(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00011)
);

ninexnine_unit ninexnine_unit_79(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01011)
);

ninexnine_unit ninexnine_unit_80(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02011)
);

assign C0011=c00011+c01011+c02011;
assign A0011=(C0011>=0)?1:0;

assign P1011=A0011;

ninexnine_unit ninexnine_unit_81(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00021)
);

ninexnine_unit ninexnine_unit_82(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01021)
);

ninexnine_unit ninexnine_unit_83(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02021)
);

assign C0021=c00021+c01021+c02021;
assign A0021=(C0021>=0)?1:0;

assign P1021=A0021;

ninexnine_unit ninexnine_unit_84(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00031)
);

ninexnine_unit ninexnine_unit_85(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01031)
);

ninexnine_unit ninexnine_unit_86(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02031)
);

assign C0031=c00031+c01031+c02031;
assign A0031=(C0031>=0)?1:0;

assign P1031=A0031;

ninexnine_unit ninexnine_unit_87(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00041)
);

ninexnine_unit ninexnine_unit_88(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01041)
);

ninexnine_unit ninexnine_unit_89(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02041)
);

assign C0041=c00041+c01041+c02041;
assign A0041=(C0041>=0)?1:0;

assign P1041=A0041;

ninexnine_unit ninexnine_unit_90(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00101)
);

ninexnine_unit ninexnine_unit_91(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01101)
);

ninexnine_unit ninexnine_unit_92(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02101)
);

assign C0101=c00101+c01101+c02101;
assign A0101=(C0101>=0)?1:0;

assign P1101=A0101;

ninexnine_unit ninexnine_unit_93(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00111)
);

ninexnine_unit ninexnine_unit_94(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01111)
);

ninexnine_unit ninexnine_unit_95(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02111)
);

assign C0111=c00111+c01111+c02111;
assign A0111=(C0111>=0)?1:0;

assign P1111=A0111;

ninexnine_unit ninexnine_unit_96(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00121)
);

ninexnine_unit ninexnine_unit_97(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01121)
);

ninexnine_unit ninexnine_unit_98(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02121)
);

assign C0121=c00121+c01121+c02121;
assign A0121=(C0121>=0)?1:0;

assign P1121=A0121;

ninexnine_unit ninexnine_unit_99(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00131)
);

ninexnine_unit ninexnine_unit_100(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01131)
);

ninexnine_unit ninexnine_unit_101(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02131)
);

assign C0131=c00131+c01131+c02131;
assign A0131=(C0131>=0)?1:0;

assign P1131=A0131;

ninexnine_unit ninexnine_unit_102(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00141)
);

ninexnine_unit ninexnine_unit_103(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01141)
);

ninexnine_unit ninexnine_unit_104(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02141)
);

assign C0141=c00141+c01141+c02141;
assign A0141=(C0141>=0)?1:0;

assign P1141=A0141;

ninexnine_unit ninexnine_unit_105(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00201)
);

ninexnine_unit ninexnine_unit_106(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01201)
);

ninexnine_unit ninexnine_unit_107(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02201)
);

assign C0201=c00201+c01201+c02201;
assign A0201=(C0201>=0)?1:0;

assign P1201=A0201;

ninexnine_unit ninexnine_unit_108(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00211)
);

ninexnine_unit ninexnine_unit_109(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01211)
);

ninexnine_unit ninexnine_unit_110(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02211)
);

assign C0211=c00211+c01211+c02211;
assign A0211=(C0211>=0)?1:0;

assign P1211=A0211;

ninexnine_unit ninexnine_unit_111(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00221)
);

ninexnine_unit ninexnine_unit_112(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01221)
);

ninexnine_unit ninexnine_unit_113(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02221)
);

assign C0221=c00221+c01221+c02221;
assign A0221=(C0221>=0)?1:0;

assign P1221=A0221;

ninexnine_unit ninexnine_unit_114(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00231)
);

ninexnine_unit ninexnine_unit_115(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01231)
);

ninexnine_unit ninexnine_unit_116(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02231)
);

assign C0231=c00231+c01231+c02231;
assign A0231=(C0231>=0)?1:0;

assign P1231=A0231;

ninexnine_unit ninexnine_unit_117(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00241)
);

ninexnine_unit ninexnine_unit_118(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01241)
);

ninexnine_unit ninexnine_unit_119(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02241)
);

assign C0241=c00241+c01241+c02241;
assign A0241=(C0241>=0)?1:0;

assign P1241=A0241;

ninexnine_unit ninexnine_unit_120(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00301)
);

ninexnine_unit ninexnine_unit_121(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01301)
);

ninexnine_unit ninexnine_unit_122(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02301)
);

assign C0301=c00301+c01301+c02301;
assign A0301=(C0301>=0)?1:0;

assign P1301=A0301;

ninexnine_unit ninexnine_unit_123(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00311)
);

ninexnine_unit ninexnine_unit_124(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01311)
);

ninexnine_unit ninexnine_unit_125(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02311)
);

assign C0311=c00311+c01311+c02311;
assign A0311=(C0311>=0)?1:0;

assign P1311=A0311;

ninexnine_unit ninexnine_unit_126(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00321)
);

ninexnine_unit ninexnine_unit_127(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01321)
);

ninexnine_unit ninexnine_unit_128(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02321)
);

assign C0321=c00321+c01321+c02321;
assign A0321=(C0321>=0)?1:0;

assign P1321=A0321;

ninexnine_unit ninexnine_unit_129(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00331)
);

ninexnine_unit ninexnine_unit_130(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01331)
);

ninexnine_unit ninexnine_unit_131(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02331)
);

assign C0331=c00331+c01331+c02331;
assign A0331=(C0331>=0)?1:0;

assign P1331=A0331;

ninexnine_unit ninexnine_unit_132(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00341)
);

ninexnine_unit ninexnine_unit_133(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01341)
);

ninexnine_unit ninexnine_unit_134(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02341)
);

assign C0341=c00341+c01341+c02341;
assign A0341=(C0341>=0)?1:0;

assign P1341=A0341;

ninexnine_unit ninexnine_unit_135(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00401)
);

ninexnine_unit ninexnine_unit_136(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01401)
);

ninexnine_unit ninexnine_unit_137(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02401)
);

assign C0401=c00401+c01401+c02401;
assign A0401=(C0401>=0)?1:0;

assign P1401=A0401;

ninexnine_unit ninexnine_unit_138(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00411)
);

ninexnine_unit ninexnine_unit_139(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01411)
);

ninexnine_unit ninexnine_unit_140(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02411)
);

assign C0411=c00411+c01411+c02411;
assign A0411=(C0411>=0)?1:0;

assign P1411=A0411;

ninexnine_unit ninexnine_unit_141(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00421)
);

ninexnine_unit ninexnine_unit_142(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01421)
);

ninexnine_unit ninexnine_unit_143(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02421)
);

assign C0421=c00421+c01421+c02421;
assign A0421=(C0421>=0)?1:0;

assign P1421=A0421;

ninexnine_unit ninexnine_unit_144(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00431)
);

ninexnine_unit ninexnine_unit_145(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01431)
);

ninexnine_unit ninexnine_unit_146(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02431)
);

assign C0431=c00431+c01431+c02431;
assign A0431=(C0431>=0)?1:0;

assign P1431=A0431;

ninexnine_unit ninexnine_unit_147(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00441)
);

ninexnine_unit ninexnine_unit_148(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01441)
);

ninexnine_unit ninexnine_unit_149(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02441)
);

assign C0441=c00441+c01441+c02441;
assign A0441=(C0441>=0)?1:0;

assign P1441=A0441;

ninexnine_unit ninexnine_unit_150(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00002)
);

ninexnine_unit ninexnine_unit_151(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01002)
);

ninexnine_unit ninexnine_unit_152(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02002)
);

assign C0002=c00002+c01002+c02002;
assign A0002=(C0002>=0)?1:0;

assign P1002=A0002;

ninexnine_unit ninexnine_unit_153(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00012)
);

ninexnine_unit ninexnine_unit_154(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01012)
);

ninexnine_unit ninexnine_unit_155(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02012)
);

assign C0012=c00012+c01012+c02012;
assign A0012=(C0012>=0)?1:0;

assign P1012=A0012;

ninexnine_unit ninexnine_unit_156(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00022)
);

ninexnine_unit ninexnine_unit_157(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01022)
);

ninexnine_unit ninexnine_unit_158(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02022)
);

assign C0022=c00022+c01022+c02022;
assign A0022=(C0022>=0)?1:0;

assign P1022=A0022;

ninexnine_unit ninexnine_unit_159(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00032)
);

ninexnine_unit ninexnine_unit_160(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01032)
);

ninexnine_unit ninexnine_unit_161(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02032)
);

assign C0032=c00032+c01032+c02032;
assign A0032=(C0032>=0)?1:0;

assign P1032=A0032;

ninexnine_unit ninexnine_unit_162(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00042)
);

ninexnine_unit ninexnine_unit_163(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01042)
);

ninexnine_unit ninexnine_unit_164(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02042)
);

assign C0042=c00042+c01042+c02042;
assign A0042=(C0042>=0)?1:0;

assign P1042=A0042;

ninexnine_unit ninexnine_unit_165(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00102)
);

ninexnine_unit ninexnine_unit_166(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01102)
);

ninexnine_unit ninexnine_unit_167(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02102)
);

assign C0102=c00102+c01102+c02102;
assign A0102=(C0102>=0)?1:0;

assign P1102=A0102;

ninexnine_unit ninexnine_unit_168(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00112)
);

ninexnine_unit ninexnine_unit_169(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01112)
);

ninexnine_unit ninexnine_unit_170(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02112)
);

assign C0112=c00112+c01112+c02112;
assign A0112=(C0112>=0)?1:0;

assign P1112=A0112;

ninexnine_unit ninexnine_unit_171(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00122)
);

ninexnine_unit ninexnine_unit_172(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01122)
);

ninexnine_unit ninexnine_unit_173(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02122)
);

assign C0122=c00122+c01122+c02122;
assign A0122=(C0122>=0)?1:0;

assign P1122=A0122;

ninexnine_unit ninexnine_unit_174(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00132)
);

ninexnine_unit ninexnine_unit_175(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01132)
);

ninexnine_unit ninexnine_unit_176(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02132)
);

assign C0132=c00132+c01132+c02132;
assign A0132=(C0132>=0)?1:0;

assign P1132=A0132;

ninexnine_unit ninexnine_unit_177(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00142)
);

ninexnine_unit ninexnine_unit_178(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01142)
);

ninexnine_unit ninexnine_unit_179(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02142)
);

assign C0142=c00142+c01142+c02142;
assign A0142=(C0142>=0)?1:0;

assign P1142=A0142;

ninexnine_unit ninexnine_unit_180(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00202)
);

ninexnine_unit ninexnine_unit_181(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01202)
);

ninexnine_unit ninexnine_unit_182(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02202)
);

assign C0202=c00202+c01202+c02202;
assign A0202=(C0202>=0)?1:0;

assign P1202=A0202;

ninexnine_unit ninexnine_unit_183(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00212)
);

ninexnine_unit ninexnine_unit_184(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01212)
);

ninexnine_unit ninexnine_unit_185(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02212)
);

assign C0212=c00212+c01212+c02212;
assign A0212=(C0212>=0)?1:0;

assign P1212=A0212;

ninexnine_unit ninexnine_unit_186(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00222)
);

ninexnine_unit ninexnine_unit_187(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01222)
);

ninexnine_unit ninexnine_unit_188(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02222)
);

assign C0222=c00222+c01222+c02222;
assign A0222=(C0222>=0)?1:0;

assign P1222=A0222;

ninexnine_unit ninexnine_unit_189(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00232)
);

ninexnine_unit ninexnine_unit_190(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01232)
);

ninexnine_unit ninexnine_unit_191(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02232)
);

assign C0232=c00232+c01232+c02232;
assign A0232=(C0232>=0)?1:0;

assign P1232=A0232;

ninexnine_unit ninexnine_unit_192(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00242)
);

ninexnine_unit ninexnine_unit_193(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01242)
);

ninexnine_unit ninexnine_unit_194(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02242)
);

assign C0242=c00242+c01242+c02242;
assign A0242=(C0242>=0)?1:0;

assign P1242=A0242;

ninexnine_unit ninexnine_unit_195(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00302)
);

ninexnine_unit ninexnine_unit_196(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01302)
);

ninexnine_unit ninexnine_unit_197(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02302)
);

assign C0302=c00302+c01302+c02302;
assign A0302=(C0302>=0)?1:0;

assign P1302=A0302;

ninexnine_unit ninexnine_unit_198(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00312)
);

ninexnine_unit ninexnine_unit_199(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01312)
);

ninexnine_unit ninexnine_unit_200(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02312)
);

assign C0312=c00312+c01312+c02312;
assign A0312=(C0312>=0)?1:0;

assign P1312=A0312;

ninexnine_unit ninexnine_unit_201(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00322)
);

ninexnine_unit ninexnine_unit_202(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01322)
);

ninexnine_unit ninexnine_unit_203(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02322)
);

assign C0322=c00322+c01322+c02322;
assign A0322=(C0322>=0)?1:0;

assign P1322=A0322;

ninexnine_unit ninexnine_unit_204(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00332)
);

ninexnine_unit ninexnine_unit_205(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01332)
);

ninexnine_unit ninexnine_unit_206(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02332)
);

assign C0332=c00332+c01332+c02332;
assign A0332=(C0332>=0)?1:0;

assign P1332=A0332;

ninexnine_unit ninexnine_unit_207(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00342)
);

ninexnine_unit ninexnine_unit_208(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01342)
);

ninexnine_unit ninexnine_unit_209(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02342)
);

assign C0342=c00342+c01342+c02342;
assign A0342=(C0342>=0)?1:0;

assign P1342=A0342;

ninexnine_unit ninexnine_unit_210(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00402)
);

ninexnine_unit ninexnine_unit_211(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01402)
);

ninexnine_unit ninexnine_unit_212(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02402)
);

assign C0402=c00402+c01402+c02402;
assign A0402=(C0402>=0)?1:0;

assign P1402=A0402;

ninexnine_unit ninexnine_unit_213(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00412)
);

ninexnine_unit ninexnine_unit_214(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01412)
);

ninexnine_unit ninexnine_unit_215(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02412)
);

assign C0412=c00412+c01412+c02412;
assign A0412=(C0412>=0)?1:0;

assign P1412=A0412;

ninexnine_unit ninexnine_unit_216(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00422)
);

ninexnine_unit ninexnine_unit_217(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01422)
);

ninexnine_unit ninexnine_unit_218(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02422)
);

assign C0422=c00422+c01422+c02422;
assign A0422=(C0422>=0)?1:0;

assign P1422=A0422;

ninexnine_unit ninexnine_unit_219(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00432)
);

ninexnine_unit ninexnine_unit_220(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01432)
);

ninexnine_unit ninexnine_unit_221(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02432)
);

assign C0432=c00432+c01432+c02432;
assign A0432=(C0432>=0)?1:0;

assign P1432=A0432;

ninexnine_unit ninexnine_unit_222(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00442)
);

ninexnine_unit ninexnine_unit_223(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01442)
);

ninexnine_unit ninexnine_unit_224(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02442)
);

assign C0442=c00442+c01442+c02442;
assign A0442=(C0442>=0)?1:0;

assign P1442=A0442;

ninexnine_unit ninexnine_unit_225(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00003)
);

ninexnine_unit ninexnine_unit_226(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01003)
);

ninexnine_unit ninexnine_unit_227(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02003)
);

assign C0003=c00003+c01003+c02003;
assign A0003=(C0003>=0)?1:0;

assign P1003=A0003;

ninexnine_unit ninexnine_unit_228(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00013)
);

ninexnine_unit ninexnine_unit_229(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01013)
);

ninexnine_unit ninexnine_unit_230(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02013)
);

assign C0013=c00013+c01013+c02013;
assign A0013=(C0013>=0)?1:0;

assign P1013=A0013;

ninexnine_unit ninexnine_unit_231(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00023)
);

ninexnine_unit ninexnine_unit_232(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01023)
);

ninexnine_unit ninexnine_unit_233(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02023)
);

assign C0023=c00023+c01023+c02023;
assign A0023=(C0023>=0)?1:0;

assign P1023=A0023;

ninexnine_unit ninexnine_unit_234(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00033)
);

ninexnine_unit ninexnine_unit_235(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01033)
);

ninexnine_unit ninexnine_unit_236(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02033)
);

assign C0033=c00033+c01033+c02033;
assign A0033=(C0033>=0)?1:0;

assign P1033=A0033;

ninexnine_unit ninexnine_unit_237(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00043)
);

ninexnine_unit ninexnine_unit_238(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01043)
);

ninexnine_unit ninexnine_unit_239(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02043)
);

assign C0043=c00043+c01043+c02043;
assign A0043=(C0043>=0)?1:0;

assign P1043=A0043;

ninexnine_unit ninexnine_unit_240(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00103)
);

ninexnine_unit ninexnine_unit_241(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01103)
);

ninexnine_unit ninexnine_unit_242(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02103)
);

assign C0103=c00103+c01103+c02103;
assign A0103=(C0103>=0)?1:0;

assign P1103=A0103;

ninexnine_unit ninexnine_unit_243(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00113)
);

ninexnine_unit ninexnine_unit_244(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01113)
);

ninexnine_unit ninexnine_unit_245(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02113)
);

assign C0113=c00113+c01113+c02113;
assign A0113=(C0113>=0)?1:0;

assign P1113=A0113;

ninexnine_unit ninexnine_unit_246(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00123)
);

ninexnine_unit ninexnine_unit_247(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01123)
);

ninexnine_unit ninexnine_unit_248(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02123)
);

assign C0123=c00123+c01123+c02123;
assign A0123=(C0123>=0)?1:0;

assign P1123=A0123;

ninexnine_unit ninexnine_unit_249(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00133)
);

ninexnine_unit ninexnine_unit_250(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01133)
);

ninexnine_unit ninexnine_unit_251(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02133)
);

assign C0133=c00133+c01133+c02133;
assign A0133=(C0133>=0)?1:0;

assign P1133=A0133;

ninexnine_unit ninexnine_unit_252(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00143)
);

ninexnine_unit ninexnine_unit_253(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01143)
);

ninexnine_unit ninexnine_unit_254(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02143)
);

assign C0143=c00143+c01143+c02143;
assign A0143=(C0143>=0)?1:0;

assign P1143=A0143;

ninexnine_unit ninexnine_unit_255(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00203)
);

ninexnine_unit ninexnine_unit_256(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01203)
);

ninexnine_unit ninexnine_unit_257(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02203)
);

assign C0203=c00203+c01203+c02203;
assign A0203=(C0203>=0)?1:0;

assign P1203=A0203;

ninexnine_unit ninexnine_unit_258(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00213)
);

ninexnine_unit ninexnine_unit_259(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01213)
);

ninexnine_unit ninexnine_unit_260(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02213)
);

assign C0213=c00213+c01213+c02213;
assign A0213=(C0213>=0)?1:0;

assign P1213=A0213;

ninexnine_unit ninexnine_unit_261(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00223)
);

ninexnine_unit ninexnine_unit_262(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01223)
);

ninexnine_unit ninexnine_unit_263(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02223)
);

assign C0223=c00223+c01223+c02223;
assign A0223=(C0223>=0)?1:0;

assign P1223=A0223;

ninexnine_unit ninexnine_unit_264(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00233)
);

ninexnine_unit ninexnine_unit_265(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01233)
);

ninexnine_unit ninexnine_unit_266(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02233)
);

assign C0233=c00233+c01233+c02233;
assign A0233=(C0233>=0)?1:0;

assign P1233=A0233;

ninexnine_unit ninexnine_unit_267(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00243)
);

ninexnine_unit ninexnine_unit_268(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01243)
);

ninexnine_unit ninexnine_unit_269(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02243)
);

assign C0243=c00243+c01243+c02243;
assign A0243=(C0243>=0)?1:0;

assign P1243=A0243;

ninexnine_unit ninexnine_unit_270(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00303)
);

ninexnine_unit ninexnine_unit_271(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01303)
);

ninexnine_unit ninexnine_unit_272(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02303)
);

assign C0303=c00303+c01303+c02303;
assign A0303=(C0303>=0)?1:0;

assign P1303=A0303;

ninexnine_unit ninexnine_unit_273(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00313)
);

ninexnine_unit ninexnine_unit_274(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01313)
);

ninexnine_unit ninexnine_unit_275(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02313)
);

assign C0313=c00313+c01313+c02313;
assign A0313=(C0313>=0)?1:0;

assign P1313=A0313;

ninexnine_unit ninexnine_unit_276(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00323)
);

ninexnine_unit ninexnine_unit_277(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01323)
);

ninexnine_unit ninexnine_unit_278(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02323)
);

assign C0323=c00323+c01323+c02323;
assign A0323=(C0323>=0)?1:0;

assign P1323=A0323;

ninexnine_unit ninexnine_unit_279(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00333)
);

ninexnine_unit ninexnine_unit_280(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01333)
);

ninexnine_unit ninexnine_unit_281(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02333)
);

assign C0333=c00333+c01333+c02333;
assign A0333=(C0333>=0)?1:0;

assign P1333=A0333;

ninexnine_unit ninexnine_unit_282(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00343)
);

ninexnine_unit ninexnine_unit_283(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01343)
);

ninexnine_unit ninexnine_unit_284(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02343)
);

assign C0343=c00343+c01343+c02343;
assign A0343=(C0343>=0)?1:0;

assign P1343=A0343;

ninexnine_unit ninexnine_unit_285(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00403)
);

ninexnine_unit ninexnine_unit_286(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01403)
);

ninexnine_unit ninexnine_unit_287(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02403)
);

assign C0403=c00403+c01403+c02403;
assign A0403=(C0403>=0)?1:0;

assign P1403=A0403;

ninexnine_unit ninexnine_unit_288(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00413)
);

ninexnine_unit ninexnine_unit_289(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01413)
);

ninexnine_unit ninexnine_unit_290(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02413)
);

assign C0413=c00413+c01413+c02413;
assign A0413=(C0413>=0)?1:0;

assign P1413=A0413;

ninexnine_unit ninexnine_unit_291(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00423)
);

ninexnine_unit ninexnine_unit_292(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01423)
);

ninexnine_unit ninexnine_unit_293(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02423)
);

assign C0423=c00423+c01423+c02423;
assign A0423=(C0423>=0)?1:0;

assign P1423=A0423;

ninexnine_unit ninexnine_unit_294(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00433)
);

ninexnine_unit ninexnine_unit_295(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01433)
);

ninexnine_unit ninexnine_unit_296(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02433)
);

assign C0433=c00433+c01433+c02433;
assign A0433=(C0433>=0)?1:0;

assign P1433=A0433;

ninexnine_unit ninexnine_unit_297(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00443)
);

ninexnine_unit ninexnine_unit_298(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01443)
);

ninexnine_unit ninexnine_unit_299(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02443)
);

assign C0443=c00443+c01443+c02443;
assign A0443=(C0443>=0)?1:0;

assign P1443=A0443;

ninexnine_unit ninexnine_unit_300(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00004)
);

ninexnine_unit ninexnine_unit_301(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01004)
);

ninexnine_unit ninexnine_unit_302(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02004)
);

assign C0004=c00004+c01004+c02004;
assign A0004=(C0004>=0)?1:0;

assign P1004=A0004;

ninexnine_unit ninexnine_unit_303(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00014)
);

ninexnine_unit ninexnine_unit_304(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01014)
);

ninexnine_unit ninexnine_unit_305(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02014)
);

assign C0014=c00014+c01014+c02014;
assign A0014=(C0014>=0)?1:0;

assign P1014=A0014;

ninexnine_unit ninexnine_unit_306(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00024)
);

ninexnine_unit ninexnine_unit_307(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01024)
);

ninexnine_unit ninexnine_unit_308(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02024)
);

assign C0024=c00024+c01024+c02024;
assign A0024=(C0024>=0)?1:0;

assign P1024=A0024;

ninexnine_unit ninexnine_unit_309(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00034)
);

ninexnine_unit ninexnine_unit_310(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01034)
);

ninexnine_unit ninexnine_unit_311(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02034)
);

assign C0034=c00034+c01034+c02034;
assign A0034=(C0034>=0)?1:0;

assign P1034=A0034;

ninexnine_unit ninexnine_unit_312(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00044)
);

ninexnine_unit ninexnine_unit_313(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01044)
);

ninexnine_unit ninexnine_unit_314(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02044)
);

assign C0044=c00044+c01044+c02044;
assign A0044=(C0044>=0)?1:0;

assign P1044=A0044;

ninexnine_unit ninexnine_unit_315(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00104)
);

ninexnine_unit ninexnine_unit_316(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01104)
);

ninexnine_unit ninexnine_unit_317(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02104)
);

assign C0104=c00104+c01104+c02104;
assign A0104=(C0104>=0)?1:0;

assign P1104=A0104;

ninexnine_unit ninexnine_unit_318(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00114)
);

ninexnine_unit ninexnine_unit_319(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01114)
);

ninexnine_unit ninexnine_unit_320(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02114)
);

assign C0114=c00114+c01114+c02114;
assign A0114=(C0114>=0)?1:0;

assign P1114=A0114;

ninexnine_unit ninexnine_unit_321(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00124)
);

ninexnine_unit ninexnine_unit_322(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01124)
);

ninexnine_unit ninexnine_unit_323(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02124)
);

assign C0124=c00124+c01124+c02124;
assign A0124=(C0124>=0)?1:0;

assign P1124=A0124;

ninexnine_unit ninexnine_unit_324(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00134)
);

ninexnine_unit ninexnine_unit_325(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01134)
);

ninexnine_unit ninexnine_unit_326(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02134)
);

assign C0134=c00134+c01134+c02134;
assign A0134=(C0134>=0)?1:0;

assign P1134=A0134;

ninexnine_unit ninexnine_unit_327(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00144)
);

ninexnine_unit ninexnine_unit_328(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01144)
);

ninexnine_unit ninexnine_unit_329(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02144)
);

assign C0144=c00144+c01144+c02144;
assign A0144=(C0144>=0)?1:0;

assign P1144=A0144;

ninexnine_unit ninexnine_unit_330(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00204)
);

ninexnine_unit ninexnine_unit_331(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01204)
);

ninexnine_unit ninexnine_unit_332(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02204)
);

assign C0204=c00204+c01204+c02204;
assign A0204=(C0204>=0)?1:0;

assign P1204=A0204;

ninexnine_unit ninexnine_unit_333(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00214)
);

ninexnine_unit ninexnine_unit_334(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01214)
);

ninexnine_unit ninexnine_unit_335(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02214)
);

assign C0214=c00214+c01214+c02214;
assign A0214=(C0214>=0)?1:0;

assign P1214=A0214;

ninexnine_unit ninexnine_unit_336(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00224)
);

ninexnine_unit ninexnine_unit_337(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01224)
);

ninexnine_unit ninexnine_unit_338(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02224)
);

assign C0224=c00224+c01224+c02224;
assign A0224=(C0224>=0)?1:0;

assign P1224=A0224;

ninexnine_unit ninexnine_unit_339(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00234)
);

ninexnine_unit ninexnine_unit_340(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01234)
);

ninexnine_unit ninexnine_unit_341(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02234)
);

assign C0234=c00234+c01234+c02234;
assign A0234=(C0234>=0)?1:0;

assign P1234=A0234;

ninexnine_unit ninexnine_unit_342(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00244)
);

ninexnine_unit ninexnine_unit_343(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01244)
);

ninexnine_unit ninexnine_unit_344(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02244)
);

assign C0244=c00244+c01244+c02244;
assign A0244=(C0244>=0)?1:0;

assign P1244=A0244;

ninexnine_unit ninexnine_unit_345(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00304)
);

ninexnine_unit ninexnine_unit_346(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01304)
);

ninexnine_unit ninexnine_unit_347(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02304)
);

assign C0304=c00304+c01304+c02304;
assign A0304=(C0304>=0)?1:0;

assign P1304=A0304;

ninexnine_unit ninexnine_unit_348(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00314)
);

ninexnine_unit ninexnine_unit_349(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01314)
);

ninexnine_unit ninexnine_unit_350(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02314)
);

assign C0314=c00314+c01314+c02314;
assign A0314=(C0314>=0)?1:0;

assign P1314=A0314;

ninexnine_unit ninexnine_unit_351(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00324)
);

ninexnine_unit ninexnine_unit_352(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01324)
);

ninexnine_unit ninexnine_unit_353(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02324)
);

assign C0324=c00324+c01324+c02324;
assign A0324=(C0324>=0)?1:0;

assign P1324=A0324;

ninexnine_unit ninexnine_unit_354(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00334)
);

ninexnine_unit ninexnine_unit_355(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01334)
);

ninexnine_unit ninexnine_unit_356(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02334)
);

assign C0334=c00334+c01334+c02334;
assign A0334=(C0334>=0)?1:0;

assign P1334=A0334;

ninexnine_unit ninexnine_unit_357(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00344)
);

ninexnine_unit ninexnine_unit_358(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01344)
);

ninexnine_unit ninexnine_unit_359(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02344)
);

assign C0344=c00344+c01344+c02344;
assign A0344=(C0344>=0)?1:0;

assign P1344=A0344;

ninexnine_unit ninexnine_unit_360(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00404)
);

ninexnine_unit ninexnine_unit_361(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01404)
);

ninexnine_unit ninexnine_unit_362(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02404)
);

assign C0404=c00404+c01404+c02404;
assign A0404=(C0404>=0)?1:0;

assign P1404=A0404;

ninexnine_unit ninexnine_unit_363(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00414)
);

ninexnine_unit ninexnine_unit_364(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01414)
);

ninexnine_unit ninexnine_unit_365(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02414)
);

assign C0414=c00414+c01414+c02414;
assign A0414=(C0414>=0)?1:0;

assign P1414=A0414;

ninexnine_unit ninexnine_unit_366(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00424)
);

ninexnine_unit ninexnine_unit_367(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01424)
);

ninexnine_unit ninexnine_unit_368(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02424)
);

assign C0424=c00424+c01424+c02424;
assign A0424=(C0424>=0)?1:0;

assign P1424=A0424;

ninexnine_unit ninexnine_unit_369(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00434)
);

ninexnine_unit ninexnine_unit_370(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01434)
);

ninexnine_unit ninexnine_unit_371(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02434)
);

assign C0434=c00434+c01434+c02434;
assign A0434=(C0434>=0)?1:0;

assign P1434=A0434;

ninexnine_unit ninexnine_unit_372(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W04000),
				.b1(W04010),
				.b2(W04020),
				.b3(W04100),
				.b4(W04110),
				.b5(W04120),
				.b6(W04200),
				.b7(W04210),
				.b8(W04220),
				.c(c00444)
);

ninexnine_unit ninexnine_unit_373(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W04001),
				.b1(W04011),
				.b2(W04021),
				.b3(W04101),
				.b4(W04111),
				.b5(W04121),
				.b6(W04201),
				.b7(W04211),
				.b8(W04221),
				.c(c01444)
);

ninexnine_unit ninexnine_unit_374(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W04002),
				.b1(W04012),
				.b2(W04022),
				.b3(W04102),
				.b4(W04112),
				.b5(W04122),
				.b6(W04202),
				.b7(W04212),
				.b8(W04222),
				.c(c02444)
);

assign C0444=c00444+c01444+c02444;
assign A0444=(C0444>=0)?1:0;

assign P1444=A0444;

ninexnine_unit ninexnine_unit_375(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00005)
);

ninexnine_unit ninexnine_unit_376(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01005)
);

ninexnine_unit ninexnine_unit_377(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02005)
);

assign C0005=c00005+c01005+c02005;
assign A0005=(C0005>=0)?1:0;

assign P1005=A0005;

ninexnine_unit ninexnine_unit_378(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00015)
);

ninexnine_unit ninexnine_unit_379(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01015)
);

ninexnine_unit ninexnine_unit_380(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02015)
);

assign C0015=c00015+c01015+c02015;
assign A0015=(C0015>=0)?1:0;

assign P1015=A0015;

ninexnine_unit ninexnine_unit_381(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00025)
);

ninexnine_unit ninexnine_unit_382(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01025)
);

ninexnine_unit ninexnine_unit_383(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02025)
);

assign C0025=c00025+c01025+c02025;
assign A0025=(C0025>=0)?1:0;

assign P1025=A0025;

ninexnine_unit ninexnine_unit_384(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00035)
);

ninexnine_unit ninexnine_unit_385(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01035)
);

ninexnine_unit ninexnine_unit_386(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02035)
);

assign C0035=c00035+c01035+c02035;
assign A0035=(C0035>=0)?1:0;

assign P1035=A0035;

ninexnine_unit ninexnine_unit_387(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00045)
);

ninexnine_unit ninexnine_unit_388(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01045)
);

ninexnine_unit ninexnine_unit_389(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02045)
);

assign C0045=c00045+c01045+c02045;
assign A0045=(C0045>=0)?1:0;

assign P1045=A0045;

ninexnine_unit ninexnine_unit_390(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00105)
);

ninexnine_unit ninexnine_unit_391(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01105)
);

ninexnine_unit ninexnine_unit_392(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02105)
);

assign C0105=c00105+c01105+c02105;
assign A0105=(C0105>=0)?1:0;

assign P1105=A0105;

ninexnine_unit ninexnine_unit_393(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00115)
);

ninexnine_unit ninexnine_unit_394(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01115)
);

ninexnine_unit ninexnine_unit_395(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02115)
);

assign C0115=c00115+c01115+c02115;
assign A0115=(C0115>=0)?1:0;

assign P1115=A0115;

ninexnine_unit ninexnine_unit_396(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00125)
);

ninexnine_unit ninexnine_unit_397(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01125)
);

ninexnine_unit ninexnine_unit_398(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02125)
);

assign C0125=c00125+c01125+c02125;
assign A0125=(C0125>=0)?1:0;

assign P1125=A0125;

ninexnine_unit ninexnine_unit_399(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00135)
);

ninexnine_unit ninexnine_unit_400(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01135)
);

ninexnine_unit ninexnine_unit_401(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02135)
);

assign C0135=c00135+c01135+c02135;
assign A0135=(C0135>=0)?1:0;

assign P1135=A0135;

ninexnine_unit ninexnine_unit_402(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00145)
);

ninexnine_unit ninexnine_unit_403(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01145)
);

ninexnine_unit ninexnine_unit_404(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02145)
);

assign C0145=c00145+c01145+c02145;
assign A0145=(C0145>=0)?1:0;

assign P1145=A0145;

ninexnine_unit ninexnine_unit_405(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00205)
);

ninexnine_unit ninexnine_unit_406(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01205)
);

ninexnine_unit ninexnine_unit_407(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02205)
);

assign C0205=c00205+c01205+c02205;
assign A0205=(C0205>=0)?1:0;

assign P1205=A0205;

ninexnine_unit ninexnine_unit_408(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00215)
);

ninexnine_unit ninexnine_unit_409(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01215)
);

ninexnine_unit ninexnine_unit_410(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02215)
);

assign C0215=c00215+c01215+c02215;
assign A0215=(C0215>=0)?1:0;

assign P1215=A0215;

ninexnine_unit ninexnine_unit_411(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00225)
);

ninexnine_unit ninexnine_unit_412(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01225)
);

ninexnine_unit ninexnine_unit_413(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02225)
);

assign C0225=c00225+c01225+c02225;
assign A0225=(C0225>=0)?1:0;

assign P1225=A0225;

ninexnine_unit ninexnine_unit_414(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00235)
);

ninexnine_unit ninexnine_unit_415(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01235)
);

ninexnine_unit ninexnine_unit_416(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02235)
);

assign C0235=c00235+c01235+c02235;
assign A0235=(C0235>=0)?1:0;

assign P1235=A0235;

ninexnine_unit ninexnine_unit_417(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00245)
);

ninexnine_unit ninexnine_unit_418(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01245)
);

ninexnine_unit ninexnine_unit_419(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02245)
);

assign C0245=c00245+c01245+c02245;
assign A0245=(C0245>=0)?1:0;

assign P1245=A0245;

ninexnine_unit ninexnine_unit_420(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00305)
);

ninexnine_unit ninexnine_unit_421(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01305)
);

ninexnine_unit ninexnine_unit_422(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02305)
);

assign C0305=c00305+c01305+c02305;
assign A0305=(C0305>=0)?1:0;

assign P1305=A0305;

ninexnine_unit ninexnine_unit_423(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00315)
);

ninexnine_unit ninexnine_unit_424(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01315)
);

ninexnine_unit ninexnine_unit_425(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02315)
);

assign C0315=c00315+c01315+c02315;
assign A0315=(C0315>=0)?1:0;

assign P1315=A0315;

ninexnine_unit ninexnine_unit_426(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00325)
);

ninexnine_unit ninexnine_unit_427(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01325)
);

ninexnine_unit ninexnine_unit_428(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02325)
);

assign C0325=c00325+c01325+c02325;
assign A0325=(C0325>=0)?1:0;

assign P1325=A0325;

ninexnine_unit ninexnine_unit_429(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00335)
);

ninexnine_unit ninexnine_unit_430(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01335)
);

ninexnine_unit ninexnine_unit_431(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02335)
);

assign C0335=c00335+c01335+c02335;
assign A0335=(C0335>=0)?1:0;

assign P1335=A0335;

ninexnine_unit ninexnine_unit_432(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00345)
);

ninexnine_unit ninexnine_unit_433(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01345)
);

ninexnine_unit ninexnine_unit_434(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02345)
);

assign C0345=c00345+c01345+c02345;
assign A0345=(C0345>=0)?1:0;

assign P1345=A0345;

ninexnine_unit ninexnine_unit_435(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00405)
);

ninexnine_unit ninexnine_unit_436(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01405)
);

ninexnine_unit ninexnine_unit_437(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02405)
);

assign C0405=c00405+c01405+c02405;
assign A0405=(C0405>=0)?1:0;

assign P1405=A0405;

ninexnine_unit ninexnine_unit_438(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00415)
);

ninexnine_unit ninexnine_unit_439(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01415)
);

ninexnine_unit ninexnine_unit_440(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02415)
);

assign C0415=c00415+c01415+c02415;
assign A0415=(C0415>=0)?1:0;

assign P1415=A0415;

ninexnine_unit ninexnine_unit_441(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00425)
);

ninexnine_unit ninexnine_unit_442(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01425)
);

ninexnine_unit ninexnine_unit_443(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02425)
);

assign C0425=c00425+c01425+c02425;
assign A0425=(C0425>=0)?1:0;

assign P1425=A0425;

ninexnine_unit ninexnine_unit_444(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00435)
);

ninexnine_unit ninexnine_unit_445(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01435)
);

ninexnine_unit ninexnine_unit_446(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02435)
);

assign C0435=c00435+c01435+c02435;
assign A0435=(C0435>=0)?1:0;

assign P1435=A0435;

ninexnine_unit ninexnine_unit_447(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W05000),
				.b1(W05010),
				.b2(W05020),
				.b3(W05100),
				.b4(W05110),
				.b5(W05120),
				.b6(W05200),
				.b7(W05210),
				.b8(W05220),
				.c(c00445)
);

ninexnine_unit ninexnine_unit_448(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W05001),
				.b1(W05011),
				.b2(W05021),
				.b3(W05101),
				.b4(W05111),
				.b5(W05121),
				.b6(W05201),
				.b7(W05211),
				.b8(W05221),
				.c(c01445)
);

ninexnine_unit ninexnine_unit_449(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W05002),
				.b1(W05012),
				.b2(W05022),
				.b3(W05102),
				.b4(W05112),
				.b5(W05122),
				.b6(W05202),
				.b7(W05212),
				.b8(W05222),
				.c(c02445)
);

assign C0445=c00445+c01445+c02445;
assign A0445=(C0445>=0)?1:0;

assign P1445=A0445;

ninexnine_unit ninexnine_unit_450(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00006)
);

ninexnine_unit ninexnine_unit_451(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01006)
);

ninexnine_unit ninexnine_unit_452(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02006)
);

assign C0006=c00006+c01006+c02006;
assign A0006=(C0006>=0)?1:0;

assign P1006=A0006;

ninexnine_unit ninexnine_unit_453(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00016)
);

ninexnine_unit ninexnine_unit_454(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01016)
);

ninexnine_unit ninexnine_unit_455(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02016)
);

assign C0016=c00016+c01016+c02016;
assign A0016=(C0016>=0)?1:0;

assign P1016=A0016;

ninexnine_unit ninexnine_unit_456(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00026)
);

ninexnine_unit ninexnine_unit_457(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01026)
);

ninexnine_unit ninexnine_unit_458(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02026)
);

assign C0026=c00026+c01026+c02026;
assign A0026=(C0026>=0)?1:0;

assign P1026=A0026;

ninexnine_unit ninexnine_unit_459(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00036)
);

ninexnine_unit ninexnine_unit_460(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01036)
);

ninexnine_unit ninexnine_unit_461(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02036)
);

assign C0036=c00036+c01036+c02036;
assign A0036=(C0036>=0)?1:0;

assign P1036=A0036;

ninexnine_unit ninexnine_unit_462(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00046)
);

ninexnine_unit ninexnine_unit_463(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01046)
);

ninexnine_unit ninexnine_unit_464(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02046)
);

assign C0046=c00046+c01046+c02046;
assign A0046=(C0046>=0)?1:0;

assign P1046=A0046;

ninexnine_unit ninexnine_unit_465(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00106)
);

ninexnine_unit ninexnine_unit_466(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01106)
);

ninexnine_unit ninexnine_unit_467(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02106)
);

assign C0106=c00106+c01106+c02106;
assign A0106=(C0106>=0)?1:0;

assign P1106=A0106;

ninexnine_unit ninexnine_unit_468(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00116)
);

ninexnine_unit ninexnine_unit_469(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01116)
);

ninexnine_unit ninexnine_unit_470(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02116)
);

assign C0116=c00116+c01116+c02116;
assign A0116=(C0116>=0)?1:0;

assign P1116=A0116;

ninexnine_unit ninexnine_unit_471(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00126)
);

ninexnine_unit ninexnine_unit_472(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01126)
);

ninexnine_unit ninexnine_unit_473(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02126)
);

assign C0126=c00126+c01126+c02126;
assign A0126=(C0126>=0)?1:0;

assign P1126=A0126;

ninexnine_unit ninexnine_unit_474(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00136)
);

ninexnine_unit ninexnine_unit_475(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01136)
);

ninexnine_unit ninexnine_unit_476(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02136)
);

assign C0136=c00136+c01136+c02136;
assign A0136=(C0136>=0)?1:0;

assign P1136=A0136;

ninexnine_unit ninexnine_unit_477(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00146)
);

ninexnine_unit ninexnine_unit_478(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01146)
);

ninexnine_unit ninexnine_unit_479(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02146)
);

assign C0146=c00146+c01146+c02146;
assign A0146=(C0146>=0)?1:0;

assign P1146=A0146;

ninexnine_unit ninexnine_unit_480(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00206)
);

ninexnine_unit ninexnine_unit_481(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01206)
);

ninexnine_unit ninexnine_unit_482(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02206)
);

assign C0206=c00206+c01206+c02206;
assign A0206=(C0206>=0)?1:0;

assign P1206=A0206;

ninexnine_unit ninexnine_unit_483(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00216)
);

ninexnine_unit ninexnine_unit_484(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01216)
);

ninexnine_unit ninexnine_unit_485(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02216)
);

assign C0216=c00216+c01216+c02216;
assign A0216=(C0216>=0)?1:0;

assign P1216=A0216;

ninexnine_unit ninexnine_unit_486(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00226)
);

ninexnine_unit ninexnine_unit_487(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01226)
);

ninexnine_unit ninexnine_unit_488(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02226)
);

assign C0226=c00226+c01226+c02226;
assign A0226=(C0226>=0)?1:0;

assign P1226=A0226;

ninexnine_unit ninexnine_unit_489(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00236)
);

ninexnine_unit ninexnine_unit_490(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01236)
);

ninexnine_unit ninexnine_unit_491(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02236)
);

assign C0236=c00236+c01236+c02236;
assign A0236=(C0236>=0)?1:0;

assign P1236=A0236;

ninexnine_unit ninexnine_unit_492(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00246)
);

ninexnine_unit ninexnine_unit_493(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01246)
);

ninexnine_unit ninexnine_unit_494(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02246)
);

assign C0246=c00246+c01246+c02246;
assign A0246=(C0246>=0)?1:0;

assign P1246=A0246;

ninexnine_unit ninexnine_unit_495(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00306)
);

ninexnine_unit ninexnine_unit_496(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01306)
);

ninexnine_unit ninexnine_unit_497(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02306)
);

assign C0306=c00306+c01306+c02306;
assign A0306=(C0306>=0)?1:0;

assign P1306=A0306;

ninexnine_unit ninexnine_unit_498(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00316)
);

ninexnine_unit ninexnine_unit_499(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01316)
);

ninexnine_unit ninexnine_unit_500(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02316)
);

assign C0316=c00316+c01316+c02316;
assign A0316=(C0316>=0)?1:0;

assign P1316=A0316;

ninexnine_unit ninexnine_unit_501(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00326)
);

ninexnine_unit ninexnine_unit_502(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01326)
);

ninexnine_unit ninexnine_unit_503(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02326)
);

assign C0326=c00326+c01326+c02326;
assign A0326=(C0326>=0)?1:0;

assign P1326=A0326;

ninexnine_unit ninexnine_unit_504(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00336)
);

ninexnine_unit ninexnine_unit_505(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01336)
);

ninexnine_unit ninexnine_unit_506(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02336)
);

assign C0336=c00336+c01336+c02336;
assign A0336=(C0336>=0)?1:0;

assign P1336=A0336;

ninexnine_unit ninexnine_unit_507(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00346)
);

ninexnine_unit ninexnine_unit_508(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01346)
);

ninexnine_unit ninexnine_unit_509(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02346)
);

assign C0346=c00346+c01346+c02346;
assign A0346=(C0346>=0)?1:0;

assign P1346=A0346;

ninexnine_unit ninexnine_unit_510(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00406)
);

ninexnine_unit ninexnine_unit_511(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01406)
);

ninexnine_unit ninexnine_unit_512(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02406)
);

assign C0406=c00406+c01406+c02406;
assign A0406=(C0406>=0)?1:0;

assign P1406=A0406;

ninexnine_unit ninexnine_unit_513(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00416)
);

ninexnine_unit ninexnine_unit_514(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01416)
);

ninexnine_unit ninexnine_unit_515(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02416)
);

assign C0416=c00416+c01416+c02416;
assign A0416=(C0416>=0)?1:0;

assign P1416=A0416;

ninexnine_unit ninexnine_unit_516(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00426)
);

ninexnine_unit ninexnine_unit_517(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01426)
);

ninexnine_unit ninexnine_unit_518(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02426)
);

assign C0426=c00426+c01426+c02426;
assign A0426=(C0426>=0)?1:0;

assign P1426=A0426;

ninexnine_unit ninexnine_unit_519(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00436)
);

ninexnine_unit ninexnine_unit_520(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01436)
);

ninexnine_unit ninexnine_unit_521(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02436)
);

assign C0436=c00436+c01436+c02436;
assign A0436=(C0436>=0)?1:0;

assign P1436=A0436;

ninexnine_unit ninexnine_unit_522(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W06000),
				.b1(W06010),
				.b2(W06020),
				.b3(W06100),
				.b4(W06110),
				.b5(W06120),
				.b6(W06200),
				.b7(W06210),
				.b8(W06220),
				.c(c00446)
);

ninexnine_unit ninexnine_unit_523(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W06001),
				.b1(W06011),
				.b2(W06021),
				.b3(W06101),
				.b4(W06111),
				.b5(W06121),
				.b6(W06201),
				.b7(W06211),
				.b8(W06221),
				.c(c01446)
);

ninexnine_unit ninexnine_unit_524(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W06002),
				.b1(W06012),
				.b2(W06022),
				.b3(W06102),
				.b4(W06112),
				.b5(W06122),
				.b6(W06202),
				.b7(W06212),
				.b8(W06222),
				.c(c02446)
);

assign C0446=c00446+c01446+c02446;
assign A0446=(C0446>=0)?1:0;

assign P1446=A0446;

ninexnine_unit ninexnine_unit_525(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00007)
);

ninexnine_unit ninexnine_unit_526(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01007)
);

ninexnine_unit ninexnine_unit_527(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02007)
);

assign C0007=c00007+c01007+c02007;
assign A0007=(C0007>=0)?1:0;

assign P1007=A0007;

ninexnine_unit ninexnine_unit_528(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00017)
);

ninexnine_unit ninexnine_unit_529(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01017)
);

ninexnine_unit ninexnine_unit_530(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02017)
);

assign C0017=c00017+c01017+c02017;
assign A0017=(C0017>=0)?1:0;

assign P1017=A0017;

ninexnine_unit ninexnine_unit_531(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00027)
);

ninexnine_unit ninexnine_unit_532(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01027)
);

ninexnine_unit ninexnine_unit_533(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02027)
);

assign C0027=c00027+c01027+c02027;
assign A0027=(C0027>=0)?1:0;

assign P1027=A0027;

ninexnine_unit ninexnine_unit_534(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00037)
);

ninexnine_unit ninexnine_unit_535(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01037)
);

ninexnine_unit ninexnine_unit_536(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02037)
);

assign C0037=c00037+c01037+c02037;
assign A0037=(C0037>=0)?1:0;

assign P1037=A0037;

ninexnine_unit ninexnine_unit_537(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00047)
);

ninexnine_unit ninexnine_unit_538(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01047)
);

ninexnine_unit ninexnine_unit_539(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02047)
);

assign C0047=c00047+c01047+c02047;
assign A0047=(C0047>=0)?1:0;

assign P1047=A0047;

ninexnine_unit ninexnine_unit_540(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00107)
);

ninexnine_unit ninexnine_unit_541(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01107)
);

ninexnine_unit ninexnine_unit_542(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02107)
);

assign C0107=c00107+c01107+c02107;
assign A0107=(C0107>=0)?1:0;

assign P1107=A0107;

ninexnine_unit ninexnine_unit_543(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00117)
);

ninexnine_unit ninexnine_unit_544(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01117)
);

ninexnine_unit ninexnine_unit_545(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02117)
);

assign C0117=c00117+c01117+c02117;
assign A0117=(C0117>=0)?1:0;

assign P1117=A0117;

ninexnine_unit ninexnine_unit_546(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00127)
);

ninexnine_unit ninexnine_unit_547(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01127)
);

ninexnine_unit ninexnine_unit_548(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02127)
);

assign C0127=c00127+c01127+c02127;
assign A0127=(C0127>=0)?1:0;

assign P1127=A0127;

ninexnine_unit ninexnine_unit_549(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00137)
);

ninexnine_unit ninexnine_unit_550(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01137)
);

ninexnine_unit ninexnine_unit_551(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02137)
);

assign C0137=c00137+c01137+c02137;
assign A0137=(C0137>=0)?1:0;

assign P1137=A0137;

ninexnine_unit ninexnine_unit_552(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00147)
);

ninexnine_unit ninexnine_unit_553(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01147)
);

ninexnine_unit ninexnine_unit_554(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02147)
);

assign C0147=c00147+c01147+c02147;
assign A0147=(C0147>=0)?1:0;

assign P1147=A0147;

ninexnine_unit ninexnine_unit_555(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00207)
);

ninexnine_unit ninexnine_unit_556(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01207)
);

ninexnine_unit ninexnine_unit_557(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02207)
);

assign C0207=c00207+c01207+c02207;
assign A0207=(C0207>=0)?1:0;

assign P1207=A0207;

ninexnine_unit ninexnine_unit_558(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00217)
);

ninexnine_unit ninexnine_unit_559(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01217)
);

ninexnine_unit ninexnine_unit_560(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02217)
);

assign C0217=c00217+c01217+c02217;
assign A0217=(C0217>=0)?1:0;

assign P1217=A0217;

ninexnine_unit ninexnine_unit_561(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00227)
);

ninexnine_unit ninexnine_unit_562(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01227)
);

ninexnine_unit ninexnine_unit_563(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02227)
);

assign C0227=c00227+c01227+c02227;
assign A0227=(C0227>=0)?1:0;

assign P1227=A0227;

ninexnine_unit ninexnine_unit_564(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00237)
);

ninexnine_unit ninexnine_unit_565(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01237)
);

ninexnine_unit ninexnine_unit_566(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02237)
);

assign C0237=c00237+c01237+c02237;
assign A0237=(C0237>=0)?1:0;

assign P1237=A0237;

ninexnine_unit ninexnine_unit_567(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00247)
);

ninexnine_unit ninexnine_unit_568(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01247)
);

ninexnine_unit ninexnine_unit_569(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02247)
);

assign C0247=c00247+c01247+c02247;
assign A0247=(C0247>=0)?1:0;

assign P1247=A0247;

ninexnine_unit ninexnine_unit_570(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00307)
);

ninexnine_unit ninexnine_unit_571(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01307)
);

ninexnine_unit ninexnine_unit_572(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02307)
);

assign C0307=c00307+c01307+c02307;
assign A0307=(C0307>=0)?1:0;

assign P1307=A0307;

ninexnine_unit ninexnine_unit_573(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00317)
);

ninexnine_unit ninexnine_unit_574(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01317)
);

ninexnine_unit ninexnine_unit_575(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02317)
);

assign C0317=c00317+c01317+c02317;
assign A0317=(C0317>=0)?1:0;

assign P1317=A0317;

ninexnine_unit ninexnine_unit_576(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00327)
);

ninexnine_unit ninexnine_unit_577(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01327)
);

ninexnine_unit ninexnine_unit_578(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02327)
);

assign C0327=c00327+c01327+c02327;
assign A0327=(C0327>=0)?1:0;

assign P1327=A0327;

ninexnine_unit ninexnine_unit_579(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00337)
);

ninexnine_unit ninexnine_unit_580(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01337)
);

ninexnine_unit ninexnine_unit_581(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02337)
);

assign C0337=c00337+c01337+c02337;
assign A0337=(C0337>=0)?1:0;

assign P1337=A0337;

ninexnine_unit ninexnine_unit_582(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00347)
);

ninexnine_unit ninexnine_unit_583(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01347)
);

ninexnine_unit ninexnine_unit_584(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02347)
);

assign C0347=c00347+c01347+c02347;
assign A0347=(C0347>=0)?1:0;

assign P1347=A0347;

ninexnine_unit ninexnine_unit_585(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00407)
);

ninexnine_unit ninexnine_unit_586(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01407)
);

ninexnine_unit ninexnine_unit_587(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02407)
);

assign C0407=c00407+c01407+c02407;
assign A0407=(C0407>=0)?1:0;

assign P1407=A0407;

ninexnine_unit ninexnine_unit_588(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00417)
);

ninexnine_unit ninexnine_unit_589(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01417)
);

ninexnine_unit ninexnine_unit_590(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02417)
);

assign C0417=c00417+c01417+c02417;
assign A0417=(C0417>=0)?1:0;

assign P1417=A0417;

ninexnine_unit ninexnine_unit_591(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00427)
);

ninexnine_unit ninexnine_unit_592(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01427)
);

ninexnine_unit ninexnine_unit_593(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02427)
);

assign C0427=c00427+c01427+c02427;
assign A0427=(C0427>=0)?1:0;

assign P1427=A0427;

ninexnine_unit ninexnine_unit_594(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00437)
);

ninexnine_unit ninexnine_unit_595(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01437)
);

ninexnine_unit ninexnine_unit_596(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02437)
);

assign C0437=c00437+c01437+c02437;
assign A0437=(C0437>=0)?1:0;

assign P1437=A0437;

ninexnine_unit ninexnine_unit_597(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W07000),
				.b1(W07010),
				.b2(W07020),
				.b3(W07100),
				.b4(W07110),
				.b5(W07120),
				.b6(W07200),
				.b7(W07210),
				.b8(W07220),
				.c(c00447)
);

ninexnine_unit ninexnine_unit_598(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W07001),
				.b1(W07011),
				.b2(W07021),
				.b3(W07101),
				.b4(W07111),
				.b5(W07121),
				.b6(W07201),
				.b7(W07211),
				.b8(W07221),
				.c(c01447)
);

ninexnine_unit ninexnine_unit_599(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W07002),
				.b1(W07012),
				.b2(W07022),
				.b3(W07102),
				.b4(W07112),
				.b5(W07122),
				.b6(W07202),
				.b7(W07212),
				.b8(W07222),
				.c(c02447)
);

assign C0447=c00447+c01447+c02447;
assign A0447=(C0447>=0)?1:0;

assign P1447=A0447;

ninexnine_unit ninexnine_unit_600(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00008)
);

ninexnine_unit ninexnine_unit_601(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01008)
);

ninexnine_unit ninexnine_unit_602(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02008)
);

assign C0008=c00008+c01008+c02008;
assign A0008=(C0008>=0)?1:0;

assign P1008=A0008;

ninexnine_unit ninexnine_unit_603(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00018)
);

ninexnine_unit ninexnine_unit_604(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01018)
);

ninexnine_unit ninexnine_unit_605(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02018)
);

assign C0018=c00018+c01018+c02018;
assign A0018=(C0018>=0)?1:0;

assign P1018=A0018;

ninexnine_unit ninexnine_unit_606(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00028)
);

ninexnine_unit ninexnine_unit_607(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01028)
);

ninexnine_unit ninexnine_unit_608(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02028)
);

assign C0028=c00028+c01028+c02028;
assign A0028=(C0028>=0)?1:0;

assign P1028=A0028;

ninexnine_unit ninexnine_unit_609(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00038)
);

ninexnine_unit ninexnine_unit_610(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01038)
);

ninexnine_unit ninexnine_unit_611(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02038)
);

assign C0038=c00038+c01038+c02038;
assign A0038=(C0038>=0)?1:0;

assign P1038=A0038;

ninexnine_unit ninexnine_unit_612(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00048)
);

ninexnine_unit ninexnine_unit_613(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01048)
);

ninexnine_unit ninexnine_unit_614(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02048)
);

assign C0048=c00048+c01048+c02048;
assign A0048=(C0048>=0)?1:0;

assign P1048=A0048;

ninexnine_unit ninexnine_unit_615(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00108)
);

ninexnine_unit ninexnine_unit_616(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01108)
);

ninexnine_unit ninexnine_unit_617(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02108)
);

assign C0108=c00108+c01108+c02108;
assign A0108=(C0108>=0)?1:0;

assign P1108=A0108;

ninexnine_unit ninexnine_unit_618(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00118)
);

ninexnine_unit ninexnine_unit_619(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01118)
);

ninexnine_unit ninexnine_unit_620(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02118)
);

assign C0118=c00118+c01118+c02118;
assign A0118=(C0118>=0)?1:0;

assign P1118=A0118;

ninexnine_unit ninexnine_unit_621(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00128)
);

ninexnine_unit ninexnine_unit_622(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01128)
);

ninexnine_unit ninexnine_unit_623(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02128)
);

assign C0128=c00128+c01128+c02128;
assign A0128=(C0128>=0)?1:0;

assign P1128=A0128;

ninexnine_unit ninexnine_unit_624(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00138)
);

ninexnine_unit ninexnine_unit_625(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01138)
);

ninexnine_unit ninexnine_unit_626(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02138)
);

assign C0138=c00138+c01138+c02138;
assign A0138=(C0138>=0)?1:0;

assign P1138=A0138;

ninexnine_unit ninexnine_unit_627(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00148)
);

ninexnine_unit ninexnine_unit_628(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01148)
);

ninexnine_unit ninexnine_unit_629(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02148)
);

assign C0148=c00148+c01148+c02148;
assign A0148=(C0148>=0)?1:0;

assign P1148=A0148;

ninexnine_unit ninexnine_unit_630(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00208)
);

ninexnine_unit ninexnine_unit_631(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01208)
);

ninexnine_unit ninexnine_unit_632(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02208)
);

assign C0208=c00208+c01208+c02208;
assign A0208=(C0208>=0)?1:0;

assign P1208=A0208;

ninexnine_unit ninexnine_unit_633(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00218)
);

ninexnine_unit ninexnine_unit_634(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01218)
);

ninexnine_unit ninexnine_unit_635(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02218)
);

assign C0218=c00218+c01218+c02218;
assign A0218=(C0218>=0)?1:0;

assign P1218=A0218;

ninexnine_unit ninexnine_unit_636(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00228)
);

ninexnine_unit ninexnine_unit_637(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01228)
);

ninexnine_unit ninexnine_unit_638(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02228)
);

assign C0228=c00228+c01228+c02228;
assign A0228=(C0228>=0)?1:0;

assign P1228=A0228;

ninexnine_unit ninexnine_unit_639(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00238)
);

ninexnine_unit ninexnine_unit_640(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01238)
);

ninexnine_unit ninexnine_unit_641(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02238)
);

assign C0238=c00238+c01238+c02238;
assign A0238=(C0238>=0)?1:0;

assign P1238=A0238;

ninexnine_unit ninexnine_unit_642(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00248)
);

ninexnine_unit ninexnine_unit_643(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01248)
);

ninexnine_unit ninexnine_unit_644(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02248)
);

assign C0248=c00248+c01248+c02248;
assign A0248=(C0248>=0)?1:0;

assign P1248=A0248;

ninexnine_unit ninexnine_unit_645(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00308)
);

ninexnine_unit ninexnine_unit_646(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01308)
);

ninexnine_unit ninexnine_unit_647(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02308)
);

assign C0308=c00308+c01308+c02308;
assign A0308=(C0308>=0)?1:0;

assign P1308=A0308;

ninexnine_unit ninexnine_unit_648(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00318)
);

ninexnine_unit ninexnine_unit_649(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01318)
);

ninexnine_unit ninexnine_unit_650(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02318)
);

assign C0318=c00318+c01318+c02318;
assign A0318=(C0318>=0)?1:0;

assign P1318=A0318;

ninexnine_unit ninexnine_unit_651(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00328)
);

ninexnine_unit ninexnine_unit_652(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01328)
);

ninexnine_unit ninexnine_unit_653(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02328)
);

assign C0328=c00328+c01328+c02328;
assign A0328=(C0328>=0)?1:0;

assign P1328=A0328;

ninexnine_unit ninexnine_unit_654(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00338)
);

ninexnine_unit ninexnine_unit_655(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01338)
);

ninexnine_unit ninexnine_unit_656(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02338)
);

assign C0338=c00338+c01338+c02338;
assign A0338=(C0338>=0)?1:0;

assign P1338=A0338;

ninexnine_unit ninexnine_unit_657(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00348)
);

ninexnine_unit ninexnine_unit_658(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01348)
);

ninexnine_unit ninexnine_unit_659(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02348)
);

assign C0348=c00348+c01348+c02348;
assign A0348=(C0348>=0)?1:0;

assign P1348=A0348;

ninexnine_unit ninexnine_unit_660(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00408)
);

ninexnine_unit ninexnine_unit_661(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01408)
);

ninexnine_unit ninexnine_unit_662(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02408)
);

assign C0408=c00408+c01408+c02408;
assign A0408=(C0408>=0)?1:0;

assign P1408=A0408;

ninexnine_unit ninexnine_unit_663(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00418)
);

ninexnine_unit ninexnine_unit_664(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01418)
);

ninexnine_unit ninexnine_unit_665(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02418)
);

assign C0418=c00418+c01418+c02418;
assign A0418=(C0418>=0)?1:0;

assign P1418=A0418;

ninexnine_unit ninexnine_unit_666(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00428)
);

ninexnine_unit ninexnine_unit_667(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01428)
);

ninexnine_unit ninexnine_unit_668(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02428)
);

assign C0428=c00428+c01428+c02428;
assign A0428=(C0428>=0)?1:0;

assign P1428=A0428;

ninexnine_unit ninexnine_unit_669(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00438)
);

ninexnine_unit ninexnine_unit_670(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01438)
);

ninexnine_unit ninexnine_unit_671(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02438)
);

assign C0438=c00438+c01438+c02438;
assign A0438=(C0438>=0)?1:0;

assign P1438=A0438;

ninexnine_unit ninexnine_unit_672(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W08000),
				.b1(W08010),
				.b2(W08020),
				.b3(W08100),
				.b4(W08110),
				.b5(W08120),
				.b6(W08200),
				.b7(W08210),
				.b8(W08220),
				.c(c00448)
);

ninexnine_unit ninexnine_unit_673(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W08001),
				.b1(W08011),
				.b2(W08021),
				.b3(W08101),
				.b4(W08111),
				.b5(W08121),
				.b6(W08201),
				.b7(W08211),
				.b8(W08221),
				.c(c01448)
);

ninexnine_unit ninexnine_unit_674(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W08002),
				.b1(W08012),
				.b2(W08022),
				.b3(W08102),
				.b4(W08112),
				.b5(W08122),
				.b6(W08202),
				.b7(W08212),
				.b8(W08222),
				.c(c02448)
);

assign C0448=c00448+c01448+c02448;
assign A0448=(C0448>=0)?1:0;

assign P1448=A0448;

ninexnine_unit ninexnine_unit_675(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00009)
);

ninexnine_unit ninexnine_unit_676(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01009)
);

ninexnine_unit ninexnine_unit_677(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02009)
);

assign C0009=c00009+c01009+c02009;
assign A0009=(C0009>=0)?1:0;

assign P1009=A0009;

ninexnine_unit ninexnine_unit_678(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00019)
);

ninexnine_unit ninexnine_unit_679(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01019)
);

ninexnine_unit ninexnine_unit_680(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02019)
);

assign C0019=c00019+c01019+c02019;
assign A0019=(C0019>=0)?1:0;

assign P1019=A0019;

ninexnine_unit ninexnine_unit_681(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00029)
);

ninexnine_unit ninexnine_unit_682(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01029)
);

ninexnine_unit ninexnine_unit_683(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02029)
);

assign C0029=c00029+c01029+c02029;
assign A0029=(C0029>=0)?1:0;

assign P1029=A0029;

ninexnine_unit ninexnine_unit_684(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00039)
);

ninexnine_unit ninexnine_unit_685(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01039)
);

ninexnine_unit ninexnine_unit_686(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02039)
);

assign C0039=c00039+c01039+c02039;
assign A0039=(C0039>=0)?1:0;

assign P1039=A0039;

ninexnine_unit ninexnine_unit_687(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00049)
);

ninexnine_unit ninexnine_unit_688(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01049)
);

ninexnine_unit ninexnine_unit_689(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02049)
);

assign C0049=c00049+c01049+c02049;
assign A0049=(C0049>=0)?1:0;

assign P1049=A0049;

ninexnine_unit ninexnine_unit_690(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00109)
);

ninexnine_unit ninexnine_unit_691(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01109)
);

ninexnine_unit ninexnine_unit_692(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02109)
);

assign C0109=c00109+c01109+c02109;
assign A0109=(C0109>=0)?1:0;

assign P1109=A0109;

ninexnine_unit ninexnine_unit_693(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00119)
);

ninexnine_unit ninexnine_unit_694(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01119)
);

ninexnine_unit ninexnine_unit_695(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02119)
);

assign C0119=c00119+c01119+c02119;
assign A0119=(C0119>=0)?1:0;

assign P1119=A0119;

ninexnine_unit ninexnine_unit_696(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00129)
);

ninexnine_unit ninexnine_unit_697(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01129)
);

ninexnine_unit ninexnine_unit_698(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02129)
);

assign C0129=c00129+c01129+c02129;
assign A0129=(C0129>=0)?1:0;

assign P1129=A0129;

ninexnine_unit ninexnine_unit_699(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00139)
);

ninexnine_unit ninexnine_unit_700(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01139)
);

ninexnine_unit ninexnine_unit_701(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02139)
);

assign C0139=c00139+c01139+c02139;
assign A0139=(C0139>=0)?1:0;

assign P1139=A0139;

ninexnine_unit ninexnine_unit_702(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00149)
);

ninexnine_unit ninexnine_unit_703(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01149)
);

ninexnine_unit ninexnine_unit_704(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02149)
);

assign C0149=c00149+c01149+c02149;
assign A0149=(C0149>=0)?1:0;

assign P1149=A0149;

ninexnine_unit ninexnine_unit_705(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00209)
);

ninexnine_unit ninexnine_unit_706(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01209)
);

ninexnine_unit ninexnine_unit_707(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02209)
);

assign C0209=c00209+c01209+c02209;
assign A0209=(C0209>=0)?1:0;

assign P1209=A0209;

ninexnine_unit ninexnine_unit_708(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00219)
);

ninexnine_unit ninexnine_unit_709(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01219)
);

ninexnine_unit ninexnine_unit_710(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02219)
);

assign C0219=c00219+c01219+c02219;
assign A0219=(C0219>=0)?1:0;

assign P1219=A0219;

ninexnine_unit ninexnine_unit_711(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00229)
);

ninexnine_unit ninexnine_unit_712(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01229)
);

ninexnine_unit ninexnine_unit_713(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02229)
);

assign C0229=c00229+c01229+c02229;
assign A0229=(C0229>=0)?1:0;

assign P1229=A0229;

ninexnine_unit ninexnine_unit_714(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00239)
);

ninexnine_unit ninexnine_unit_715(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01239)
);

ninexnine_unit ninexnine_unit_716(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02239)
);

assign C0239=c00239+c01239+c02239;
assign A0239=(C0239>=0)?1:0;

assign P1239=A0239;

ninexnine_unit ninexnine_unit_717(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00249)
);

ninexnine_unit ninexnine_unit_718(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01249)
);

ninexnine_unit ninexnine_unit_719(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02249)
);

assign C0249=c00249+c01249+c02249;
assign A0249=(C0249>=0)?1:0;

assign P1249=A0249;

ninexnine_unit ninexnine_unit_720(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00309)
);

ninexnine_unit ninexnine_unit_721(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01309)
);

ninexnine_unit ninexnine_unit_722(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02309)
);

assign C0309=c00309+c01309+c02309;
assign A0309=(C0309>=0)?1:0;

assign P1309=A0309;

ninexnine_unit ninexnine_unit_723(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00319)
);

ninexnine_unit ninexnine_unit_724(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01319)
);

ninexnine_unit ninexnine_unit_725(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02319)
);

assign C0319=c00319+c01319+c02319;
assign A0319=(C0319>=0)?1:0;

assign P1319=A0319;

ninexnine_unit ninexnine_unit_726(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00329)
);

ninexnine_unit ninexnine_unit_727(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01329)
);

ninexnine_unit ninexnine_unit_728(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02329)
);

assign C0329=c00329+c01329+c02329;
assign A0329=(C0329>=0)?1:0;

assign P1329=A0329;

ninexnine_unit ninexnine_unit_729(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00339)
);

ninexnine_unit ninexnine_unit_730(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01339)
);

ninexnine_unit ninexnine_unit_731(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02339)
);

assign C0339=c00339+c01339+c02339;
assign A0339=(C0339>=0)?1:0;

assign P1339=A0339;

ninexnine_unit ninexnine_unit_732(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00349)
);

ninexnine_unit ninexnine_unit_733(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01349)
);

ninexnine_unit ninexnine_unit_734(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02349)
);

assign C0349=c00349+c01349+c02349;
assign A0349=(C0349>=0)?1:0;

assign P1349=A0349;

ninexnine_unit ninexnine_unit_735(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00409)
);

ninexnine_unit ninexnine_unit_736(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01409)
);

ninexnine_unit ninexnine_unit_737(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02409)
);

assign C0409=c00409+c01409+c02409;
assign A0409=(C0409>=0)?1:0;

assign P1409=A0409;

ninexnine_unit ninexnine_unit_738(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00419)
);

ninexnine_unit ninexnine_unit_739(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01419)
);

ninexnine_unit ninexnine_unit_740(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02419)
);

assign C0419=c00419+c01419+c02419;
assign A0419=(C0419>=0)?1:0;

assign P1419=A0419;

ninexnine_unit ninexnine_unit_741(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00429)
);

ninexnine_unit ninexnine_unit_742(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01429)
);

ninexnine_unit ninexnine_unit_743(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02429)
);

assign C0429=c00429+c01429+c02429;
assign A0429=(C0429>=0)?1:0;

assign P1429=A0429;

ninexnine_unit ninexnine_unit_744(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00439)
);

ninexnine_unit ninexnine_unit_745(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01439)
);

ninexnine_unit ninexnine_unit_746(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02439)
);

assign C0439=c00439+c01439+c02439;
assign A0439=(C0439>=0)?1:0;

assign P1439=A0439;

ninexnine_unit ninexnine_unit_747(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W09000),
				.b1(W09010),
				.b2(W09020),
				.b3(W09100),
				.b4(W09110),
				.b5(W09120),
				.b6(W09200),
				.b7(W09210),
				.b8(W09220),
				.c(c00449)
);

ninexnine_unit ninexnine_unit_748(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W09001),
				.b1(W09011),
				.b2(W09021),
				.b3(W09101),
				.b4(W09111),
				.b5(W09121),
				.b6(W09201),
				.b7(W09211),
				.b8(W09221),
				.c(c01449)
);

ninexnine_unit ninexnine_unit_749(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W09002),
				.b1(W09012),
				.b2(W09022),
				.b3(W09102),
				.b4(W09112),
				.b5(W09122),
				.b6(W09202),
				.b7(W09212),
				.b8(W09222),
				.c(c02449)
);

assign C0449=c00449+c01449+c02449;
assign A0449=(C0449>=0)?1:0;

assign P1449=A0449;

ninexnine_unit ninexnine_unit_750(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0000A)
);

ninexnine_unit ninexnine_unit_751(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0100A)
);

ninexnine_unit ninexnine_unit_752(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0200A)
);

assign C000A=c0000A+c0100A+c0200A;
assign A000A=(C000A>=0)?1:0;

assign P100A=A000A;

ninexnine_unit ninexnine_unit_753(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0001A)
);

ninexnine_unit ninexnine_unit_754(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0101A)
);

ninexnine_unit ninexnine_unit_755(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0201A)
);

assign C001A=c0001A+c0101A+c0201A;
assign A001A=(C001A>=0)?1:0;

assign P101A=A001A;

ninexnine_unit ninexnine_unit_756(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0002A)
);

ninexnine_unit ninexnine_unit_757(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0102A)
);

ninexnine_unit ninexnine_unit_758(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0202A)
);

assign C002A=c0002A+c0102A+c0202A;
assign A002A=(C002A>=0)?1:0;

assign P102A=A002A;

ninexnine_unit ninexnine_unit_759(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0003A)
);

ninexnine_unit ninexnine_unit_760(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0103A)
);

ninexnine_unit ninexnine_unit_761(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0203A)
);

assign C003A=c0003A+c0103A+c0203A;
assign A003A=(C003A>=0)?1:0;

assign P103A=A003A;

ninexnine_unit ninexnine_unit_762(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0004A)
);

ninexnine_unit ninexnine_unit_763(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0104A)
);

ninexnine_unit ninexnine_unit_764(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0204A)
);

assign C004A=c0004A+c0104A+c0204A;
assign A004A=(C004A>=0)?1:0;

assign P104A=A004A;

ninexnine_unit ninexnine_unit_765(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0010A)
);

ninexnine_unit ninexnine_unit_766(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0110A)
);

ninexnine_unit ninexnine_unit_767(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0210A)
);

assign C010A=c0010A+c0110A+c0210A;
assign A010A=(C010A>=0)?1:0;

assign P110A=A010A;

ninexnine_unit ninexnine_unit_768(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0011A)
);

ninexnine_unit ninexnine_unit_769(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0111A)
);

ninexnine_unit ninexnine_unit_770(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0211A)
);

assign C011A=c0011A+c0111A+c0211A;
assign A011A=(C011A>=0)?1:0;

assign P111A=A011A;

ninexnine_unit ninexnine_unit_771(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0012A)
);

ninexnine_unit ninexnine_unit_772(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0112A)
);

ninexnine_unit ninexnine_unit_773(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0212A)
);

assign C012A=c0012A+c0112A+c0212A;
assign A012A=(C012A>=0)?1:0;

assign P112A=A012A;

ninexnine_unit ninexnine_unit_774(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0013A)
);

ninexnine_unit ninexnine_unit_775(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0113A)
);

ninexnine_unit ninexnine_unit_776(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0213A)
);

assign C013A=c0013A+c0113A+c0213A;
assign A013A=(C013A>=0)?1:0;

assign P113A=A013A;

ninexnine_unit ninexnine_unit_777(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0014A)
);

ninexnine_unit ninexnine_unit_778(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0114A)
);

ninexnine_unit ninexnine_unit_779(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0214A)
);

assign C014A=c0014A+c0114A+c0214A;
assign A014A=(C014A>=0)?1:0;

assign P114A=A014A;

ninexnine_unit ninexnine_unit_780(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0020A)
);

ninexnine_unit ninexnine_unit_781(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0120A)
);

ninexnine_unit ninexnine_unit_782(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0220A)
);

assign C020A=c0020A+c0120A+c0220A;
assign A020A=(C020A>=0)?1:0;

assign P120A=A020A;

ninexnine_unit ninexnine_unit_783(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0021A)
);

ninexnine_unit ninexnine_unit_784(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0121A)
);

ninexnine_unit ninexnine_unit_785(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0221A)
);

assign C021A=c0021A+c0121A+c0221A;
assign A021A=(C021A>=0)?1:0;

assign P121A=A021A;

ninexnine_unit ninexnine_unit_786(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0022A)
);

ninexnine_unit ninexnine_unit_787(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0122A)
);

ninexnine_unit ninexnine_unit_788(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0222A)
);

assign C022A=c0022A+c0122A+c0222A;
assign A022A=(C022A>=0)?1:0;

assign P122A=A022A;

ninexnine_unit ninexnine_unit_789(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0023A)
);

ninexnine_unit ninexnine_unit_790(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0123A)
);

ninexnine_unit ninexnine_unit_791(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0223A)
);

assign C023A=c0023A+c0123A+c0223A;
assign A023A=(C023A>=0)?1:0;

assign P123A=A023A;

ninexnine_unit ninexnine_unit_792(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0024A)
);

ninexnine_unit ninexnine_unit_793(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0124A)
);

ninexnine_unit ninexnine_unit_794(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0224A)
);

assign C024A=c0024A+c0124A+c0224A;
assign A024A=(C024A>=0)?1:0;

assign P124A=A024A;

ninexnine_unit ninexnine_unit_795(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0030A)
);

ninexnine_unit ninexnine_unit_796(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0130A)
);

ninexnine_unit ninexnine_unit_797(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0230A)
);

assign C030A=c0030A+c0130A+c0230A;
assign A030A=(C030A>=0)?1:0;

assign P130A=A030A;

ninexnine_unit ninexnine_unit_798(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0031A)
);

ninexnine_unit ninexnine_unit_799(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0131A)
);

ninexnine_unit ninexnine_unit_800(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0231A)
);

assign C031A=c0031A+c0131A+c0231A;
assign A031A=(C031A>=0)?1:0;

assign P131A=A031A;

ninexnine_unit ninexnine_unit_801(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0032A)
);

ninexnine_unit ninexnine_unit_802(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0132A)
);

ninexnine_unit ninexnine_unit_803(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0232A)
);

assign C032A=c0032A+c0132A+c0232A;
assign A032A=(C032A>=0)?1:0;

assign P132A=A032A;

ninexnine_unit ninexnine_unit_804(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0033A)
);

ninexnine_unit ninexnine_unit_805(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0133A)
);

ninexnine_unit ninexnine_unit_806(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0233A)
);

assign C033A=c0033A+c0133A+c0233A;
assign A033A=(C033A>=0)?1:0;

assign P133A=A033A;

ninexnine_unit ninexnine_unit_807(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0034A)
);

ninexnine_unit ninexnine_unit_808(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0134A)
);

ninexnine_unit ninexnine_unit_809(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0234A)
);

assign C034A=c0034A+c0134A+c0234A;
assign A034A=(C034A>=0)?1:0;

assign P134A=A034A;

ninexnine_unit ninexnine_unit_810(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0040A)
);

ninexnine_unit ninexnine_unit_811(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0140A)
);

ninexnine_unit ninexnine_unit_812(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0240A)
);

assign C040A=c0040A+c0140A+c0240A;
assign A040A=(C040A>=0)?1:0;

assign P140A=A040A;

ninexnine_unit ninexnine_unit_813(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0041A)
);

ninexnine_unit ninexnine_unit_814(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0141A)
);

ninexnine_unit ninexnine_unit_815(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0241A)
);

assign C041A=c0041A+c0141A+c0241A;
assign A041A=(C041A>=0)?1:0;

assign P141A=A041A;

ninexnine_unit ninexnine_unit_816(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0042A)
);

ninexnine_unit ninexnine_unit_817(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0142A)
);

ninexnine_unit ninexnine_unit_818(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0242A)
);

assign C042A=c0042A+c0142A+c0242A;
assign A042A=(C042A>=0)?1:0;

assign P142A=A042A;

ninexnine_unit ninexnine_unit_819(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0043A)
);

ninexnine_unit ninexnine_unit_820(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0143A)
);

ninexnine_unit ninexnine_unit_821(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0243A)
);

assign C043A=c0043A+c0143A+c0243A;
assign A043A=(C043A>=0)?1:0;

assign P143A=A043A;

ninexnine_unit ninexnine_unit_822(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W0A000),
				.b1(W0A010),
				.b2(W0A020),
				.b3(W0A100),
				.b4(W0A110),
				.b5(W0A120),
				.b6(W0A200),
				.b7(W0A210),
				.b8(W0A220),
				.c(c0044A)
);

ninexnine_unit ninexnine_unit_823(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W0A001),
				.b1(W0A011),
				.b2(W0A021),
				.b3(W0A101),
				.b4(W0A111),
				.b5(W0A121),
				.b6(W0A201),
				.b7(W0A211),
				.b8(W0A221),
				.c(c0144A)
);

ninexnine_unit ninexnine_unit_824(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W0A002),
				.b1(W0A012),
				.b2(W0A022),
				.b3(W0A102),
				.b4(W0A112),
				.b5(W0A122),
				.b6(W0A202),
				.b7(W0A212),
				.b8(W0A222),
				.c(c0244A)
);

assign C044A=c0044A+c0144A+c0244A;
assign A044A=(C044A>=0)?1:0;

assign P144A=A044A;

ninexnine_unit ninexnine_unit_825(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0000B)
);

ninexnine_unit ninexnine_unit_826(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0100B)
);

ninexnine_unit ninexnine_unit_827(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0200B)
);

assign C000B=c0000B+c0100B+c0200B;
assign A000B=(C000B>=0)?1:0;

assign P100B=A000B;

ninexnine_unit ninexnine_unit_828(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0001B)
);

ninexnine_unit ninexnine_unit_829(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0101B)
);

ninexnine_unit ninexnine_unit_830(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0201B)
);

assign C001B=c0001B+c0101B+c0201B;
assign A001B=(C001B>=0)?1:0;

assign P101B=A001B;

ninexnine_unit ninexnine_unit_831(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0002B)
);

ninexnine_unit ninexnine_unit_832(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0102B)
);

ninexnine_unit ninexnine_unit_833(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0202B)
);

assign C002B=c0002B+c0102B+c0202B;
assign A002B=(C002B>=0)?1:0;

assign P102B=A002B;

ninexnine_unit ninexnine_unit_834(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0003B)
);

ninexnine_unit ninexnine_unit_835(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0103B)
);

ninexnine_unit ninexnine_unit_836(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0203B)
);

assign C003B=c0003B+c0103B+c0203B;
assign A003B=(C003B>=0)?1:0;

assign P103B=A003B;

ninexnine_unit ninexnine_unit_837(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0004B)
);

ninexnine_unit ninexnine_unit_838(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0104B)
);

ninexnine_unit ninexnine_unit_839(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0204B)
);

assign C004B=c0004B+c0104B+c0204B;
assign A004B=(C004B>=0)?1:0;

assign P104B=A004B;

ninexnine_unit ninexnine_unit_840(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0010B)
);

ninexnine_unit ninexnine_unit_841(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0110B)
);

ninexnine_unit ninexnine_unit_842(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0210B)
);

assign C010B=c0010B+c0110B+c0210B;
assign A010B=(C010B>=0)?1:0;

assign P110B=A010B;

ninexnine_unit ninexnine_unit_843(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0011B)
);

ninexnine_unit ninexnine_unit_844(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0111B)
);

ninexnine_unit ninexnine_unit_845(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0211B)
);

assign C011B=c0011B+c0111B+c0211B;
assign A011B=(C011B>=0)?1:0;

assign P111B=A011B;

ninexnine_unit ninexnine_unit_846(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0012B)
);

ninexnine_unit ninexnine_unit_847(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0112B)
);

ninexnine_unit ninexnine_unit_848(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0212B)
);

assign C012B=c0012B+c0112B+c0212B;
assign A012B=(C012B>=0)?1:0;

assign P112B=A012B;

ninexnine_unit ninexnine_unit_849(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0013B)
);

ninexnine_unit ninexnine_unit_850(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0113B)
);

ninexnine_unit ninexnine_unit_851(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0213B)
);

assign C013B=c0013B+c0113B+c0213B;
assign A013B=(C013B>=0)?1:0;

assign P113B=A013B;

ninexnine_unit ninexnine_unit_852(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0014B)
);

ninexnine_unit ninexnine_unit_853(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0114B)
);

ninexnine_unit ninexnine_unit_854(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0214B)
);

assign C014B=c0014B+c0114B+c0214B;
assign A014B=(C014B>=0)?1:0;

assign P114B=A014B;

ninexnine_unit ninexnine_unit_855(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0020B)
);

ninexnine_unit ninexnine_unit_856(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0120B)
);

ninexnine_unit ninexnine_unit_857(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0220B)
);

assign C020B=c0020B+c0120B+c0220B;
assign A020B=(C020B>=0)?1:0;

assign P120B=A020B;

ninexnine_unit ninexnine_unit_858(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0021B)
);

ninexnine_unit ninexnine_unit_859(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0121B)
);

ninexnine_unit ninexnine_unit_860(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0221B)
);

assign C021B=c0021B+c0121B+c0221B;
assign A021B=(C021B>=0)?1:0;

assign P121B=A021B;

ninexnine_unit ninexnine_unit_861(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0022B)
);

ninexnine_unit ninexnine_unit_862(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0122B)
);

ninexnine_unit ninexnine_unit_863(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0222B)
);

assign C022B=c0022B+c0122B+c0222B;
assign A022B=(C022B>=0)?1:0;

assign P122B=A022B;

ninexnine_unit ninexnine_unit_864(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0023B)
);

ninexnine_unit ninexnine_unit_865(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0123B)
);

ninexnine_unit ninexnine_unit_866(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0223B)
);

assign C023B=c0023B+c0123B+c0223B;
assign A023B=(C023B>=0)?1:0;

assign P123B=A023B;

ninexnine_unit ninexnine_unit_867(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0024B)
);

ninexnine_unit ninexnine_unit_868(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0124B)
);

ninexnine_unit ninexnine_unit_869(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0224B)
);

assign C024B=c0024B+c0124B+c0224B;
assign A024B=(C024B>=0)?1:0;

assign P124B=A024B;

ninexnine_unit ninexnine_unit_870(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0030B)
);

ninexnine_unit ninexnine_unit_871(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0130B)
);

ninexnine_unit ninexnine_unit_872(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0230B)
);

assign C030B=c0030B+c0130B+c0230B;
assign A030B=(C030B>=0)?1:0;

assign P130B=A030B;

ninexnine_unit ninexnine_unit_873(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0031B)
);

ninexnine_unit ninexnine_unit_874(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0131B)
);

ninexnine_unit ninexnine_unit_875(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0231B)
);

assign C031B=c0031B+c0131B+c0231B;
assign A031B=(C031B>=0)?1:0;

assign P131B=A031B;

ninexnine_unit ninexnine_unit_876(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0032B)
);

ninexnine_unit ninexnine_unit_877(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0132B)
);

ninexnine_unit ninexnine_unit_878(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0232B)
);

assign C032B=c0032B+c0132B+c0232B;
assign A032B=(C032B>=0)?1:0;

assign P132B=A032B;

ninexnine_unit ninexnine_unit_879(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0033B)
);

ninexnine_unit ninexnine_unit_880(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0133B)
);

ninexnine_unit ninexnine_unit_881(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0233B)
);

assign C033B=c0033B+c0133B+c0233B;
assign A033B=(C033B>=0)?1:0;

assign P133B=A033B;

ninexnine_unit ninexnine_unit_882(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0034B)
);

ninexnine_unit ninexnine_unit_883(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0134B)
);

ninexnine_unit ninexnine_unit_884(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0234B)
);

assign C034B=c0034B+c0134B+c0234B;
assign A034B=(C034B>=0)?1:0;

assign P134B=A034B;

ninexnine_unit ninexnine_unit_885(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0040B)
);

ninexnine_unit ninexnine_unit_886(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0140B)
);

ninexnine_unit ninexnine_unit_887(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0240B)
);

assign C040B=c0040B+c0140B+c0240B;
assign A040B=(C040B>=0)?1:0;

assign P140B=A040B;

ninexnine_unit ninexnine_unit_888(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0041B)
);

ninexnine_unit ninexnine_unit_889(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0141B)
);

ninexnine_unit ninexnine_unit_890(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0241B)
);

assign C041B=c0041B+c0141B+c0241B;
assign A041B=(C041B>=0)?1:0;

assign P141B=A041B;

ninexnine_unit ninexnine_unit_891(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0042B)
);

ninexnine_unit ninexnine_unit_892(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0142B)
);

ninexnine_unit ninexnine_unit_893(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0242B)
);

assign C042B=c0042B+c0142B+c0242B;
assign A042B=(C042B>=0)?1:0;

assign P142B=A042B;

ninexnine_unit ninexnine_unit_894(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0043B)
);

ninexnine_unit ninexnine_unit_895(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0143B)
);

ninexnine_unit ninexnine_unit_896(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0243B)
);

assign C043B=c0043B+c0143B+c0243B;
assign A043B=(C043B>=0)?1:0;

assign P143B=A043B;

ninexnine_unit ninexnine_unit_897(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W0B000),
				.b1(W0B010),
				.b2(W0B020),
				.b3(W0B100),
				.b4(W0B110),
				.b5(W0B120),
				.b6(W0B200),
				.b7(W0B210),
				.b8(W0B220),
				.c(c0044B)
);

ninexnine_unit ninexnine_unit_898(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W0B001),
				.b1(W0B011),
				.b2(W0B021),
				.b3(W0B101),
				.b4(W0B111),
				.b5(W0B121),
				.b6(W0B201),
				.b7(W0B211),
				.b8(W0B221),
				.c(c0144B)
);

ninexnine_unit ninexnine_unit_899(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W0B002),
				.b1(W0B012),
				.b2(W0B022),
				.b3(W0B102),
				.b4(W0B112),
				.b5(W0B122),
				.b6(W0B202),
				.b7(W0B212),
				.b8(W0B222),
				.c(c0244B)
);

assign C044B=c0044B+c0144B+c0244B;
assign A044B=(C044B>=0)?1:0;

assign P144B=A044B;

ninexnine_unit ninexnine_unit_900(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0000C)
);

ninexnine_unit ninexnine_unit_901(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0100C)
);

ninexnine_unit ninexnine_unit_902(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0200C)
);

assign C000C=c0000C+c0100C+c0200C;
assign A000C=(C000C>=0)?1:0;

assign P100C=A000C;

ninexnine_unit ninexnine_unit_903(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0001C)
);

ninexnine_unit ninexnine_unit_904(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0101C)
);

ninexnine_unit ninexnine_unit_905(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0201C)
);

assign C001C=c0001C+c0101C+c0201C;
assign A001C=(C001C>=0)?1:0;

assign P101C=A001C;

ninexnine_unit ninexnine_unit_906(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0002C)
);

ninexnine_unit ninexnine_unit_907(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0102C)
);

ninexnine_unit ninexnine_unit_908(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0202C)
);

assign C002C=c0002C+c0102C+c0202C;
assign A002C=(C002C>=0)?1:0;

assign P102C=A002C;

ninexnine_unit ninexnine_unit_909(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0003C)
);

ninexnine_unit ninexnine_unit_910(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0103C)
);

ninexnine_unit ninexnine_unit_911(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0203C)
);

assign C003C=c0003C+c0103C+c0203C;
assign A003C=(C003C>=0)?1:0;

assign P103C=A003C;

ninexnine_unit ninexnine_unit_912(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0004C)
);

ninexnine_unit ninexnine_unit_913(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0104C)
);

ninexnine_unit ninexnine_unit_914(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0204C)
);

assign C004C=c0004C+c0104C+c0204C;
assign A004C=(C004C>=0)?1:0;

assign P104C=A004C;

ninexnine_unit ninexnine_unit_915(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0010C)
);

ninexnine_unit ninexnine_unit_916(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0110C)
);

ninexnine_unit ninexnine_unit_917(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0210C)
);

assign C010C=c0010C+c0110C+c0210C;
assign A010C=(C010C>=0)?1:0;

assign P110C=A010C;

ninexnine_unit ninexnine_unit_918(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0011C)
);

ninexnine_unit ninexnine_unit_919(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0111C)
);

ninexnine_unit ninexnine_unit_920(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0211C)
);

assign C011C=c0011C+c0111C+c0211C;
assign A011C=(C011C>=0)?1:0;

assign P111C=A011C;

ninexnine_unit ninexnine_unit_921(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0012C)
);

ninexnine_unit ninexnine_unit_922(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0112C)
);

ninexnine_unit ninexnine_unit_923(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0212C)
);

assign C012C=c0012C+c0112C+c0212C;
assign A012C=(C012C>=0)?1:0;

assign P112C=A012C;

ninexnine_unit ninexnine_unit_924(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0013C)
);

ninexnine_unit ninexnine_unit_925(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0113C)
);

ninexnine_unit ninexnine_unit_926(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0213C)
);

assign C013C=c0013C+c0113C+c0213C;
assign A013C=(C013C>=0)?1:0;

assign P113C=A013C;

ninexnine_unit ninexnine_unit_927(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0014C)
);

ninexnine_unit ninexnine_unit_928(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0114C)
);

ninexnine_unit ninexnine_unit_929(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0214C)
);

assign C014C=c0014C+c0114C+c0214C;
assign A014C=(C014C>=0)?1:0;

assign P114C=A014C;

ninexnine_unit ninexnine_unit_930(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0020C)
);

ninexnine_unit ninexnine_unit_931(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0120C)
);

ninexnine_unit ninexnine_unit_932(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0220C)
);

assign C020C=c0020C+c0120C+c0220C;
assign A020C=(C020C>=0)?1:0;

assign P120C=A020C;

ninexnine_unit ninexnine_unit_933(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0021C)
);

ninexnine_unit ninexnine_unit_934(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0121C)
);

ninexnine_unit ninexnine_unit_935(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0221C)
);

assign C021C=c0021C+c0121C+c0221C;
assign A021C=(C021C>=0)?1:0;

assign P121C=A021C;

ninexnine_unit ninexnine_unit_936(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0022C)
);

ninexnine_unit ninexnine_unit_937(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0122C)
);

ninexnine_unit ninexnine_unit_938(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0222C)
);

assign C022C=c0022C+c0122C+c0222C;
assign A022C=(C022C>=0)?1:0;

assign P122C=A022C;

ninexnine_unit ninexnine_unit_939(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0023C)
);

ninexnine_unit ninexnine_unit_940(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0123C)
);

ninexnine_unit ninexnine_unit_941(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0223C)
);

assign C023C=c0023C+c0123C+c0223C;
assign A023C=(C023C>=0)?1:0;

assign P123C=A023C;

ninexnine_unit ninexnine_unit_942(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0024C)
);

ninexnine_unit ninexnine_unit_943(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0124C)
);

ninexnine_unit ninexnine_unit_944(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0224C)
);

assign C024C=c0024C+c0124C+c0224C;
assign A024C=(C024C>=0)?1:0;

assign P124C=A024C;

ninexnine_unit ninexnine_unit_945(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0030C)
);

ninexnine_unit ninexnine_unit_946(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0130C)
);

ninexnine_unit ninexnine_unit_947(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0230C)
);

assign C030C=c0030C+c0130C+c0230C;
assign A030C=(C030C>=0)?1:0;

assign P130C=A030C;

ninexnine_unit ninexnine_unit_948(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0031C)
);

ninexnine_unit ninexnine_unit_949(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0131C)
);

ninexnine_unit ninexnine_unit_950(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0231C)
);

assign C031C=c0031C+c0131C+c0231C;
assign A031C=(C031C>=0)?1:0;

assign P131C=A031C;

ninexnine_unit ninexnine_unit_951(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0032C)
);

ninexnine_unit ninexnine_unit_952(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0132C)
);

ninexnine_unit ninexnine_unit_953(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0232C)
);

assign C032C=c0032C+c0132C+c0232C;
assign A032C=(C032C>=0)?1:0;

assign P132C=A032C;

ninexnine_unit ninexnine_unit_954(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0033C)
);

ninexnine_unit ninexnine_unit_955(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0133C)
);

ninexnine_unit ninexnine_unit_956(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0233C)
);

assign C033C=c0033C+c0133C+c0233C;
assign A033C=(C033C>=0)?1:0;

assign P133C=A033C;

ninexnine_unit ninexnine_unit_957(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0034C)
);

ninexnine_unit ninexnine_unit_958(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0134C)
);

ninexnine_unit ninexnine_unit_959(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0234C)
);

assign C034C=c0034C+c0134C+c0234C;
assign A034C=(C034C>=0)?1:0;

assign P134C=A034C;

ninexnine_unit ninexnine_unit_960(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0040C)
);

ninexnine_unit ninexnine_unit_961(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0140C)
);

ninexnine_unit ninexnine_unit_962(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0240C)
);

assign C040C=c0040C+c0140C+c0240C;
assign A040C=(C040C>=0)?1:0;

assign P140C=A040C;

ninexnine_unit ninexnine_unit_963(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0041C)
);

ninexnine_unit ninexnine_unit_964(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0141C)
);

ninexnine_unit ninexnine_unit_965(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0241C)
);

assign C041C=c0041C+c0141C+c0241C;
assign A041C=(C041C>=0)?1:0;

assign P141C=A041C;

ninexnine_unit ninexnine_unit_966(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0042C)
);

ninexnine_unit ninexnine_unit_967(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0142C)
);

ninexnine_unit ninexnine_unit_968(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0242C)
);

assign C042C=c0042C+c0142C+c0242C;
assign A042C=(C042C>=0)?1:0;

assign P142C=A042C;

ninexnine_unit ninexnine_unit_969(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0043C)
);

ninexnine_unit ninexnine_unit_970(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0143C)
);

ninexnine_unit ninexnine_unit_971(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0243C)
);

assign C043C=c0043C+c0143C+c0243C;
assign A043C=(C043C>=0)?1:0;

assign P143C=A043C;

ninexnine_unit ninexnine_unit_972(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W0C000),
				.b1(W0C010),
				.b2(W0C020),
				.b3(W0C100),
				.b4(W0C110),
				.b5(W0C120),
				.b6(W0C200),
				.b7(W0C210),
				.b8(W0C220),
				.c(c0044C)
);

ninexnine_unit ninexnine_unit_973(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W0C001),
				.b1(W0C011),
				.b2(W0C021),
				.b3(W0C101),
				.b4(W0C111),
				.b5(W0C121),
				.b6(W0C201),
				.b7(W0C211),
				.b8(W0C221),
				.c(c0144C)
);

ninexnine_unit ninexnine_unit_974(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W0C002),
				.b1(W0C012),
				.b2(W0C022),
				.b3(W0C102),
				.b4(W0C112),
				.b5(W0C122),
				.b6(W0C202),
				.b7(W0C212),
				.b8(W0C222),
				.c(c0244C)
);

assign C044C=c0044C+c0144C+c0244C;
assign A044C=(C044C>=0)?1:0;

assign P144C=A044C;

ninexnine_unit ninexnine_unit_975(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0000D)
);

ninexnine_unit ninexnine_unit_976(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0100D)
);

ninexnine_unit ninexnine_unit_977(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0200D)
);

assign C000D=c0000D+c0100D+c0200D;
assign A000D=(C000D>=0)?1:0;

assign P100D=A000D;

ninexnine_unit ninexnine_unit_978(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0001D)
);

ninexnine_unit ninexnine_unit_979(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0101D)
);

ninexnine_unit ninexnine_unit_980(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0201D)
);

assign C001D=c0001D+c0101D+c0201D;
assign A001D=(C001D>=0)?1:0;

assign P101D=A001D;

ninexnine_unit ninexnine_unit_981(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0002D)
);

ninexnine_unit ninexnine_unit_982(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0102D)
);

ninexnine_unit ninexnine_unit_983(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0202D)
);

assign C002D=c0002D+c0102D+c0202D;
assign A002D=(C002D>=0)?1:0;

assign P102D=A002D;

ninexnine_unit ninexnine_unit_984(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0003D)
);

ninexnine_unit ninexnine_unit_985(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0103D)
);

ninexnine_unit ninexnine_unit_986(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0203D)
);

assign C003D=c0003D+c0103D+c0203D;
assign A003D=(C003D>=0)?1:0;

assign P103D=A003D;

ninexnine_unit ninexnine_unit_987(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0004D)
);

ninexnine_unit ninexnine_unit_988(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0104D)
);

ninexnine_unit ninexnine_unit_989(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0204D)
);

assign C004D=c0004D+c0104D+c0204D;
assign A004D=(C004D>=0)?1:0;

assign P104D=A004D;

ninexnine_unit ninexnine_unit_990(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0010D)
);

ninexnine_unit ninexnine_unit_991(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0110D)
);

ninexnine_unit ninexnine_unit_992(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0210D)
);

assign C010D=c0010D+c0110D+c0210D;
assign A010D=(C010D>=0)?1:0;

assign P110D=A010D;

ninexnine_unit ninexnine_unit_993(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0011D)
);

ninexnine_unit ninexnine_unit_994(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0111D)
);

ninexnine_unit ninexnine_unit_995(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0211D)
);

assign C011D=c0011D+c0111D+c0211D;
assign A011D=(C011D>=0)?1:0;

assign P111D=A011D;

ninexnine_unit ninexnine_unit_996(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0012D)
);

ninexnine_unit ninexnine_unit_997(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0112D)
);

ninexnine_unit ninexnine_unit_998(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0212D)
);

assign C012D=c0012D+c0112D+c0212D;
assign A012D=(C012D>=0)?1:0;

assign P112D=A012D;

ninexnine_unit ninexnine_unit_999(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0013D)
);

ninexnine_unit ninexnine_unit_1000(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0113D)
);

ninexnine_unit ninexnine_unit_1001(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0213D)
);

assign C013D=c0013D+c0113D+c0213D;
assign A013D=(C013D>=0)?1:0;

assign P113D=A013D;

ninexnine_unit ninexnine_unit_1002(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0014D)
);

ninexnine_unit ninexnine_unit_1003(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0114D)
);

ninexnine_unit ninexnine_unit_1004(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0214D)
);

assign C014D=c0014D+c0114D+c0214D;
assign A014D=(C014D>=0)?1:0;

assign P114D=A014D;

ninexnine_unit ninexnine_unit_1005(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0020D)
);

ninexnine_unit ninexnine_unit_1006(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0120D)
);

ninexnine_unit ninexnine_unit_1007(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0220D)
);

assign C020D=c0020D+c0120D+c0220D;
assign A020D=(C020D>=0)?1:0;

assign P120D=A020D;

ninexnine_unit ninexnine_unit_1008(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0021D)
);

ninexnine_unit ninexnine_unit_1009(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0121D)
);

ninexnine_unit ninexnine_unit_1010(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0221D)
);

assign C021D=c0021D+c0121D+c0221D;
assign A021D=(C021D>=0)?1:0;

assign P121D=A021D;

ninexnine_unit ninexnine_unit_1011(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0022D)
);

ninexnine_unit ninexnine_unit_1012(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0122D)
);

ninexnine_unit ninexnine_unit_1013(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0222D)
);

assign C022D=c0022D+c0122D+c0222D;
assign A022D=(C022D>=0)?1:0;

assign P122D=A022D;

ninexnine_unit ninexnine_unit_1014(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0023D)
);

ninexnine_unit ninexnine_unit_1015(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0123D)
);

ninexnine_unit ninexnine_unit_1016(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0223D)
);

assign C023D=c0023D+c0123D+c0223D;
assign A023D=(C023D>=0)?1:0;

assign P123D=A023D;

ninexnine_unit ninexnine_unit_1017(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0024D)
);

ninexnine_unit ninexnine_unit_1018(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0124D)
);

ninexnine_unit ninexnine_unit_1019(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0224D)
);

assign C024D=c0024D+c0124D+c0224D;
assign A024D=(C024D>=0)?1:0;

assign P124D=A024D;

ninexnine_unit ninexnine_unit_1020(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0030D)
);

ninexnine_unit ninexnine_unit_1021(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0130D)
);

ninexnine_unit ninexnine_unit_1022(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0230D)
);

assign C030D=c0030D+c0130D+c0230D;
assign A030D=(C030D>=0)?1:0;

assign P130D=A030D;

ninexnine_unit ninexnine_unit_1023(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0031D)
);

ninexnine_unit ninexnine_unit_1024(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0131D)
);

ninexnine_unit ninexnine_unit_1025(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0231D)
);

assign C031D=c0031D+c0131D+c0231D;
assign A031D=(C031D>=0)?1:0;

assign P131D=A031D;

ninexnine_unit ninexnine_unit_1026(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0032D)
);

ninexnine_unit ninexnine_unit_1027(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0132D)
);

ninexnine_unit ninexnine_unit_1028(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0232D)
);

assign C032D=c0032D+c0132D+c0232D;
assign A032D=(C032D>=0)?1:0;

assign P132D=A032D;

ninexnine_unit ninexnine_unit_1029(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0033D)
);

ninexnine_unit ninexnine_unit_1030(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0133D)
);

ninexnine_unit ninexnine_unit_1031(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0233D)
);

assign C033D=c0033D+c0133D+c0233D;
assign A033D=(C033D>=0)?1:0;

assign P133D=A033D;

ninexnine_unit ninexnine_unit_1032(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0034D)
);

ninexnine_unit ninexnine_unit_1033(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0134D)
);

ninexnine_unit ninexnine_unit_1034(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0234D)
);

assign C034D=c0034D+c0134D+c0234D;
assign A034D=(C034D>=0)?1:0;

assign P134D=A034D;

ninexnine_unit ninexnine_unit_1035(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0040D)
);

ninexnine_unit ninexnine_unit_1036(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0140D)
);

ninexnine_unit ninexnine_unit_1037(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0240D)
);

assign C040D=c0040D+c0140D+c0240D;
assign A040D=(C040D>=0)?1:0;

assign P140D=A040D;

ninexnine_unit ninexnine_unit_1038(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0041D)
);

ninexnine_unit ninexnine_unit_1039(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0141D)
);

ninexnine_unit ninexnine_unit_1040(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0241D)
);

assign C041D=c0041D+c0141D+c0241D;
assign A041D=(C041D>=0)?1:0;

assign P141D=A041D;

ninexnine_unit ninexnine_unit_1041(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0042D)
);

ninexnine_unit ninexnine_unit_1042(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0142D)
);

ninexnine_unit ninexnine_unit_1043(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0242D)
);

assign C042D=c0042D+c0142D+c0242D;
assign A042D=(C042D>=0)?1:0;

assign P142D=A042D;

ninexnine_unit ninexnine_unit_1044(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0043D)
);

ninexnine_unit ninexnine_unit_1045(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0143D)
);

ninexnine_unit ninexnine_unit_1046(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0243D)
);

assign C043D=c0043D+c0143D+c0243D;
assign A043D=(C043D>=0)?1:0;

assign P143D=A043D;

ninexnine_unit ninexnine_unit_1047(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W0D000),
				.b1(W0D010),
				.b2(W0D020),
				.b3(W0D100),
				.b4(W0D110),
				.b5(W0D120),
				.b6(W0D200),
				.b7(W0D210),
				.b8(W0D220),
				.c(c0044D)
);

ninexnine_unit ninexnine_unit_1048(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W0D001),
				.b1(W0D011),
				.b2(W0D021),
				.b3(W0D101),
				.b4(W0D111),
				.b5(W0D121),
				.b6(W0D201),
				.b7(W0D211),
				.b8(W0D221),
				.c(c0144D)
);

ninexnine_unit ninexnine_unit_1049(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W0D002),
				.b1(W0D012),
				.b2(W0D022),
				.b3(W0D102),
				.b4(W0D112),
				.b5(W0D122),
				.b6(W0D202),
				.b7(W0D212),
				.b8(W0D222),
				.c(c0244D)
);

assign C044D=c0044D+c0144D+c0244D;
assign A044D=(C044D>=0)?1:0;

assign P144D=A044D;

ninexnine_unit ninexnine_unit_1050(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0000E)
);

ninexnine_unit ninexnine_unit_1051(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0100E)
);

ninexnine_unit ninexnine_unit_1052(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0200E)
);

assign C000E=c0000E+c0100E+c0200E;
assign A000E=(C000E>=0)?1:0;

assign P100E=A000E;

ninexnine_unit ninexnine_unit_1053(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0001E)
);

ninexnine_unit ninexnine_unit_1054(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0101E)
);

ninexnine_unit ninexnine_unit_1055(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0201E)
);

assign C001E=c0001E+c0101E+c0201E;
assign A001E=(C001E>=0)?1:0;

assign P101E=A001E;

ninexnine_unit ninexnine_unit_1056(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0002E)
);

ninexnine_unit ninexnine_unit_1057(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0102E)
);

ninexnine_unit ninexnine_unit_1058(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0202E)
);

assign C002E=c0002E+c0102E+c0202E;
assign A002E=(C002E>=0)?1:0;

assign P102E=A002E;

ninexnine_unit ninexnine_unit_1059(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0003E)
);

ninexnine_unit ninexnine_unit_1060(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0103E)
);

ninexnine_unit ninexnine_unit_1061(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0203E)
);

assign C003E=c0003E+c0103E+c0203E;
assign A003E=(C003E>=0)?1:0;

assign P103E=A003E;

ninexnine_unit ninexnine_unit_1062(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0004E)
);

ninexnine_unit ninexnine_unit_1063(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0104E)
);

ninexnine_unit ninexnine_unit_1064(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0204E)
);

assign C004E=c0004E+c0104E+c0204E;
assign A004E=(C004E>=0)?1:0;

assign P104E=A004E;

ninexnine_unit ninexnine_unit_1065(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0010E)
);

ninexnine_unit ninexnine_unit_1066(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0110E)
);

ninexnine_unit ninexnine_unit_1067(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0210E)
);

assign C010E=c0010E+c0110E+c0210E;
assign A010E=(C010E>=0)?1:0;

assign P110E=A010E;

ninexnine_unit ninexnine_unit_1068(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0011E)
);

ninexnine_unit ninexnine_unit_1069(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0111E)
);

ninexnine_unit ninexnine_unit_1070(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0211E)
);

assign C011E=c0011E+c0111E+c0211E;
assign A011E=(C011E>=0)?1:0;

assign P111E=A011E;

ninexnine_unit ninexnine_unit_1071(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0012E)
);

ninexnine_unit ninexnine_unit_1072(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0112E)
);

ninexnine_unit ninexnine_unit_1073(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0212E)
);

assign C012E=c0012E+c0112E+c0212E;
assign A012E=(C012E>=0)?1:0;

assign P112E=A012E;

ninexnine_unit ninexnine_unit_1074(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0013E)
);

ninexnine_unit ninexnine_unit_1075(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0113E)
);

ninexnine_unit ninexnine_unit_1076(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0213E)
);

assign C013E=c0013E+c0113E+c0213E;
assign A013E=(C013E>=0)?1:0;

assign P113E=A013E;

ninexnine_unit ninexnine_unit_1077(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0014E)
);

ninexnine_unit ninexnine_unit_1078(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0114E)
);

ninexnine_unit ninexnine_unit_1079(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0214E)
);

assign C014E=c0014E+c0114E+c0214E;
assign A014E=(C014E>=0)?1:0;

assign P114E=A014E;

ninexnine_unit ninexnine_unit_1080(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0020E)
);

ninexnine_unit ninexnine_unit_1081(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0120E)
);

ninexnine_unit ninexnine_unit_1082(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0220E)
);

assign C020E=c0020E+c0120E+c0220E;
assign A020E=(C020E>=0)?1:0;

assign P120E=A020E;

ninexnine_unit ninexnine_unit_1083(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0021E)
);

ninexnine_unit ninexnine_unit_1084(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0121E)
);

ninexnine_unit ninexnine_unit_1085(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0221E)
);

assign C021E=c0021E+c0121E+c0221E;
assign A021E=(C021E>=0)?1:0;

assign P121E=A021E;

ninexnine_unit ninexnine_unit_1086(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0022E)
);

ninexnine_unit ninexnine_unit_1087(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0122E)
);

ninexnine_unit ninexnine_unit_1088(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0222E)
);

assign C022E=c0022E+c0122E+c0222E;
assign A022E=(C022E>=0)?1:0;

assign P122E=A022E;

ninexnine_unit ninexnine_unit_1089(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0023E)
);

ninexnine_unit ninexnine_unit_1090(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0123E)
);

ninexnine_unit ninexnine_unit_1091(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0223E)
);

assign C023E=c0023E+c0123E+c0223E;
assign A023E=(C023E>=0)?1:0;

assign P123E=A023E;

ninexnine_unit ninexnine_unit_1092(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0024E)
);

ninexnine_unit ninexnine_unit_1093(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0124E)
);

ninexnine_unit ninexnine_unit_1094(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0224E)
);

assign C024E=c0024E+c0124E+c0224E;
assign A024E=(C024E>=0)?1:0;

assign P124E=A024E;

ninexnine_unit ninexnine_unit_1095(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0030E)
);

ninexnine_unit ninexnine_unit_1096(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0130E)
);

ninexnine_unit ninexnine_unit_1097(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0230E)
);

assign C030E=c0030E+c0130E+c0230E;
assign A030E=(C030E>=0)?1:0;

assign P130E=A030E;

ninexnine_unit ninexnine_unit_1098(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0031E)
);

ninexnine_unit ninexnine_unit_1099(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0131E)
);

ninexnine_unit ninexnine_unit_1100(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0231E)
);

assign C031E=c0031E+c0131E+c0231E;
assign A031E=(C031E>=0)?1:0;

assign P131E=A031E;

ninexnine_unit ninexnine_unit_1101(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0032E)
);

ninexnine_unit ninexnine_unit_1102(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0132E)
);

ninexnine_unit ninexnine_unit_1103(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0232E)
);

assign C032E=c0032E+c0132E+c0232E;
assign A032E=(C032E>=0)?1:0;

assign P132E=A032E;

ninexnine_unit ninexnine_unit_1104(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0033E)
);

ninexnine_unit ninexnine_unit_1105(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0133E)
);

ninexnine_unit ninexnine_unit_1106(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0233E)
);

assign C033E=c0033E+c0133E+c0233E;
assign A033E=(C033E>=0)?1:0;

assign P133E=A033E;

ninexnine_unit ninexnine_unit_1107(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0034E)
);

ninexnine_unit ninexnine_unit_1108(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0134E)
);

ninexnine_unit ninexnine_unit_1109(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0234E)
);

assign C034E=c0034E+c0134E+c0234E;
assign A034E=(C034E>=0)?1:0;

assign P134E=A034E;

ninexnine_unit ninexnine_unit_1110(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0040E)
);

ninexnine_unit ninexnine_unit_1111(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0140E)
);

ninexnine_unit ninexnine_unit_1112(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0240E)
);

assign C040E=c0040E+c0140E+c0240E;
assign A040E=(C040E>=0)?1:0;

assign P140E=A040E;

ninexnine_unit ninexnine_unit_1113(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0041E)
);

ninexnine_unit ninexnine_unit_1114(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0141E)
);

ninexnine_unit ninexnine_unit_1115(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0241E)
);

assign C041E=c0041E+c0141E+c0241E;
assign A041E=(C041E>=0)?1:0;

assign P141E=A041E;

ninexnine_unit ninexnine_unit_1116(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0042E)
);

ninexnine_unit ninexnine_unit_1117(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0142E)
);

ninexnine_unit ninexnine_unit_1118(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0242E)
);

assign C042E=c0042E+c0142E+c0242E;
assign A042E=(C042E>=0)?1:0;

assign P142E=A042E;

ninexnine_unit ninexnine_unit_1119(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0043E)
);

ninexnine_unit ninexnine_unit_1120(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0143E)
);

ninexnine_unit ninexnine_unit_1121(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0243E)
);

assign C043E=c0043E+c0143E+c0243E;
assign A043E=(C043E>=0)?1:0;

assign P143E=A043E;

ninexnine_unit ninexnine_unit_1122(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W0E000),
				.b1(W0E010),
				.b2(W0E020),
				.b3(W0E100),
				.b4(W0E110),
				.b5(W0E120),
				.b6(W0E200),
				.b7(W0E210),
				.b8(W0E220),
				.c(c0044E)
);

ninexnine_unit ninexnine_unit_1123(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W0E001),
				.b1(W0E011),
				.b2(W0E021),
				.b3(W0E101),
				.b4(W0E111),
				.b5(W0E121),
				.b6(W0E201),
				.b7(W0E211),
				.b8(W0E221),
				.c(c0144E)
);

ninexnine_unit ninexnine_unit_1124(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W0E002),
				.b1(W0E012),
				.b2(W0E022),
				.b3(W0E102),
				.b4(W0E112),
				.b5(W0E122),
				.b6(W0E202),
				.b7(W0E212),
				.b8(W0E222),
				.c(c0244E)
);

assign C044E=c0044E+c0144E+c0244E;
assign A044E=(C044E>=0)?1:0;

assign P144E=A044E;

ninexnine_unit ninexnine_unit_1125(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0000F)
);

ninexnine_unit ninexnine_unit_1126(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0100F)
);

ninexnine_unit ninexnine_unit_1127(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0200F)
);

assign C000F=c0000F+c0100F+c0200F;
assign A000F=(C000F>=0)?1:0;

assign P100F=A000F;

ninexnine_unit ninexnine_unit_1128(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0001F)
);

ninexnine_unit ninexnine_unit_1129(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0101F)
);

ninexnine_unit ninexnine_unit_1130(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0201F)
);

assign C001F=c0001F+c0101F+c0201F;
assign A001F=(C001F>=0)?1:0;

assign P101F=A001F;

ninexnine_unit ninexnine_unit_1131(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0002F)
);

ninexnine_unit ninexnine_unit_1132(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0102F)
);

ninexnine_unit ninexnine_unit_1133(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0202F)
);

assign C002F=c0002F+c0102F+c0202F;
assign A002F=(C002F>=0)?1:0;

assign P102F=A002F;

ninexnine_unit ninexnine_unit_1134(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0003F)
);

ninexnine_unit ninexnine_unit_1135(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0103F)
);

ninexnine_unit ninexnine_unit_1136(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0203F)
);

assign C003F=c0003F+c0103F+c0203F;
assign A003F=(C003F>=0)?1:0;

assign P103F=A003F;

ninexnine_unit ninexnine_unit_1137(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0004F)
);

ninexnine_unit ninexnine_unit_1138(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0104F)
);

ninexnine_unit ninexnine_unit_1139(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0204F)
);

assign C004F=c0004F+c0104F+c0204F;
assign A004F=(C004F>=0)?1:0;

assign P104F=A004F;

ninexnine_unit ninexnine_unit_1140(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0010F)
);

ninexnine_unit ninexnine_unit_1141(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0110F)
);

ninexnine_unit ninexnine_unit_1142(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0210F)
);

assign C010F=c0010F+c0110F+c0210F;
assign A010F=(C010F>=0)?1:0;

assign P110F=A010F;

ninexnine_unit ninexnine_unit_1143(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0011F)
);

ninexnine_unit ninexnine_unit_1144(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0111F)
);

ninexnine_unit ninexnine_unit_1145(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0211F)
);

assign C011F=c0011F+c0111F+c0211F;
assign A011F=(C011F>=0)?1:0;

assign P111F=A011F;

ninexnine_unit ninexnine_unit_1146(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0012F)
);

ninexnine_unit ninexnine_unit_1147(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0112F)
);

ninexnine_unit ninexnine_unit_1148(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0212F)
);

assign C012F=c0012F+c0112F+c0212F;
assign A012F=(C012F>=0)?1:0;

assign P112F=A012F;

ninexnine_unit ninexnine_unit_1149(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0013F)
);

ninexnine_unit ninexnine_unit_1150(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0113F)
);

ninexnine_unit ninexnine_unit_1151(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0213F)
);

assign C013F=c0013F+c0113F+c0213F;
assign A013F=(C013F>=0)?1:0;

assign P113F=A013F;

ninexnine_unit ninexnine_unit_1152(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0014F)
);

ninexnine_unit ninexnine_unit_1153(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0114F)
);

ninexnine_unit ninexnine_unit_1154(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0214F)
);

assign C014F=c0014F+c0114F+c0214F;
assign A014F=(C014F>=0)?1:0;

assign P114F=A014F;

ninexnine_unit ninexnine_unit_1155(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0020F)
);

ninexnine_unit ninexnine_unit_1156(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0120F)
);

ninexnine_unit ninexnine_unit_1157(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0220F)
);

assign C020F=c0020F+c0120F+c0220F;
assign A020F=(C020F>=0)?1:0;

assign P120F=A020F;

ninexnine_unit ninexnine_unit_1158(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0021F)
);

ninexnine_unit ninexnine_unit_1159(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0121F)
);

ninexnine_unit ninexnine_unit_1160(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0221F)
);

assign C021F=c0021F+c0121F+c0221F;
assign A021F=(C021F>=0)?1:0;

assign P121F=A021F;

ninexnine_unit ninexnine_unit_1161(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0022F)
);

ninexnine_unit ninexnine_unit_1162(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0122F)
);

ninexnine_unit ninexnine_unit_1163(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0222F)
);

assign C022F=c0022F+c0122F+c0222F;
assign A022F=(C022F>=0)?1:0;

assign P122F=A022F;

ninexnine_unit ninexnine_unit_1164(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0023F)
);

ninexnine_unit ninexnine_unit_1165(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0123F)
);

ninexnine_unit ninexnine_unit_1166(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0223F)
);

assign C023F=c0023F+c0123F+c0223F;
assign A023F=(C023F>=0)?1:0;

assign P123F=A023F;

ninexnine_unit ninexnine_unit_1167(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0024F)
);

ninexnine_unit ninexnine_unit_1168(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0124F)
);

ninexnine_unit ninexnine_unit_1169(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0224F)
);

assign C024F=c0024F+c0124F+c0224F;
assign A024F=(C024F>=0)?1:0;

assign P124F=A024F;

ninexnine_unit ninexnine_unit_1170(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0030F)
);

ninexnine_unit ninexnine_unit_1171(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0130F)
);

ninexnine_unit ninexnine_unit_1172(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0230F)
);

assign C030F=c0030F+c0130F+c0230F;
assign A030F=(C030F>=0)?1:0;

assign P130F=A030F;

ninexnine_unit ninexnine_unit_1173(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0031F)
);

ninexnine_unit ninexnine_unit_1174(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0131F)
);

ninexnine_unit ninexnine_unit_1175(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0231F)
);

assign C031F=c0031F+c0131F+c0231F;
assign A031F=(C031F>=0)?1:0;

assign P131F=A031F;

ninexnine_unit ninexnine_unit_1176(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0032F)
);

ninexnine_unit ninexnine_unit_1177(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0132F)
);

ninexnine_unit ninexnine_unit_1178(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0232F)
);

assign C032F=c0032F+c0132F+c0232F;
assign A032F=(C032F>=0)?1:0;

assign P132F=A032F;

ninexnine_unit ninexnine_unit_1179(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0033F)
);

ninexnine_unit ninexnine_unit_1180(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0133F)
);

ninexnine_unit ninexnine_unit_1181(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0233F)
);

assign C033F=c0033F+c0133F+c0233F;
assign A033F=(C033F>=0)?1:0;

assign P133F=A033F;

ninexnine_unit ninexnine_unit_1182(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0034F)
);

ninexnine_unit ninexnine_unit_1183(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0134F)
);

ninexnine_unit ninexnine_unit_1184(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0234F)
);

assign C034F=c0034F+c0134F+c0234F;
assign A034F=(C034F>=0)?1:0;

assign P134F=A034F;

ninexnine_unit ninexnine_unit_1185(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0040F)
);

ninexnine_unit ninexnine_unit_1186(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0140F)
);

ninexnine_unit ninexnine_unit_1187(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0240F)
);

assign C040F=c0040F+c0140F+c0240F;
assign A040F=(C040F>=0)?1:0;

assign P140F=A040F;

ninexnine_unit ninexnine_unit_1188(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0041F)
);

ninexnine_unit ninexnine_unit_1189(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0141F)
);

ninexnine_unit ninexnine_unit_1190(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0241F)
);

assign C041F=c0041F+c0141F+c0241F;
assign A041F=(C041F>=0)?1:0;

assign P141F=A041F;

ninexnine_unit ninexnine_unit_1191(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0042F)
);

ninexnine_unit ninexnine_unit_1192(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0142F)
);

ninexnine_unit ninexnine_unit_1193(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0242F)
);

assign C042F=c0042F+c0142F+c0242F;
assign A042F=(C042F>=0)?1:0;

assign P142F=A042F;

ninexnine_unit ninexnine_unit_1194(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0043F)
);

ninexnine_unit ninexnine_unit_1195(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0143F)
);

ninexnine_unit ninexnine_unit_1196(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0243F)
);

assign C043F=c0043F+c0143F+c0243F;
assign A043F=(C043F>=0)?1:0;

assign P143F=A043F;

ninexnine_unit ninexnine_unit_1197(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W0F000),
				.b1(W0F010),
				.b2(W0F020),
				.b3(W0F100),
				.b4(W0F110),
				.b5(W0F120),
				.b6(W0F200),
				.b7(W0F210),
				.b8(W0F220),
				.c(c0044F)
);

ninexnine_unit ninexnine_unit_1198(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W0F001),
				.b1(W0F011),
				.b2(W0F021),
				.b3(W0F101),
				.b4(W0F111),
				.b5(W0F121),
				.b6(W0F201),
				.b7(W0F211),
				.b8(W0F221),
				.c(c0144F)
);

ninexnine_unit ninexnine_unit_1199(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W0F002),
				.b1(W0F012),
				.b2(W0F022),
				.b3(W0F102),
				.b4(W0F112),
				.b5(W0F122),
				.b6(W0F202),
				.b7(W0F212),
				.b8(W0F222),
				.c(c0244F)
);

assign C044F=c0044F+c0144F+c0244F;
assign A044F=(C044F>=0)?1:0;

assign P144F=A044F;

//layer2 done, begain next layer
wire P2000;
wire P2010;
wire P2020;
wire P2100;
wire P2110;
wire P2120;
wire P2200;
wire P2210;
wire P2220;
wire P2001;
wire P2011;
wire P2021;
wire P2101;
wire P2111;
wire P2121;
wire P2201;
wire P2211;
wire P2221;
wire P2002;
wire P2012;
wire P2022;
wire P2102;
wire P2112;
wire P2122;
wire P2202;
wire P2212;
wire P2222;
wire P2003;
wire P2013;
wire P2023;
wire P2103;
wire P2113;
wire P2123;
wire P2203;
wire P2213;
wire P2223;
wire P2004;
wire P2014;
wire P2024;
wire P2104;
wire P2114;
wire P2124;
wire P2204;
wire P2214;
wire P2224;
wire P2005;
wire P2015;
wire P2025;
wire P2105;
wire P2115;
wire P2125;
wire P2205;
wire P2215;
wire P2225;
wire P2006;
wire P2016;
wire P2026;
wire P2106;
wire P2116;
wire P2126;
wire P2206;
wire P2216;
wire P2226;
wire P2007;
wire P2017;
wire P2027;
wire P2107;
wire P2117;
wire P2127;
wire P2207;
wire P2217;
wire P2227;
wire P2008;
wire P2018;
wire P2028;
wire P2108;
wire P2118;
wire P2128;
wire P2208;
wire P2218;
wire P2228;
wire P2009;
wire P2019;
wire P2029;
wire P2109;
wire P2119;
wire P2129;
wire P2209;
wire P2219;
wire P2229;
wire P200A;
wire P201A;
wire P202A;
wire P210A;
wire P211A;
wire P212A;
wire P220A;
wire P221A;
wire P222A;
wire P200B;
wire P201B;
wire P202B;
wire P210B;
wire P211B;
wire P212B;
wire P220B;
wire P221B;
wire P222B;
wire P200C;
wire P201C;
wire P202C;
wire P210C;
wire P211C;
wire P212C;
wire P220C;
wire P221C;
wire P222C;
wire P200D;
wire P201D;
wire P202D;
wire P210D;
wire P211D;
wire P212D;
wire P220D;
wire P221D;
wire P222D;
wire P200E;
wire P201E;
wire P202E;
wire P210E;
wire P211E;
wire P212E;
wire P220E;
wire P221E;
wire P222E;
wire P200F;
wire P201F;
wire P202F;
wire P210F;
wire P211F;
wire P212F;
wire P220F;
wire P221F;
wire P222F;
wire P200G;
wire P201G;
wire P202G;
wire P210G;
wire P211G;
wire P212G;
wire P220G;
wire P221G;
wire P222G;
wire P200H;
wire P201H;
wire P202H;
wire P210H;
wire P211H;
wire P212H;
wire P220H;
wire P221H;
wire P222H;
wire P200I;
wire P201I;
wire P202I;
wire P210I;
wire P211I;
wire P212I;
wire P220I;
wire P221I;
wire P222I;
wire P200J;
wire P201J;
wire P202J;
wire P210J;
wire P211J;
wire P212J;
wire P220J;
wire P221J;
wire P222J;
wire P200K;
wire P201K;
wire P202K;
wire P210K;
wire P211K;
wire P212K;
wire P220K;
wire P221K;
wire P222K;
wire P200L;
wire P201L;
wire P202L;
wire P210L;
wire P211L;
wire P212L;
wire P220L;
wire P221L;
wire P222L;
wire P200M;
wire P201M;
wire P202M;
wire P210M;
wire P211M;
wire P212M;
wire P220M;
wire P221M;
wire P222M;
wire W10000,W10010,W10020,W10100,W10110,W10120,W10200,W10210,W10220;
wire W10001,W10011,W10021,W10101,W10111,W10121,W10201,W10211,W10221;
wire W10002,W10012,W10022,W10102,W10112,W10122,W10202,W10212,W10222;
wire W10003,W10013,W10023,W10103,W10113,W10123,W10203,W10213,W10223;
wire W10004,W10014,W10024,W10104,W10114,W10124,W10204,W10214,W10224;
wire W10005,W10015,W10025,W10105,W10115,W10125,W10205,W10215,W10225;
wire W10006,W10016,W10026,W10106,W10116,W10126,W10206,W10216,W10226;
wire W10007,W10017,W10027,W10107,W10117,W10127,W10207,W10217,W10227;
wire W10008,W10018,W10028,W10108,W10118,W10128,W10208,W10218,W10228;
wire W10009,W10019,W10029,W10109,W10119,W10129,W10209,W10219,W10229;
wire W1000A,W1001A,W1002A,W1010A,W1011A,W1012A,W1020A,W1021A,W1022A;
wire W1000B,W1001B,W1002B,W1010B,W1011B,W1012B,W1020B,W1021B,W1022B;
wire W1000C,W1001C,W1002C,W1010C,W1011C,W1012C,W1020C,W1021C,W1022C;
wire W1000D,W1001D,W1002D,W1010D,W1011D,W1012D,W1020D,W1021D,W1022D;
wire W1000E,W1001E,W1002E,W1010E,W1011E,W1012E,W1020E,W1021E,W1022E;
wire W1000F,W1001F,W1002F,W1010F,W1011F,W1012F,W1020F,W1021F,W1022F;
wire W11000,W11010,W11020,W11100,W11110,W11120,W11200,W11210,W11220;
wire W11001,W11011,W11021,W11101,W11111,W11121,W11201,W11211,W11221;
wire W11002,W11012,W11022,W11102,W11112,W11122,W11202,W11212,W11222;
wire W11003,W11013,W11023,W11103,W11113,W11123,W11203,W11213,W11223;
wire W11004,W11014,W11024,W11104,W11114,W11124,W11204,W11214,W11224;
wire W11005,W11015,W11025,W11105,W11115,W11125,W11205,W11215,W11225;
wire W11006,W11016,W11026,W11106,W11116,W11126,W11206,W11216,W11226;
wire W11007,W11017,W11027,W11107,W11117,W11127,W11207,W11217,W11227;
wire W11008,W11018,W11028,W11108,W11118,W11128,W11208,W11218,W11228;
wire W11009,W11019,W11029,W11109,W11119,W11129,W11209,W11219,W11229;
wire W1100A,W1101A,W1102A,W1110A,W1111A,W1112A,W1120A,W1121A,W1122A;
wire W1100B,W1101B,W1102B,W1110B,W1111B,W1112B,W1120B,W1121B,W1122B;
wire W1100C,W1101C,W1102C,W1110C,W1111C,W1112C,W1120C,W1121C,W1122C;
wire W1100D,W1101D,W1102D,W1110D,W1111D,W1112D,W1120D,W1121D,W1122D;
wire W1100E,W1101E,W1102E,W1110E,W1111E,W1112E,W1120E,W1121E,W1122E;
wire W1100F,W1101F,W1102F,W1110F,W1111F,W1112F,W1120F,W1121F,W1122F;
wire W12000,W12010,W12020,W12100,W12110,W12120,W12200,W12210,W12220;
wire W12001,W12011,W12021,W12101,W12111,W12121,W12201,W12211,W12221;
wire W12002,W12012,W12022,W12102,W12112,W12122,W12202,W12212,W12222;
wire W12003,W12013,W12023,W12103,W12113,W12123,W12203,W12213,W12223;
wire W12004,W12014,W12024,W12104,W12114,W12124,W12204,W12214,W12224;
wire W12005,W12015,W12025,W12105,W12115,W12125,W12205,W12215,W12225;
wire W12006,W12016,W12026,W12106,W12116,W12126,W12206,W12216,W12226;
wire W12007,W12017,W12027,W12107,W12117,W12127,W12207,W12217,W12227;
wire W12008,W12018,W12028,W12108,W12118,W12128,W12208,W12218,W12228;
wire W12009,W12019,W12029,W12109,W12119,W12129,W12209,W12219,W12229;
wire W1200A,W1201A,W1202A,W1210A,W1211A,W1212A,W1220A,W1221A,W1222A;
wire W1200B,W1201B,W1202B,W1210B,W1211B,W1212B,W1220B,W1221B,W1222B;
wire W1200C,W1201C,W1202C,W1210C,W1211C,W1212C,W1220C,W1221C,W1222C;
wire W1200D,W1201D,W1202D,W1210D,W1211D,W1212D,W1220D,W1221D,W1222D;
wire W1200E,W1201E,W1202E,W1210E,W1211E,W1212E,W1220E,W1221E,W1222E;
wire W1200F,W1201F,W1202F,W1210F,W1211F,W1212F,W1220F,W1221F,W1222F;
wire W13000,W13010,W13020,W13100,W13110,W13120,W13200,W13210,W13220;
wire W13001,W13011,W13021,W13101,W13111,W13121,W13201,W13211,W13221;
wire W13002,W13012,W13022,W13102,W13112,W13122,W13202,W13212,W13222;
wire W13003,W13013,W13023,W13103,W13113,W13123,W13203,W13213,W13223;
wire W13004,W13014,W13024,W13104,W13114,W13124,W13204,W13214,W13224;
wire W13005,W13015,W13025,W13105,W13115,W13125,W13205,W13215,W13225;
wire W13006,W13016,W13026,W13106,W13116,W13126,W13206,W13216,W13226;
wire W13007,W13017,W13027,W13107,W13117,W13127,W13207,W13217,W13227;
wire W13008,W13018,W13028,W13108,W13118,W13128,W13208,W13218,W13228;
wire W13009,W13019,W13029,W13109,W13119,W13129,W13209,W13219,W13229;
wire W1300A,W1301A,W1302A,W1310A,W1311A,W1312A,W1320A,W1321A,W1322A;
wire W1300B,W1301B,W1302B,W1310B,W1311B,W1312B,W1320B,W1321B,W1322B;
wire W1300C,W1301C,W1302C,W1310C,W1311C,W1312C,W1320C,W1321C,W1322C;
wire W1300D,W1301D,W1302D,W1310D,W1311D,W1312D,W1320D,W1321D,W1322D;
wire W1300E,W1301E,W1302E,W1310E,W1311E,W1312E,W1320E,W1321E,W1322E;
wire W1300F,W1301F,W1302F,W1310F,W1311F,W1312F,W1320F,W1321F,W1322F;
wire W14000,W14010,W14020,W14100,W14110,W14120,W14200,W14210,W14220;
wire W14001,W14011,W14021,W14101,W14111,W14121,W14201,W14211,W14221;
wire W14002,W14012,W14022,W14102,W14112,W14122,W14202,W14212,W14222;
wire W14003,W14013,W14023,W14103,W14113,W14123,W14203,W14213,W14223;
wire W14004,W14014,W14024,W14104,W14114,W14124,W14204,W14214,W14224;
wire W14005,W14015,W14025,W14105,W14115,W14125,W14205,W14215,W14225;
wire W14006,W14016,W14026,W14106,W14116,W14126,W14206,W14216,W14226;
wire W14007,W14017,W14027,W14107,W14117,W14127,W14207,W14217,W14227;
wire W14008,W14018,W14028,W14108,W14118,W14128,W14208,W14218,W14228;
wire W14009,W14019,W14029,W14109,W14119,W14129,W14209,W14219,W14229;
wire W1400A,W1401A,W1402A,W1410A,W1411A,W1412A,W1420A,W1421A,W1422A;
wire W1400B,W1401B,W1402B,W1410B,W1411B,W1412B,W1420B,W1421B,W1422B;
wire W1400C,W1401C,W1402C,W1410C,W1411C,W1412C,W1420C,W1421C,W1422C;
wire W1400D,W1401D,W1402D,W1410D,W1411D,W1412D,W1420D,W1421D,W1422D;
wire W1400E,W1401E,W1402E,W1410E,W1411E,W1412E,W1420E,W1421E,W1422E;
wire W1400F,W1401F,W1402F,W1410F,W1411F,W1412F,W1420F,W1421F,W1422F;
wire W15000,W15010,W15020,W15100,W15110,W15120,W15200,W15210,W15220;
wire W15001,W15011,W15021,W15101,W15111,W15121,W15201,W15211,W15221;
wire W15002,W15012,W15022,W15102,W15112,W15122,W15202,W15212,W15222;
wire W15003,W15013,W15023,W15103,W15113,W15123,W15203,W15213,W15223;
wire W15004,W15014,W15024,W15104,W15114,W15124,W15204,W15214,W15224;
wire W15005,W15015,W15025,W15105,W15115,W15125,W15205,W15215,W15225;
wire W15006,W15016,W15026,W15106,W15116,W15126,W15206,W15216,W15226;
wire W15007,W15017,W15027,W15107,W15117,W15127,W15207,W15217,W15227;
wire W15008,W15018,W15028,W15108,W15118,W15128,W15208,W15218,W15228;
wire W15009,W15019,W15029,W15109,W15119,W15129,W15209,W15219,W15229;
wire W1500A,W1501A,W1502A,W1510A,W1511A,W1512A,W1520A,W1521A,W1522A;
wire W1500B,W1501B,W1502B,W1510B,W1511B,W1512B,W1520B,W1521B,W1522B;
wire W1500C,W1501C,W1502C,W1510C,W1511C,W1512C,W1520C,W1521C,W1522C;
wire W1500D,W1501D,W1502D,W1510D,W1511D,W1512D,W1520D,W1521D,W1522D;
wire W1500E,W1501E,W1502E,W1510E,W1511E,W1512E,W1520E,W1521E,W1522E;
wire W1500F,W1501F,W1502F,W1510F,W1511F,W1512F,W1520F,W1521F,W1522F;
wire W16000,W16010,W16020,W16100,W16110,W16120,W16200,W16210,W16220;
wire W16001,W16011,W16021,W16101,W16111,W16121,W16201,W16211,W16221;
wire W16002,W16012,W16022,W16102,W16112,W16122,W16202,W16212,W16222;
wire W16003,W16013,W16023,W16103,W16113,W16123,W16203,W16213,W16223;
wire W16004,W16014,W16024,W16104,W16114,W16124,W16204,W16214,W16224;
wire W16005,W16015,W16025,W16105,W16115,W16125,W16205,W16215,W16225;
wire W16006,W16016,W16026,W16106,W16116,W16126,W16206,W16216,W16226;
wire W16007,W16017,W16027,W16107,W16117,W16127,W16207,W16217,W16227;
wire W16008,W16018,W16028,W16108,W16118,W16128,W16208,W16218,W16228;
wire W16009,W16019,W16029,W16109,W16119,W16129,W16209,W16219,W16229;
wire W1600A,W1601A,W1602A,W1610A,W1611A,W1612A,W1620A,W1621A,W1622A;
wire W1600B,W1601B,W1602B,W1610B,W1611B,W1612B,W1620B,W1621B,W1622B;
wire W1600C,W1601C,W1602C,W1610C,W1611C,W1612C,W1620C,W1621C,W1622C;
wire W1600D,W1601D,W1602D,W1610D,W1611D,W1612D,W1620D,W1621D,W1622D;
wire W1600E,W1601E,W1602E,W1610E,W1611E,W1612E,W1620E,W1621E,W1622E;
wire W1600F,W1601F,W1602F,W1610F,W1611F,W1612F,W1620F,W1621F,W1622F;
wire W17000,W17010,W17020,W17100,W17110,W17120,W17200,W17210,W17220;
wire W17001,W17011,W17021,W17101,W17111,W17121,W17201,W17211,W17221;
wire W17002,W17012,W17022,W17102,W17112,W17122,W17202,W17212,W17222;
wire W17003,W17013,W17023,W17103,W17113,W17123,W17203,W17213,W17223;
wire W17004,W17014,W17024,W17104,W17114,W17124,W17204,W17214,W17224;
wire W17005,W17015,W17025,W17105,W17115,W17125,W17205,W17215,W17225;
wire W17006,W17016,W17026,W17106,W17116,W17126,W17206,W17216,W17226;
wire W17007,W17017,W17027,W17107,W17117,W17127,W17207,W17217,W17227;
wire W17008,W17018,W17028,W17108,W17118,W17128,W17208,W17218,W17228;
wire W17009,W17019,W17029,W17109,W17119,W17129,W17209,W17219,W17229;
wire W1700A,W1701A,W1702A,W1710A,W1711A,W1712A,W1720A,W1721A,W1722A;
wire W1700B,W1701B,W1702B,W1710B,W1711B,W1712B,W1720B,W1721B,W1722B;
wire W1700C,W1701C,W1702C,W1710C,W1711C,W1712C,W1720C,W1721C,W1722C;
wire W1700D,W1701D,W1702D,W1710D,W1711D,W1712D,W1720D,W1721D,W1722D;
wire W1700E,W1701E,W1702E,W1710E,W1711E,W1712E,W1720E,W1721E,W1722E;
wire W1700F,W1701F,W1702F,W1710F,W1711F,W1712F,W1720F,W1721F,W1722F;
wire W18000,W18010,W18020,W18100,W18110,W18120,W18200,W18210,W18220;
wire W18001,W18011,W18021,W18101,W18111,W18121,W18201,W18211,W18221;
wire W18002,W18012,W18022,W18102,W18112,W18122,W18202,W18212,W18222;
wire W18003,W18013,W18023,W18103,W18113,W18123,W18203,W18213,W18223;
wire W18004,W18014,W18024,W18104,W18114,W18124,W18204,W18214,W18224;
wire W18005,W18015,W18025,W18105,W18115,W18125,W18205,W18215,W18225;
wire W18006,W18016,W18026,W18106,W18116,W18126,W18206,W18216,W18226;
wire W18007,W18017,W18027,W18107,W18117,W18127,W18207,W18217,W18227;
wire W18008,W18018,W18028,W18108,W18118,W18128,W18208,W18218,W18228;
wire W18009,W18019,W18029,W18109,W18119,W18129,W18209,W18219,W18229;
wire W1800A,W1801A,W1802A,W1810A,W1811A,W1812A,W1820A,W1821A,W1822A;
wire W1800B,W1801B,W1802B,W1810B,W1811B,W1812B,W1820B,W1821B,W1822B;
wire W1800C,W1801C,W1802C,W1810C,W1811C,W1812C,W1820C,W1821C,W1822C;
wire W1800D,W1801D,W1802D,W1810D,W1811D,W1812D,W1820D,W1821D,W1822D;
wire W1800E,W1801E,W1802E,W1810E,W1811E,W1812E,W1820E,W1821E,W1822E;
wire W1800F,W1801F,W1802F,W1810F,W1811F,W1812F,W1820F,W1821F,W1822F;
wire W19000,W19010,W19020,W19100,W19110,W19120,W19200,W19210,W19220;
wire W19001,W19011,W19021,W19101,W19111,W19121,W19201,W19211,W19221;
wire W19002,W19012,W19022,W19102,W19112,W19122,W19202,W19212,W19222;
wire W19003,W19013,W19023,W19103,W19113,W19123,W19203,W19213,W19223;
wire W19004,W19014,W19024,W19104,W19114,W19124,W19204,W19214,W19224;
wire W19005,W19015,W19025,W19105,W19115,W19125,W19205,W19215,W19225;
wire W19006,W19016,W19026,W19106,W19116,W19126,W19206,W19216,W19226;
wire W19007,W19017,W19027,W19107,W19117,W19127,W19207,W19217,W19227;
wire W19008,W19018,W19028,W19108,W19118,W19128,W19208,W19218,W19228;
wire W19009,W19019,W19029,W19109,W19119,W19129,W19209,W19219,W19229;
wire W1900A,W1901A,W1902A,W1910A,W1911A,W1912A,W1920A,W1921A,W1922A;
wire W1900B,W1901B,W1902B,W1910B,W1911B,W1912B,W1920B,W1921B,W1922B;
wire W1900C,W1901C,W1902C,W1910C,W1911C,W1912C,W1920C,W1921C,W1922C;
wire W1900D,W1901D,W1902D,W1910D,W1911D,W1912D,W1920D,W1921D,W1922D;
wire W1900E,W1901E,W1902E,W1910E,W1911E,W1912E,W1920E,W1921E,W1922E;
wire W1900F,W1901F,W1902F,W1910F,W1911F,W1912F,W1920F,W1921F,W1922F;
wire W1A000,W1A010,W1A020,W1A100,W1A110,W1A120,W1A200,W1A210,W1A220;
wire W1A001,W1A011,W1A021,W1A101,W1A111,W1A121,W1A201,W1A211,W1A221;
wire W1A002,W1A012,W1A022,W1A102,W1A112,W1A122,W1A202,W1A212,W1A222;
wire W1A003,W1A013,W1A023,W1A103,W1A113,W1A123,W1A203,W1A213,W1A223;
wire W1A004,W1A014,W1A024,W1A104,W1A114,W1A124,W1A204,W1A214,W1A224;
wire W1A005,W1A015,W1A025,W1A105,W1A115,W1A125,W1A205,W1A215,W1A225;
wire W1A006,W1A016,W1A026,W1A106,W1A116,W1A126,W1A206,W1A216,W1A226;
wire W1A007,W1A017,W1A027,W1A107,W1A117,W1A127,W1A207,W1A217,W1A227;
wire W1A008,W1A018,W1A028,W1A108,W1A118,W1A128,W1A208,W1A218,W1A228;
wire W1A009,W1A019,W1A029,W1A109,W1A119,W1A129,W1A209,W1A219,W1A229;
wire W1A00A,W1A01A,W1A02A,W1A10A,W1A11A,W1A12A,W1A20A,W1A21A,W1A22A;
wire W1A00B,W1A01B,W1A02B,W1A10B,W1A11B,W1A12B,W1A20B,W1A21B,W1A22B;
wire W1A00C,W1A01C,W1A02C,W1A10C,W1A11C,W1A12C,W1A20C,W1A21C,W1A22C;
wire W1A00D,W1A01D,W1A02D,W1A10D,W1A11D,W1A12D,W1A20D,W1A21D,W1A22D;
wire W1A00E,W1A01E,W1A02E,W1A10E,W1A11E,W1A12E,W1A20E,W1A21E,W1A22E;
wire W1A00F,W1A01F,W1A02F,W1A10F,W1A11F,W1A12F,W1A20F,W1A21F,W1A22F;
wire W1B000,W1B010,W1B020,W1B100,W1B110,W1B120,W1B200,W1B210,W1B220;
wire W1B001,W1B011,W1B021,W1B101,W1B111,W1B121,W1B201,W1B211,W1B221;
wire W1B002,W1B012,W1B022,W1B102,W1B112,W1B122,W1B202,W1B212,W1B222;
wire W1B003,W1B013,W1B023,W1B103,W1B113,W1B123,W1B203,W1B213,W1B223;
wire W1B004,W1B014,W1B024,W1B104,W1B114,W1B124,W1B204,W1B214,W1B224;
wire W1B005,W1B015,W1B025,W1B105,W1B115,W1B125,W1B205,W1B215,W1B225;
wire W1B006,W1B016,W1B026,W1B106,W1B116,W1B126,W1B206,W1B216,W1B226;
wire W1B007,W1B017,W1B027,W1B107,W1B117,W1B127,W1B207,W1B217,W1B227;
wire W1B008,W1B018,W1B028,W1B108,W1B118,W1B128,W1B208,W1B218,W1B228;
wire W1B009,W1B019,W1B029,W1B109,W1B119,W1B129,W1B209,W1B219,W1B229;
wire W1B00A,W1B01A,W1B02A,W1B10A,W1B11A,W1B12A,W1B20A,W1B21A,W1B22A;
wire W1B00B,W1B01B,W1B02B,W1B10B,W1B11B,W1B12B,W1B20B,W1B21B,W1B22B;
wire W1B00C,W1B01C,W1B02C,W1B10C,W1B11C,W1B12C,W1B20C,W1B21C,W1B22C;
wire W1B00D,W1B01D,W1B02D,W1B10D,W1B11D,W1B12D,W1B20D,W1B21D,W1B22D;
wire W1B00E,W1B01E,W1B02E,W1B10E,W1B11E,W1B12E,W1B20E,W1B21E,W1B22E;
wire W1B00F,W1B01F,W1B02F,W1B10F,W1B11F,W1B12F,W1B20F,W1B21F,W1B22F;
wire W1C000,W1C010,W1C020,W1C100,W1C110,W1C120,W1C200,W1C210,W1C220;
wire W1C001,W1C011,W1C021,W1C101,W1C111,W1C121,W1C201,W1C211,W1C221;
wire W1C002,W1C012,W1C022,W1C102,W1C112,W1C122,W1C202,W1C212,W1C222;
wire W1C003,W1C013,W1C023,W1C103,W1C113,W1C123,W1C203,W1C213,W1C223;
wire W1C004,W1C014,W1C024,W1C104,W1C114,W1C124,W1C204,W1C214,W1C224;
wire W1C005,W1C015,W1C025,W1C105,W1C115,W1C125,W1C205,W1C215,W1C225;
wire W1C006,W1C016,W1C026,W1C106,W1C116,W1C126,W1C206,W1C216,W1C226;
wire W1C007,W1C017,W1C027,W1C107,W1C117,W1C127,W1C207,W1C217,W1C227;
wire W1C008,W1C018,W1C028,W1C108,W1C118,W1C128,W1C208,W1C218,W1C228;
wire W1C009,W1C019,W1C029,W1C109,W1C119,W1C129,W1C209,W1C219,W1C229;
wire W1C00A,W1C01A,W1C02A,W1C10A,W1C11A,W1C12A,W1C20A,W1C21A,W1C22A;
wire W1C00B,W1C01B,W1C02B,W1C10B,W1C11B,W1C12B,W1C20B,W1C21B,W1C22B;
wire W1C00C,W1C01C,W1C02C,W1C10C,W1C11C,W1C12C,W1C20C,W1C21C,W1C22C;
wire W1C00D,W1C01D,W1C02D,W1C10D,W1C11D,W1C12D,W1C20D,W1C21D,W1C22D;
wire W1C00E,W1C01E,W1C02E,W1C10E,W1C11E,W1C12E,W1C20E,W1C21E,W1C22E;
wire W1C00F,W1C01F,W1C02F,W1C10F,W1C11F,W1C12F,W1C20F,W1C21F,W1C22F;
wire W1D000,W1D010,W1D020,W1D100,W1D110,W1D120,W1D200,W1D210,W1D220;
wire W1D001,W1D011,W1D021,W1D101,W1D111,W1D121,W1D201,W1D211,W1D221;
wire W1D002,W1D012,W1D022,W1D102,W1D112,W1D122,W1D202,W1D212,W1D222;
wire W1D003,W1D013,W1D023,W1D103,W1D113,W1D123,W1D203,W1D213,W1D223;
wire W1D004,W1D014,W1D024,W1D104,W1D114,W1D124,W1D204,W1D214,W1D224;
wire W1D005,W1D015,W1D025,W1D105,W1D115,W1D125,W1D205,W1D215,W1D225;
wire W1D006,W1D016,W1D026,W1D106,W1D116,W1D126,W1D206,W1D216,W1D226;
wire W1D007,W1D017,W1D027,W1D107,W1D117,W1D127,W1D207,W1D217,W1D227;
wire W1D008,W1D018,W1D028,W1D108,W1D118,W1D128,W1D208,W1D218,W1D228;
wire W1D009,W1D019,W1D029,W1D109,W1D119,W1D129,W1D209,W1D219,W1D229;
wire W1D00A,W1D01A,W1D02A,W1D10A,W1D11A,W1D12A,W1D20A,W1D21A,W1D22A;
wire W1D00B,W1D01B,W1D02B,W1D10B,W1D11B,W1D12B,W1D20B,W1D21B,W1D22B;
wire W1D00C,W1D01C,W1D02C,W1D10C,W1D11C,W1D12C,W1D20C,W1D21C,W1D22C;
wire W1D00D,W1D01D,W1D02D,W1D10D,W1D11D,W1D12D,W1D20D,W1D21D,W1D22D;
wire W1D00E,W1D01E,W1D02E,W1D10E,W1D11E,W1D12E,W1D20E,W1D21E,W1D22E;
wire W1D00F,W1D01F,W1D02F,W1D10F,W1D11F,W1D12F,W1D20F,W1D21F,W1D22F;
wire W1E000,W1E010,W1E020,W1E100,W1E110,W1E120,W1E200,W1E210,W1E220;
wire W1E001,W1E011,W1E021,W1E101,W1E111,W1E121,W1E201,W1E211,W1E221;
wire W1E002,W1E012,W1E022,W1E102,W1E112,W1E122,W1E202,W1E212,W1E222;
wire W1E003,W1E013,W1E023,W1E103,W1E113,W1E123,W1E203,W1E213,W1E223;
wire W1E004,W1E014,W1E024,W1E104,W1E114,W1E124,W1E204,W1E214,W1E224;
wire W1E005,W1E015,W1E025,W1E105,W1E115,W1E125,W1E205,W1E215,W1E225;
wire W1E006,W1E016,W1E026,W1E106,W1E116,W1E126,W1E206,W1E216,W1E226;
wire W1E007,W1E017,W1E027,W1E107,W1E117,W1E127,W1E207,W1E217,W1E227;
wire W1E008,W1E018,W1E028,W1E108,W1E118,W1E128,W1E208,W1E218,W1E228;
wire W1E009,W1E019,W1E029,W1E109,W1E119,W1E129,W1E209,W1E219,W1E229;
wire W1E00A,W1E01A,W1E02A,W1E10A,W1E11A,W1E12A,W1E20A,W1E21A,W1E22A;
wire W1E00B,W1E01B,W1E02B,W1E10B,W1E11B,W1E12B,W1E20B,W1E21B,W1E22B;
wire W1E00C,W1E01C,W1E02C,W1E10C,W1E11C,W1E12C,W1E20C,W1E21C,W1E22C;
wire W1E00D,W1E01D,W1E02D,W1E10D,W1E11D,W1E12D,W1E20D,W1E21D,W1E22D;
wire W1E00E,W1E01E,W1E02E,W1E10E,W1E11E,W1E12E,W1E20E,W1E21E,W1E22E;
wire W1E00F,W1E01F,W1E02F,W1E10F,W1E11F,W1E12F,W1E20F,W1E21F,W1E22F;
wire W1F000,W1F010,W1F020,W1F100,W1F110,W1F120,W1F200,W1F210,W1F220;
wire W1F001,W1F011,W1F021,W1F101,W1F111,W1F121,W1F201,W1F211,W1F221;
wire W1F002,W1F012,W1F022,W1F102,W1F112,W1F122,W1F202,W1F212,W1F222;
wire W1F003,W1F013,W1F023,W1F103,W1F113,W1F123,W1F203,W1F213,W1F223;
wire W1F004,W1F014,W1F024,W1F104,W1F114,W1F124,W1F204,W1F214,W1F224;
wire W1F005,W1F015,W1F025,W1F105,W1F115,W1F125,W1F205,W1F215,W1F225;
wire W1F006,W1F016,W1F026,W1F106,W1F116,W1F126,W1F206,W1F216,W1F226;
wire W1F007,W1F017,W1F027,W1F107,W1F117,W1F127,W1F207,W1F217,W1F227;
wire W1F008,W1F018,W1F028,W1F108,W1F118,W1F128,W1F208,W1F218,W1F228;
wire W1F009,W1F019,W1F029,W1F109,W1F119,W1F129,W1F209,W1F219,W1F229;
wire W1F00A,W1F01A,W1F02A,W1F10A,W1F11A,W1F12A,W1F20A,W1F21A,W1F22A;
wire W1F00B,W1F01B,W1F02B,W1F10B,W1F11B,W1F12B,W1F20B,W1F21B,W1F22B;
wire W1F00C,W1F01C,W1F02C,W1F10C,W1F11C,W1F12C,W1F20C,W1F21C,W1F22C;
wire W1F00D,W1F01D,W1F02D,W1F10D,W1F11D,W1F12D,W1F20D,W1F21D,W1F22D;
wire W1F00E,W1F01E,W1F02E,W1F10E,W1F11E,W1F12E,W1F20E,W1F21E,W1F22E;
wire W1F00F,W1F01F,W1F02F,W1F10F,W1F11F,W1F12F,W1F20F,W1F21F,W1F22F;
wire W1G000,W1G010,W1G020,W1G100,W1G110,W1G120,W1G200,W1G210,W1G220;
wire W1G001,W1G011,W1G021,W1G101,W1G111,W1G121,W1G201,W1G211,W1G221;
wire W1G002,W1G012,W1G022,W1G102,W1G112,W1G122,W1G202,W1G212,W1G222;
wire W1G003,W1G013,W1G023,W1G103,W1G113,W1G123,W1G203,W1G213,W1G223;
wire W1G004,W1G014,W1G024,W1G104,W1G114,W1G124,W1G204,W1G214,W1G224;
wire W1G005,W1G015,W1G025,W1G105,W1G115,W1G125,W1G205,W1G215,W1G225;
wire W1G006,W1G016,W1G026,W1G106,W1G116,W1G126,W1G206,W1G216,W1G226;
wire W1G007,W1G017,W1G027,W1G107,W1G117,W1G127,W1G207,W1G217,W1G227;
wire W1G008,W1G018,W1G028,W1G108,W1G118,W1G128,W1G208,W1G218,W1G228;
wire W1G009,W1G019,W1G029,W1G109,W1G119,W1G129,W1G209,W1G219,W1G229;
wire W1G00A,W1G01A,W1G02A,W1G10A,W1G11A,W1G12A,W1G20A,W1G21A,W1G22A;
wire W1G00B,W1G01B,W1G02B,W1G10B,W1G11B,W1G12B,W1G20B,W1G21B,W1G22B;
wire W1G00C,W1G01C,W1G02C,W1G10C,W1G11C,W1G12C,W1G20C,W1G21C,W1G22C;
wire W1G00D,W1G01D,W1G02D,W1G10D,W1G11D,W1G12D,W1G20D,W1G21D,W1G22D;
wire W1G00E,W1G01E,W1G02E,W1G10E,W1G11E,W1G12E,W1G20E,W1G21E,W1G22E;
wire W1G00F,W1G01F,W1G02F,W1G10F,W1G11F,W1G12F,W1G20F,W1G21F,W1G22F;
wire W1H000,W1H010,W1H020,W1H100,W1H110,W1H120,W1H200,W1H210,W1H220;
wire W1H001,W1H011,W1H021,W1H101,W1H111,W1H121,W1H201,W1H211,W1H221;
wire W1H002,W1H012,W1H022,W1H102,W1H112,W1H122,W1H202,W1H212,W1H222;
wire W1H003,W1H013,W1H023,W1H103,W1H113,W1H123,W1H203,W1H213,W1H223;
wire W1H004,W1H014,W1H024,W1H104,W1H114,W1H124,W1H204,W1H214,W1H224;
wire W1H005,W1H015,W1H025,W1H105,W1H115,W1H125,W1H205,W1H215,W1H225;
wire W1H006,W1H016,W1H026,W1H106,W1H116,W1H126,W1H206,W1H216,W1H226;
wire W1H007,W1H017,W1H027,W1H107,W1H117,W1H127,W1H207,W1H217,W1H227;
wire W1H008,W1H018,W1H028,W1H108,W1H118,W1H128,W1H208,W1H218,W1H228;
wire W1H009,W1H019,W1H029,W1H109,W1H119,W1H129,W1H209,W1H219,W1H229;
wire W1H00A,W1H01A,W1H02A,W1H10A,W1H11A,W1H12A,W1H20A,W1H21A,W1H22A;
wire W1H00B,W1H01B,W1H02B,W1H10B,W1H11B,W1H12B,W1H20B,W1H21B,W1H22B;
wire W1H00C,W1H01C,W1H02C,W1H10C,W1H11C,W1H12C,W1H20C,W1H21C,W1H22C;
wire W1H00D,W1H01D,W1H02D,W1H10D,W1H11D,W1H12D,W1H20D,W1H21D,W1H22D;
wire W1H00E,W1H01E,W1H02E,W1H10E,W1H11E,W1H12E,W1H20E,W1H21E,W1H22E;
wire W1H00F,W1H01F,W1H02F,W1H10F,W1H11F,W1H12F,W1H20F,W1H21F,W1H22F;
wire W1I000,W1I010,W1I020,W1I100,W1I110,W1I120,W1I200,W1I210,W1I220;
wire W1I001,W1I011,W1I021,W1I101,W1I111,W1I121,W1I201,W1I211,W1I221;
wire W1I002,W1I012,W1I022,W1I102,W1I112,W1I122,W1I202,W1I212,W1I222;
wire W1I003,W1I013,W1I023,W1I103,W1I113,W1I123,W1I203,W1I213,W1I223;
wire W1I004,W1I014,W1I024,W1I104,W1I114,W1I124,W1I204,W1I214,W1I224;
wire W1I005,W1I015,W1I025,W1I105,W1I115,W1I125,W1I205,W1I215,W1I225;
wire W1I006,W1I016,W1I026,W1I106,W1I116,W1I126,W1I206,W1I216,W1I226;
wire W1I007,W1I017,W1I027,W1I107,W1I117,W1I127,W1I207,W1I217,W1I227;
wire W1I008,W1I018,W1I028,W1I108,W1I118,W1I128,W1I208,W1I218,W1I228;
wire W1I009,W1I019,W1I029,W1I109,W1I119,W1I129,W1I209,W1I219,W1I229;
wire W1I00A,W1I01A,W1I02A,W1I10A,W1I11A,W1I12A,W1I20A,W1I21A,W1I22A;
wire W1I00B,W1I01B,W1I02B,W1I10B,W1I11B,W1I12B,W1I20B,W1I21B,W1I22B;
wire W1I00C,W1I01C,W1I02C,W1I10C,W1I11C,W1I12C,W1I20C,W1I21C,W1I22C;
wire W1I00D,W1I01D,W1I02D,W1I10D,W1I11D,W1I12D,W1I20D,W1I21D,W1I22D;
wire W1I00E,W1I01E,W1I02E,W1I10E,W1I11E,W1I12E,W1I20E,W1I21E,W1I22E;
wire W1I00F,W1I01F,W1I02F,W1I10F,W1I11F,W1I12F,W1I20F,W1I21F,W1I22F;
wire W1J000,W1J010,W1J020,W1J100,W1J110,W1J120,W1J200,W1J210,W1J220;
wire W1J001,W1J011,W1J021,W1J101,W1J111,W1J121,W1J201,W1J211,W1J221;
wire W1J002,W1J012,W1J022,W1J102,W1J112,W1J122,W1J202,W1J212,W1J222;
wire W1J003,W1J013,W1J023,W1J103,W1J113,W1J123,W1J203,W1J213,W1J223;
wire W1J004,W1J014,W1J024,W1J104,W1J114,W1J124,W1J204,W1J214,W1J224;
wire W1J005,W1J015,W1J025,W1J105,W1J115,W1J125,W1J205,W1J215,W1J225;
wire W1J006,W1J016,W1J026,W1J106,W1J116,W1J126,W1J206,W1J216,W1J226;
wire W1J007,W1J017,W1J027,W1J107,W1J117,W1J127,W1J207,W1J217,W1J227;
wire W1J008,W1J018,W1J028,W1J108,W1J118,W1J128,W1J208,W1J218,W1J228;
wire W1J009,W1J019,W1J029,W1J109,W1J119,W1J129,W1J209,W1J219,W1J229;
wire W1J00A,W1J01A,W1J02A,W1J10A,W1J11A,W1J12A,W1J20A,W1J21A,W1J22A;
wire W1J00B,W1J01B,W1J02B,W1J10B,W1J11B,W1J12B,W1J20B,W1J21B,W1J22B;
wire W1J00C,W1J01C,W1J02C,W1J10C,W1J11C,W1J12C,W1J20C,W1J21C,W1J22C;
wire W1J00D,W1J01D,W1J02D,W1J10D,W1J11D,W1J12D,W1J20D,W1J21D,W1J22D;
wire W1J00E,W1J01E,W1J02E,W1J10E,W1J11E,W1J12E,W1J20E,W1J21E,W1J22E;
wire W1J00F,W1J01F,W1J02F,W1J10F,W1J11F,W1J12F,W1J20F,W1J21F,W1J22F;
wire W1K000,W1K010,W1K020,W1K100,W1K110,W1K120,W1K200,W1K210,W1K220;
wire W1K001,W1K011,W1K021,W1K101,W1K111,W1K121,W1K201,W1K211,W1K221;
wire W1K002,W1K012,W1K022,W1K102,W1K112,W1K122,W1K202,W1K212,W1K222;
wire W1K003,W1K013,W1K023,W1K103,W1K113,W1K123,W1K203,W1K213,W1K223;
wire W1K004,W1K014,W1K024,W1K104,W1K114,W1K124,W1K204,W1K214,W1K224;
wire W1K005,W1K015,W1K025,W1K105,W1K115,W1K125,W1K205,W1K215,W1K225;
wire W1K006,W1K016,W1K026,W1K106,W1K116,W1K126,W1K206,W1K216,W1K226;
wire W1K007,W1K017,W1K027,W1K107,W1K117,W1K127,W1K207,W1K217,W1K227;
wire W1K008,W1K018,W1K028,W1K108,W1K118,W1K128,W1K208,W1K218,W1K228;
wire W1K009,W1K019,W1K029,W1K109,W1K119,W1K129,W1K209,W1K219,W1K229;
wire W1K00A,W1K01A,W1K02A,W1K10A,W1K11A,W1K12A,W1K20A,W1K21A,W1K22A;
wire W1K00B,W1K01B,W1K02B,W1K10B,W1K11B,W1K12B,W1K20B,W1K21B,W1K22B;
wire W1K00C,W1K01C,W1K02C,W1K10C,W1K11C,W1K12C,W1K20C,W1K21C,W1K22C;
wire W1K00D,W1K01D,W1K02D,W1K10D,W1K11D,W1K12D,W1K20D,W1K21D,W1K22D;
wire W1K00E,W1K01E,W1K02E,W1K10E,W1K11E,W1K12E,W1K20E,W1K21E,W1K22E;
wire W1K00F,W1K01F,W1K02F,W1K10F,W1K11F,W1K12F,W1K20F,W1K21F,W1K22F;
wire W1L000,W1L010,W1L020,W1L100,W1L110,W1L120,W1L200,W1L210,W1L220;
wire W1L001,W1L011,W1L021,W1L101,W1L111,W1L121,W1L201,W1L211,W1L221;
wire W1L002,W1L012,W1L022,W1L102,W1L112,W1L122,W1L202,W1L212,W1L222;
wire W1L003,W1L013,W1L023,W1L103,W1L113,W1L123,W1L203,W1L213,W1L223;
wire W1L004,W1L014,W1L024,W1L104,W1L114,W1L124,W1L204,W1L214,W1L224;
wire W1L005,W1L015,W1L025,W1L105,W1L115,W1L125,W1L205,W1L215,W1L225;
wire W1L006,W1L016,W1L026,W1L106,W1L116,W1L126,W1L206,W1L216,W1L226;
wire W1L007,W1L017,W1L027,W1L107,W1L117,W1L127,W1L207,W1L217,W1L227;
wire W1L008,W1L018,W1L028,W1L108,W1L118,W1L128,W1L208,W1L218,W1L228;
wire W1L009,W1L019,W1L029,W1L109,W1L119,W1L129,W1L209,W1L219,W1L229;
wire W1L00A,W1L01A,W1L02A,W1L10A,W1L11A,W1L12A,W1L20A,W1L21A,W1L22A;
wire W1L00B,W1L01B,W1L02B,W1L10B,W1L11B,W1L12B,W1L20B,W1L21B,W1L22B;
wire W1L00C,W1L01C,W1L02C,W1L10C,W1L11C,W1L12C,W1L20C,W1L21C,W1L22C;
wire W1L00D,W1L01D,W1L02D,W1L10D,W1L11D,W1L12D,W1L20D,W1L21D,W1L22D;
wire W1L00E,W1L01E,W1L02E,W1L10E,W1L11E,W1L12E,W1L20E,W1L21E,W1L22E;
wire W1L00F,W1L01F,W1L02F,W1L10F,W1L11F,W1L12F,W1L20F,W1L21F,W1L22F;
wire W1M000,W1M010,W1M020,W1M100,W1M110,W1M120,W1M200,W1M210,W1M220;
wire W1M001,W1M011,W1M021,W1M101,W1M111,W1M121,W1M201,W1M211,W1M221;
wire W1M002,W1M012,W1M022,W1M102,W1M112,W1M122,W1M202,W1M212,W1M222;
wire W1M003,W1M013,W1M023,W1M103,W1M113,W1M123,W1M203,W1M213,W1M223;
wire W1M004,W1M014,W1M024,W1M104,W1M114,W1M124,W1M204,W1M214,W1M224;
wire W1M005,W1M015,W1M025,W1M105,W1M115,W1M125,W1M205,W1M215,W1M225;
wire W1M006,W1M016,W1M026,W1M106,W1M116,W1M126,W1M206,W1M216,W1M226;
wire W1M007,W1M017,W1M027,W1M107,W1M117,W1M127,W1M207,W1M217,W1M227;
wire W1M008,W1M018,W1M028,W1M108,W1M118,W1M128,W1M208,W1M218,W1M228;
wire W1M009,W1M019,W1M029,W1M109,W1M119,W1M129,W1M209,W1M219,W1M229;
wire W1M00A,W1M01A,W1M02A,W1M10A,W1M11A,W1M12A,W1M20A,W1M21A,W1M22A;
wire W1M00B,W1M01B,W1M02B,W1M10B,W1M11B,W1M12B,W1M20B,W1M21B,W1M22B;
wire W1M00C,W1M01C,W1M02C,W1M10C,W1M11C,W1M12C,W1M20C,W1M21C,W1M22C;
wire W1M00D,W1M01D,W1M02D,W1M10D,W1M11D,W1M12D,W1M20D,W1M21D,W1M22D;
wire W1M00E,W1M01E,W1M02E,W1M10E,W1M11E,W1M12E,W1M20E,W1M21E,W1M22E;
wire W1M00F,W1M01F,W1M02F,W1M10F,W1M11F,W1M12F,W1M20F,W1M21F,W1M22F;
wire signed [4:0] c10000,c11000,c12000,c13000,c14000,c15000,c16000,c17000,c18000,c19000,c1A000,c1B000,c1C000,c1D000,c1E000,c1F000;
wire signed [4:0] c10010,c11010,c12010,c13010,c14010,c15010,c16010,c17010,c18010,c19010,c1A010,c1B010,c1C010,c1D010,c1E010,c1F010;
wire signed [4:0] c10020,c11020,c12020,c13020,c14020,c15020,c16020,c17020,c18020,c19020,c1A020,c1B020,c1C020,c1D020,c1E020,c1F020;
wire signed [4:0] c10100,c11100,c12100,c13100,c14100,c15100,c16100,c17100,c18100,c19100,c1A100,c1B100,c1C100,c1D100,c1E100,c1F100;
wire signed [4:0] c10110,c11110,c12110,c13110,c14110,c15110,c16110,c17110,c18110,c19110,c1A110,c1B110,c1C110,c1D110,c1E110,c1F110;
wire signed [4:0] c10120,c11120,c12120,c13120,c14120,c15120,c16120,c17120,c18120,c19120,c1A120,c1B120,c1C120,c1D120,c1E120,c1F120;
wire signed [4:0] c10200,c11200,c12200,c13200,c14200,c15200,c16200,c17200,c18200,c19200,c1A200,c1B200,c1C200,c1D200,c1E200,c1F200;
wire signed [4:0] c10210,c11210,c12210,c13210,c14210,c15210,c16210,c17210,c18210,c19210,c1A210,c1B210,c1C210,c1D210,c1E210,c1F210;
wire signed [4:0] c10220,c11220,c12220,c13220,c14220,c15220,c16220,c17220,c18220,c19220,c1A220,c1B220,c1C220,c1D220,c1E220,c1F220;
wire signed [4:0] c10001,c11001,c12001,c13001,c14001,c15001,c16001,c17001,c18001,c19001,c1A001,c1B001,c1C001,c1D001,c1E001,c1F001;
wire signed [4:0] c10011,c11011,c12011,c13011,c14011,c15011,c16011,c17011,c18011,c19011,c1A011,c1B011,c1C011,c1D011,c1E011,c1F011;
wire signed [4:0] c10021,c11021,c12021,c13021,c14021,c15021,c16021,c17021,c18021,c19021,c1A021,c1B021,c1C021,c1D021,c1E021,c1F021;
wire signed [4:0] c10101,c11101,c12101,c13101,c14101,c15101,c16101,c17101,c18101,c19101,c1A101,c1B101,c1C101,c1D101,c1E101,c1F101;
wire signed [4:0] c10111,c11111,c12111,c13111,c14111,c15111,c16111,c17111,c18111,c19111,c1A111,c1B111,c1C111,c1D111,c1E111,c1F111;
wire signed [4:0] c10121,c11121,c12121,c13121,c14121,c15121,c16121,c17121,c18121,c19121,c1A121,c1B121,c1C121,c1D121,c1E121,c1F121;
wire signed [4:0] c10201,c11201,c12201,c13201,c14201,c15201,c16201,c17201,c18201,c19201,c1A201,c1B201,c1C201,c1D201,c1E201,c1F201;
wire signed [4:0] c10211,c11211,c12211,c13211,c14211,c15211,c16211,c17211,c18211,c19211,c1A211,c1B211,c1C211,c1D211,c1E211,c1F211;
wire signed [4:0] c10221,c11221,c12221,c13221,c14221,c15221,c16221,c17221,c18221,c19221,c1A221,c1B221,c1C221,c1D221,c1E221,c1F221;
wire signed [4:0] c10002,c11002,c12002,c13002,c14002,c15002,c16002,c17002,c18002,c19002,c1A002,c1B002,c1C002,c1D002,c1E002,c1F002;
wire signed [4:0] c10012,c11012,c12012,c13012,c14012,c15012,c16012,c17012,c18012,c19012,c1A012,c1B012,c1C012,c1D012,c1E012,c1F012;
wire signed [4:0] c10022,c11022,c12022,c13022,c14022,c15022,c16022,c17022,c18022,c19022,c1A022,c1B022,c1C022,c1D022,c1E022,c1F022;
wire signed [4:0] c10102,c11102,c12102,c13102,c14102,c15102,c16102,c17102,c18102,c19102,c1A102,c1B102,c1C102,c1D102,c1E102,c1F102;
wire signed [4:0] c10112,c11112,c12112,c13112,c14112,c15112,c16112,c17112,c18112,c19112,c1A112,c1B112,c1C112,c1D112,c1E112,c1F112;
wire signed [4:0] c10122,c11122,c12122,c13122,c14122,c15122,c16122,c17122,c18122,c19122,c1A122,c1B122,c1C122,c1D122,c1E122,c1F122;
wire signed [4:0] c10202,c11202,c12202,c13202,c14202,c15202,c16202,c17202,c18202,c19202,c1A202,c1B202,c1C202,c1D202,c1E202,c1F202;
wire signed [4:0] c10212,c11212,c12212,c13212,c14212,c15212,c16212,c17212,c18212,c19212,c1A212,c1B212,c1C212,c1D212,c1E212,c1F212;
wire signed [4:0] c10222,c11222,c12222,c13222,c14222,c15222,c16222,c17222,c18222,c19222,c1A222,c1B222,c1C222,c1D222,c1E222,c1F222;
wire signed [4:0] c10003,c11003,c12003,c13003,c14003,c15003,c16003,c17003,c18003,c19003,c1A003,c1B003,c1C003,c1D003,c1E003,c1F003;
wire signed [4:0] c10013,c11013,c12013,c13013,c14013,c15013,c16013,c17013,c18013,c19013,c1A013,c1B013,c1C013,c1D013,c1E013,c1F013;
wire signed [4:0] c10023,c11023,c12023,c13023,c14023,c15023,c16023,c17023,c18023,c19023,c1A023,c1B023,c1C023,c1D023,c1E023,c1F023;
wire signed [4:0] c10103,c11103,c12103,c13103,c14103,c15103,c16103,c17103,c18103,c19103,c1A103,c1B103,c1C103,c1D103,c1E103,c1F103;
wire signed [4:0] c10113,c11113,c12113,c13113,c14113,c15113,c16113,c17113,c18113,c19113,c1A113,c1B113,c1C113,c1D113,c1E113,c1F113;
wire signed [4:0] c10123,c11123,c12123,c13123,c14123,c15123,c16123,c17123,c18123,c19123,c1A123,c1B123,c1C123,c1D123,c1E123,c1F123;
wire signed [4:0] c10203,c11203,c12203,c13203,c14203,c15203,c16203,c17203,c18203,c19203,c1A203,c1B203,c1C203,c1D203,c1E203,c1F203;
wire signed [4:0] c10213,c11213,c12213,c13213,c14213,c15213,c16213,c17213,c18213,c19213,c1A213,c1B213,c1C213,c1D213,c1E213,c1F213;
wire signed [4:0] c10223,c11223,c12223,c13223,c14223,c15223,c16223,c17223,c18223,c19223,c1A223,c1B223,c1C223,c1D223,c1E223,c1F223;
wire signed [4:0] c10004,c11004,c12004,c13004,c14004,c15004,c16004,c17004,c18004,c19004,c1A004,c1B004,c1C004,c1D004,c1E004,c1F004;
wire signed [4:0] c10014,c11014,c12014,c13014,c14014,c15014,c16014,c17014,c18014,c19014,c1A014,c1B014,c1C014,c1D014,c1E014,c1F014;
wire signed [4:0] c10024,c11024,c12024,c13024,c14024,c15024,c16024,c17024,c18024,c19024,c1A024,c1B024,c1C024,c1D024,c1E024,c1F024;
wire signed [4:0] c10104,c11104,c12104,c13104,c14104,c15104,c16104,c17104,c18104,c19104,c1A104,c1B104,c1C104,c1D104,c1E104,c1F104;
wire signed [4:0] c10114,c11114,c12114,c13114,c14114,c15114,c16114,c17114,c18114,c19114,c1A114,c1B114,c1C114,c1D114,c1E114,c1F114;
wire signed [4:0] c10124,c11124,c12124,c13124,c14124,c15124,c16124,c17124,c18124,c19124,c1A124,c1B124,c1C124,c1D124,c1E124,c1F124;
wire signed [4:0] c10204,c11204,c12204,c13204,c14204,c15204,c16204,c17204,c18204,c19204,c1A204,c1B204,c1C204,c1D204,c1E204,c1F204;
wire signed [4:0] c10214,c11214,c12214,c13214,c14214,c15214,c16214,c17214,c18214,c19214,c1A214,c1B214,c1C214,c1D214,c1E214,c1F214;
wire signed [4:0] c10224,c11224,c12224,c13224,c14224,c15224,c16224,c17224,c18224,c19224,c1A224,c1B224,c1C224,c1D224,c1E224,c1F224;
wire signed [4:0] c10005,c11005,c12005,c13005,c14005,c15005,c16005,c17005,c18005,c19005,c1A005,c1B005,c1C005,c1D005,c1E005,c1F005;
wire signed [4:0] c10015,c11015,c12015,c13015,c14015,c15015,c16015,c17015,c18015,c19015,c1A015,c1B015,c1C015,c1D015,c1E015,c1F015;
wire signed [4:0] c10025,c11025,c12025,c13025,c14025,c15025,c16025,c17025,c18025,c19025,c1A025,c1B025,c1C025,c1D025,c1E025,c1F025;
wire signed [4:0] c10105,c11105,c12105,c13105,c14105,c15105,c16105,c17105,c18105,c19105,c1A105,c1B105,c1C105,c1D105,c1E105,c1F105;
wire signed [4:0] c10115,c11115,c12115,c13115,c14115,c15115,c16115,c17115,c18115,c19115,c1A115,c1B115,c1C115,c1D115,c1E115,c1F115;
wire signed [4:0] c10125,c11125,c12125,c13125,c14125,c15125,c16125,c17125,c18125,c19125,c1A125,c1B125,c1C125,c1D125,c1E125,c1F125;
wire signed [4:0] c10205,c11205,c12205,c13205,c14205,c15205,c16205,c17205,c18205,c19205,c1A205,c1B205,c1C205,c1D205,c1E205,c1F205;
wire signed [4:0] c10215,c11215,c12215,c13215,c14215,c15215,c16215,c17215,c18215,c19215,c1A215,c1B215,c1C215,c1D215,c1E215,c1F215;
wire signed [4:0] c10225,c11225,c12225,c13225,c14225,c15225,c16225,c17225,c18225,c19225,c1A225,c1B225,c1C225,c1D225,c1E225,c1F225;
wire signed [4:0] c10006,c11006,c12006,c13006,c14006,c15006,c16006,c17006,c18006,c19006,c1A006,c1B006,c1C006,c1D006,c1E006,c1F006;
wire signed [4:0] c10016,c11016,c12016,c13016,c14016,c15016,c16016,c17016,c18016,c19016,c1A016,c1B016,c1C016,c1D016,c1E016,c1F016;
wire signed [4:0] c10026,c11026,c12026,c13026,c14026,c15026,c16026,c17026,c18026,c19026,c1A026,c1B026,c1C026,c1D026,c1E026,c1F026;
wire signed [4:0] c10106,c11106,c12106,c13106,c14106,c15106,c16106,c17106,c18106,c19106,c1A106,c1B106,c1C106,c1D106,c1E106,c1F106;
wire signed [4:0] c10116,c11116,c12116,c13116,c14116,c15116,c16116,c17116,c18116,c19116,c1A116,c1B116,c1C116,c1D116,c1E116,c1F116;
wire signed [4:0] c10126,c11126,c12126,c13126,c14126,c15126,c16126,c17126,c18126,c19126,c1A126,c1B126,c1C126,c1D126,c1E126,c1F126;
wire signed [4:0] c10206,c11206,c12206,c13206,c14206,c15206,c16206,c17206,c18206,c19206,c1A206,c1B206,c1C206,c1D206,c1E206,c1F206;
wire signed [4:0] c10216,c11216,c12216,c13216,c14216,c15216,c16216,c17216,c18216,c19216,c1A216,c1B216,c1C216,c1D216,c1E216,c1F216;
wire signed [4:0] c10226,c11226,c12226,c13226,c14226,c15226,c16226,c17226,c18226,c19226,c1A226,c1B226,c1C226,c1D226,c1E226,c1F226;
wire signed [4:0] c10007,c11007,c12007,c13007,c14007,c15007,c16007,c17007,c18007,c19007,c1A007,c1B007,c1C007,c1D007,c1E007,c1F007;
wire signed [4:0] c10017,c11017,c12017,c13017,c14017,c15017,c16017,c17017,c18017,c19017,c1A017,c1B017,c1C017,c1D017,c1E017,c1F017;
wire signed [4:0] c10027,c11027,c12027,c13027,c14027,c15027,c16027,c17027,c18027,c19027,c1A027,c1B027,c1C027,c1D027,c1E027,c1F027;
wire signed [4:0] c10107,c11107,c12107,c13107,c14107,c15107,c16107,c17107,c18107,c19107,c1A107,c1B107,c1C107,c1D107,c1E107,c1F107;
wire signed [4:0] c10117,c11117,c12117,c13117,c14117,c15117,c16117,c17117,c18117,c19117,c1A117,c1B117,c1C117,c1D117,c1E117,c1F117;
wire signed [4:0] c10127,c11127,c12127,c13127,c14127,c15127,c16127,c17127,c18127,c19127,c1A127,c1B127,c1C127,c1D127,c1E127,c1F127;
wire signed [4:0] c10207,c11207,c12207,c13207,c14207,c15207,c16207,c17207,c18207,c19207,c1A207,c1B207,c1C207,c1D207,c1E207,c1F207;
wire signed [4:0] c10217,c11217,c12217,c13217,c14217,c15217,c16217,c17217,c18217,c19217,c1A217,c1B217,c1C217,c1D217,c1E217,c1F217;
wire signed [4:0] c10227,c11227,c12227,c13227,c14227,c15227,c16227,c17227,c18227,c19227,c1A227,c1B227,c1C227,c1D227,c1E227,c1F227;
wire signed [4:0] c10008,c11008,c12008,c13008,c14008,c15008,c16008,c17008,c18008,c19008,c1A008,c1B008,c1C008,c1D008,c1E008,c1F008;
wire signed [4:0] c10018,c11018,c12018,c13018,c14018,c15018,c16018,c17018,c18018,c19018,c1A018,c1B018,c1C018,c1D018,c1E018,c1F018;
wire signed [4:0] c10028,c11028,c12028,c13028,c14028,c15028,c16028,c17028,c18028,c19028,c1A028,c1B028,c1C028,c1D028,c1E028,c1F028;
wire signed [4:0] c10108,c11108,c12108,c13108,c14108,c15108,c16108,c17108,c18108,c19108,c1A108,c1B108,c1C108,c1D108,c1E108,c1F108;
wire signed [4:0] c10118,c11118,c12118,c13118,c14118,c15118,c16118,c17118,c18118,c19118,c1A118,c1B118,c1C118,c1D118,c1E118,c1F118;
wire signed [4:0] c10128,c11128,c12128,c13128,c14128,c15128,c16128,c17128,c18128,c19128,c1A128,c1B128,c1C128,c1D128,c1E128,c1F128;
wire signed [4:0] c10208,c11208,c12208,c13208,c14208,c15208,c16208,c17208,c18208,c19208,c1A208,c1B208,c1C208,c1D208,c1E208,c1F208;
wire signed [4:0] c10218,c11218,c12218,c13218,c14218,c15218,c16218,c17218,c18218,c19218,c1A218,c1B218,c1C218,c1D218,c1E218,c1F218;
wire signed [4:0] c10228,c11228,c12228,c13228,c14228,c15228,c16228,c17228,c18228,c19228,c1A228,c1B228,c1C228,c1D228,c1E228,c1F228;
wire signed [4:0] c10009,c11009,c12009,c13009,c14009,c15009,c16009,c17009,c18009,c19009,c1A009,c1B009,c1C009,c1D009,c1E009,c1F009;
wire signed [4:0] c10019,c11019,c12019,c13019,c14019,c15019,c16019,c17019,c18019,c19019,c1A019,c1B019,c1C019,c1D019,c1E019,c1F019;
wire signed [4:0] c10029,c11029,c12029,c13029,c14029,c15029,c16029,c17029,c18029,c19029,c1A029,c1B029,c1C029,c1D029,c1E029,c1F029;
wire signed [4:0] c10109,c11109,c12109,c13109,c14109,c15109,c16109,c17109,c18109,c19109,c1A109,c1B109,c1C109,c1D109,c1E109,c1F109;
wire signed [4:0] c10119,c11119,c12119,c13119,c14119,c15119,c16119,c17119,c18119,c19119,c1A119,c1B119,c1C119,c1D119,c1E119,c1F119;
wire signed [4:0] c10129,c11129,c12129,c13129,c14129,c15129,c16129,c17129,c18129,c19129,c1A129,c1B129,c1C129,c1D129,c1E129,c1F129;
wire signed [4:0] c10209,c11209,c12209,c13209,c14209,c15209,c16209,c17209,c18209,c19209,c1A209,c1B209,c1C209,c1D209,c1E209,c1F209;
wire signed [4:0] c10219,c11219,c12219,c13219,c14219,c15219,c16219,c17219,c18219,c19219,c1A219,c1B219,c1C219,c1D219,c1E219,c1F219;
wire signed [4:0] c10229,c11229,c12229,c13229,c14229,c15229,c16229,c17229,c18229,c19229,c1A229,c1B229,c1C229,c1D229,c1E229,c1F229;
wire signed [4:0] c1000A,c1100A,c1200A,c1300A,c1400A,c1500A,c1600A,c1700A,c1800A,c1900A,c1A00A,c1B00A,c1C00A,c1D00A,c1E00A,c1F00A;
wire signed [4:0] c1001A,c1101A,c1201A,c1301A,c1401A,c1501A,c1601A,c1701A,c1801A,c1901A,c1A01A,c1B01A,c1C01A,c1D01A,c1E01A,c1F01A;
wire signed [4:0] c1002A,c1102A,c1202A,c1302A,c1402A,c1502A,c1602A,c1702A,c1802A,c1902A,c1A02A,c1B02A,c1C02A,c1D02A,c1E02A,c1F02A;
wire signed [4:0] c1010A,c1110A,c1210A,c1310A,c1410A,c1510A,c1610A,c1710A,c1810A,c1910A,c1A10A,c1B10A,c1C10A,c1D10A,c1E10A,c1F10A;
wire signed [4:0] c1011A,c1111A,c1211A,c1311A,c1411A,c1511A,c1611A,c1711A,c1811A,c1911A,c1A11A,c1B11A,c1C11A,c1D11A,c1E11A,c1F11A;
wire signed [4:0] c1012A,c1112A,c1212A,c1312A,c1412A,c1512A,c1612A,c1712A,c1812A,c1912A,c1A12A,c1B12A,c1C12A,c1D12A,c1E12A,c1F12A;
wire signed [4:0] c1020A,c1120A,c1220A,c1320A,c1420A,c1520A,c1620A,c1720A,c1820A,c1920A,c1A20A,c1B20A,c1C20A,c1D20A,c1E20A,c1F20A;
wire signed [4:0] c1021A,c1121A,c1221A,c1321A,c1421A,c1521A,c1621A,c1721A,c1821A,c1921A,c1A21A,c1B21A,c1C21A,c1D21A,c1E21A,c1F21A;
wire signed [4:0] c1022A,c1122A,c1222A,c1322A,c1422A,c1522A,c1622A,c1722A,c1822A,c1922A,c1A22A,c1B22A,c1C22A,c1D22A,c1E22A,c1F22A;
wire signed [4:0] c1000B,c1100B,c1200B,c1300B,c1400B,c1500B,c1600B,c1700B,c1800B,c1900B,c1A00B,c1B00B,c1C00B,c1D00B,c1E00B,c1F00B;
wire signed [4:0] c1001B,c1101B,c1201B,c1301B,c1401B,c1501B,c1601B,c1701B,c1801B,c1901B,c1A01B,c1B01B,c1C01B,c1D01B,c1E01B,c1F01B;
wire signed [4:0] c1002B,c1102B,c1202B,c1302B,c1402B,c1502B,c1602B,c1702B,c1802B,c1902B,c1A02B,c1B02B,c1C02B,c1D02B,c1E02B,c1F02B;
wire signed [4:0] c1010B,c1110B,c1210B,c1310B,c1410B,c1510B,c1610B,c1710B,c1810B,c1910B,c1A10B,c1B10B,c1C10B,c1D10B,c1E10B,c1F10B;
wire signed [4:0] c1011B,c1111B,c1211B,c1311B,c1411B,c1511B,c1611B,c1711B,c1811B,c1911B,c1A11B,c1B11B,c1C11B,c1D11B,c1E11B,c1F11B;
wire signed [4:0] c1012B,c1112B,c1212B,c1312B,c1412B,c1512B,c1612B,c1712B,c1812B,c1912B,c1A12B,c1B12B,c1C12B,c1D12B,c1E12B,c1F12B;
wire signed [4:0] c1020B,c1120B,c1220B,c1320B,c1420B,c1520B,c1620B,c1720B,c1820B,c1920B,c1A20B,c1B20B,c1C20B,c1D20B,c1E20B,c1F20B;
wire signed [4:0] c1021B,c1121B,c1221B,c1321B,c1421B,c1521B,c1621B,c1721B,c1821B,c1921B,c1A21B,c1B21B,c1C21B,c1D21B,c1E21B,c1F21B;
wire signed [4:0] c1022B,c1122B,c1222B,c1322B,c1422B,c1522B,c1622B,c1722B,c1822B,c1922B,c1A22B,c1B22B,c1C22B,c1D22B,c1E22B,c1F22B;
wire signed [4:0] c1000C,c1100C,c1200C,c1300C,c1400C,c1500C,c1600C,c1700C,c1800C,c1900C,c1A00C,c1B00C,c1C00C,c1D00C,c1E00C,c1F00C;
wire signed [4:0] c1001C,c1101C,c1201C,c1301C,c1401C,c1501C,c1601C,c1701C,c1801C,c1901C,c1A01C,c1B01C,c1C01C,c1D01C,c1E01C,c1F01C;
wire signed [4:0] c1002C,c1102C,c1202C,c1302C,c1402C,c1502C,c1602C,c1702C,c1802C,c1902C,c1A02C,c1B02C,c1C02C,c1D02C,c1E02C,c1F02C;
wire signed [4:0] c1010C,c1110C,c1210C,c1310C,c1410C,c1510C,c1610C,c1710C,c1810C,c1910C,c1A10C,c1B10C,c1C10C,c1D10C,c1E10C,c1F10C;
wire signed [4:0] c1011C,c1111C,c1211C,c1311C,c1411C,c1511C,c1611C,c1711C,c1811C,c1911C,c1A11C,c1B11C,c1C11C,c1D11C,c1E11C,c1F11C;
wire signed [4:0] c1012C,c1112C,c1212C,c1312C,c1412C,c1512C,c1612C,c1712C,c1812C,c1912C,c1A12C,c1B12C,c1C12C,c1D12C,c1E12C,c1F12C;
wire signed [4:0] c1020C,c1120C,c1220C,c1320C,c1420C,c1520C,c1620C,c1720C,c1820C,c1920C,c1A20C,c1B20C,c1C20C,c1D20C,c1E20C,c1F20C;
wire signed [4:0] c1021C,c1121C,c1221C,c1321C,c1421C,c1521C,c1621C,c1721C,c1821C,c1921C,c1A21C,c1B21C,c1C21C,c1D21C,c1E21C,c1F21C;
wire signed [4:0] c1022C,c1122C,c1222C,c1322C,c1422C,c1522C,c1622C,c1722C,c1822C,c1922C,c1A22C,c1B22C,c1C22C,c1D22C,c1E22C,c1F22C;
wire signed [4:0] c1000D,c1100D,c1200D,c1300D,c1400D,c1500D,c1600D,c1700D,c1800D,c1900D,c1A00D,c1B00D,c1C00D,c1D00D,c1E00D,c1F00D;
wire signed [4:0] c1001D,c1101D,c1201D,c1301D,c1401D,c1501D,c1601D,c1701D,c1801D,c1901D,c1A01D,c1B01D,c1C01D,c1D01D,c1E01D,c1F01D;
wire signed [4:0] c1002D,c1102D,c1202D,c1302D,c1402D,c1502D,c1602D,c1702D,c1802D,c1902D,c1A02D,c1B02D,c1C02D,c1D02D,c1E02D,c1F02D;
wire signed [4:0] c1010D,c1110D,c1210D,c1310D,c1410D,c1510D,c1610D,c1710D,c1810D,c1910D,c1A10D,c1B10D,c1C10D,c1D10D,c1E10D,c1F10D;
wire signed [4:0] c1011D,c1111D,c1211D,c1311D,c1411D,c1511D,c1611D,c1711D,c1811D,c1911D,c1A11D,c1B11D,c1C11D,c1D11D,c1E11D,c1F11D;
wire signed [4:0] c1012D,c1112D,c1212D,c1312D,c1412D,c1512D,c1612D,c1712D,c1812D,c1912D,c1A12D,c1B12D,c1C12D,c1D12D,c1E12D,c1F12D;
wire signed [4:0] c1020D,c1120D,c1220D,c1320D,c1420D,c1520D,c1620D,c1720D,c1820D,c1920D,c1A20D,c1B20D,c1C20D,c1D20D,c1E20D,c1F20D;
wire signed [4:0] c1021D,c1121D,c1221D,c1321D,c1421D,c1521D,c1621D,c1721D,c1821D,c1921D,c1A21D,c1B21D,c1C21D,c1D21D,c1E21D,c1F21D;
wire signed [4:0] c1022D,c1122D,c1222D,c1322D,c1422D,c1522D,c1622D,c1722D,c1822D,c1922D,c1A22D,c1B22D,c1C22D,c1D22D,c1E22D,c1F22D;
wire signed [4:0] c1000E,c1100E,c1200E,c1300E,c1400E,c1500E,c1600E,c1700E,c1800E,c1900E,c1A00E,c1B00E,c1C00E,c1D00E,c1E00E,c1F00E;
wire signed [4:0] c1001E,c1101E,c1201E,c1301E,c1401E,c1501E,c1601E,c1701E,c1801E,c1901E,c1A01E,c1B01E,c1C01E,c1D01E,c1E01E,c1F01E;
wire signed [4:0] c1002E,c1102E,c1202E,c1302E,c1402E,c1502E,c1602E,c1702E,c1802E,c1902E,c1A02E,c1B02E,c1C02E,c1D02E,c1E02E,c1F02E;
wire signed [4:0] c1010E,c1110E,c1210E,c1310E,c1410E,c1510E,c1610E,c1710E,c1810E,c1910E,c1A10E,c1B10E,c1C10E,c1D10E,c1E10E,c1F10E;
wire signed [4:0] c1011E,c1111E,c1211E,c1311E,c1411E,c1511E,c1611E,c1711E,c1811E,c1911E,c1A11E,c1B11E,c1C11E,c1D11E,c1E11E,c1F11E;
wire signed [4:0] c1012E,c1112E,c1212E,c1312E,c1412E,c1512E,c1612E,c1712E,c1812E,c1912E,c1A12E,c1B12E,c1C12E,c1D12E,c1E12E,c1F12E;
wire signed [4:0] c1020E,c1120E,c1220E,c1320E,c1420E,c1520E,c1620E,c1720E,c1820E,c1920E,c1A20E,c1B20E,c1C20E,c1D20E,c1E20E,c1F20E;
wire signed [4:0] c1021E,c1121E,c1221E,c1321E,c1421E,c1521E,c1621E,c1721E,c1821E,c1921E,c1A21E,c1B21E,c1C21E,c1D21E,c1E21E,c1F21E;
wire signed [4:0] c1022E,c1122E,c1222E,c1322E,c1422E,c1522E,c1622E,c1722E,c1822E,c1922E,c1A22E,c1B22E,c1C22E,c1D22E,c1E22E,c1F22E;
wire signed [4:0] c1000F,c1100F,c1200F,c1300F,c1400F,c1500F,c1600F,c1700F,c1800F,c1900F,c1A00F,c1B00F,c1C00F,c1D00F,c1E00F,c1F00F;
wire signed [4:0] c1001F,c1101F,c1201F,c1301F,c1401F,c1501F,c1601F,c1701F,c1801F,c1901F,c1A01F,c1B01F,c1C01F,c1D01F,c1E01F,c1F01F;
wire signed [4:0] c1002F,c1102F,c1202F,c1302F,c1402F,c1502F,c1602F,c1702F,c1802F,c1902F,c1A02F,c1B02F,c1C02F,c1D02F,c1E02F,c1F02F;
wire signed [4:0] c1010F,c1110F,c1210F,c1310F,c1410F,c1510F,c1610F,c1710F,c1810F,c1910F,c1A10F,c1B10F,c1C10F,c1D10F,c1E10F,c1F10F;
wire signed [4:0] c1011F,c1111F,c1211F,c1311F,c1411F,c1511F,c1611F,c1711F,c1811F,c1911F,c1A11F,c1B11F,c1C11F,c1D11F,c1E11F,c1F11F;
wire signed [4:0] c1012F,c1112F,c1212F,c1312F,c1412F,c1512F,c1612F,c1712F,c1812F,c1912F,c1A12F,c1B12F,c1C12F,c1D12F,c1E12F,c1F12F;
wire signed [4:0] c1020F,c1120F,c1220F,c1320F,c1420F,c1520F,c1620F,c1720F,c1820F,c1920F,c1A20F,c1B20F,c1C20F,c1D20F,c1E20F,c1F20F;
wire signed [4:0] c1021F,c1121F,c1221F,c1321F,c1421F,c1521F,c1621F,c1721F,c1821F,c1921F,c1A21F,c1B21F,c1C21F,c1D21F,c1E21F,c1F21F;
wire signed [4:0] c1022F,c1122F,c1222F,c1322F,c1422F,c1522F,c1622F,c1722F,c1822F,c1922F,c1A22F,c1B22F,c1C22F,c1D22F,c1E22F,c1F22F;
wire signed [4:0] c1000G,c1100G,c1200G,c1300G,c1400G,c1500G,c1600G,c1700G,c1800G,c1900G,c1A00G,c1B00G,c1C00G,c1D00G,c1E00G,c1F00G;
wire signed [4:0] c1001G,c1101G,c1201G,c1301G,c1401G,c1501G,c1601G,c1701G,c1801G,c1901G,c1A01G,c1B01G,c1C01G,c1D01G,c1E01G,c1F01G;
wire signed [4:0] c1002G,c1102G,c1202G,c1302G,c1402G,c1502G,c1602G,c1702G,c1802G,c1902G,c1A02G,c1B02G,c1C02G,c1D02G,c1E02G,c1F02G;
wire signed [4:0] c1010G,c1110G,c1210G,c1310G,c1410G,c1510G,c1610G,c1710G,c1810G,c1910G,c1A10G,c1B10G,c1C10G,c1D10G,c1E10G,c1F10G;
wire signed [4:0] c1011G,c1111G,c1211G,c1311G,c1411G,c1511G,c1611G,c1711G,c1811G,c1911G,c1A11G,c1B11G,c1C11G,c1D11G,c1E11G,c1F11G;
wire signed [4:0] c1012G,c1112G,c1212G,c1312G,c1412G,c1512G,c1612G,c1712G,c1812G,c1912G,c1A12G,c1B12G,c1C12G,c1D12G,c1E12G,c1F12G;
wire signed [4:0] c1020G,c1120G,c1220G,c1320G,c1420G,c1520G,c1620G,c1720G,c1820G,c1920G,c1A20G,c1B20G,c1C20G,c1D20G,c1E20G,c1F20G;
wire signed [4:0] c1021G,c1121G,c1221G,c1321G,c1421G,c1521G,c1621G,c1721G,c1821G,c1921G,c1A21G,c1B21G,c1C21G,c1D21G,c1E21G,c1F21G;
wire signed [4:0] c1022G,c1122G,c1222G,c1322G,c1422G,c1522G,c1622G,c1722G,c1822G,c1922G,c1A22G,c1B22G,c1C22G,c1D22G,c1E22G,c1F22G;
wire signed [4:0] c1000H,c1100H,c1200H,c1300H,c1400H,c1500H,c1600H,c1700H,c1800H,c1900H,c1A00H,c1B00H,c1C00H,c1D00H,c1E00H,c1F00H;
wire signed [4:0] c1001H,c1101H,c1201H,c1301H,c1401H,c1501H,c1601H,c1701H,c1801H,c1901H,c1A01H,c1B01H,c1C01H,c1D01H,c1E01H,c1F01H;
wire signed [4:0] c1002H,c1102H,c1202H,c1302H,c1402H,c1502H,c1602H,c1702H,c1802H,c1902H,c1A02H,c1B02H,c1C02H,c1D02H,c1E02H,c1F02H;
wire signed [4:0] c1010H,c1110H,c1210H,c1310H,c1410H,c1510H,c1610H,c1710H,c1810H,c1910H,c1A10H,c1B10H,c1C10H,c1D10H,c1E10H,c1F10H;
wire signed [4:0] c1011H,c1111H,c1211H,c1311H,c1411H,c1511H,c1611H,c1711H,c1811H,c1911H,c1A11H,c1B11H,c1C11H,c1D11H,c1E11H,c1F11H;
wire signed [4:0] c1012H,c1112H,c1212H,c1312H,c1412H,c1512H,c1612H,c1712H,c1812H,c1912H,c1A12H,c1B12H,c1C12H,c1D12H,c1E12H,c1F12H;
wire signed [4:0] c1020H,c1120H,c1220H,c1320H,c1420H,c1520H,c1620H,c1720H,c1820H,c1920H,c1A20H,c1B20H,c1C20H,c1D20H,c1E20H,c1F20H;
wire signed [4:0] c1021H,c1121H,c1221H,c1321H,c1421H,c1521H,c1621H,c1721H,c1821H,c1921H,c1A21H,c1B21H,c1C21H,c1D21H,c1E21H,c1F21H;
wire signed [4:0] c1022H,c1122H,c1222H,c1322H,c1422H,c1522H,c1622H,c1722H,c1822H,c1922H,c1A22H,c1B22H,c1C22H,c1D22H,c1E22H,c1F22H;
wire signed [4:0] c1000I,c1100I,c1200I,c1300I,c1400I,c1500I,c1600I,c1700I,c1800I,c1900I,c1A00I,c1B00I,c1C00I,c1D00I,c1E00I,c1F00I;
wire signed [4:0] c1001I,c1101I,c1201I,c1301I,c1401I,c1501I,c1601I,c1701I,c1801I,c1901I,c1A01I,c1B01I,c1C01I,c1D01I,c1E01I,c1F01I;
wire signed [4:0] c1002I,c1102I,c1202I,c1302I,c1402I,c1502I,c1602I,c1702I,c1802I,c1902I,c1A02I,c1B02I,c1C02I,c1D02I,c1E02I,c1F02I;
wire signed [4:0] c1010I,c1110I,c1210I,c1310I,c1410I,c1510I,c1610I,c1710I,c1810I,c1910I,c1A10I,c1B10I,c1C10I,c1D10I,c1E10I,c1F10I;
wire signed [4:0] c1011I,c1111I,c1211I,c1311I,c1411I,c1511I,c1611I,c1711I,c1811I,c1911I,c1A11I,c1B11I,c1C11I,c1D11I,c1E11I,c1F11I;
wire signed [4:0] c1012I,c1112I,c1212I,c1312I,c1412I,c1512I,c1612I,c1712I,c1812I,c1912I,c1A12I,c1B12I,c1C12I,c1D12I,c1E12I,c1F12I;
wire signed [4:0] c1020I,c1120I,c1220I,c1320I,c1420I,c1520I,c1620I,c1720I,c1820I,c1920I,c1A20I,c1B20I,c1C20I,c1D20I,c1E20I,c1F20I;
wire signed [4:0] c1021I,c1121I,c1221I,c1321I,c1421I,c1521I,c1621I,c1721I,c1821I,c1921I,c1A21I,c1B21I,c1C21I,c1D21I,c1E21I,c1F21I;
wire signed [4:0] c1022I,c1122I,c1222I,c1322I,c1422I,c1522I,c1622I,c1722I,c1822I,c1922I,c1A22I,c1B22I,c1C22I,c1D22I,c1E22I,c1F22I;
wire signed [4:0] c1000J,c1100J,c1200J,c1300J,c1400J,c1500J,c1600J,c1700J,c1800J,c1900J,c1A00J,c1B00J,c1C00J,c1D00J,c1E00J,c1F00J;
wire signed [4:0] c1001J,c1101J,c1201J,c1301J,c1401J,c1501J,c1601J,c1701J,c1801J,c1901J,c1A01J,c1B01J,c1C01J,c1D01J,c1E01J,c1F01J;
wire signed [4:0] c1002J,c1102J,c1202J,c1302J,c1402J,c1502J,c1602J,c1702J,c1802J,c1902J,c1A02J,c1B02J,c1C02J,c1D02J,c1E02J,c1F02J;
wire signed [4:0] c1010J,c1110J,c1210J,c1310J,c1410J,c1510J,c1610J,c1710J,c1810J,c1910J,c1A10J,c1B10J,c1C10J,c1D10J,c1E10J,c1F10J;
wire signed [4:0] c1011J,c1111J,c1211J,c1311J,c1411J,c1511J,c1611J,c1711J,c1811J,c1911J,c1A11J,c1B11J,c1C11J,c1D11J,c1E11J,c1F11J;
wire signed [4:0] c1012J,c1112J,c1212J,c1312J,c1412J,c1512J,c1612J,c1712J,c1812J,c1912J,c1A12J,c1B12J,c1C12J,c1D12J,c1E12J,c1F12J;
wire signed [4:0] c1020J,c1120J,c1220J,c1320J,c1420J,c1520J,c1620J,c1720J,c1820J,c1920J,c1A20J,c1B20J,c1C20J,c1D20J,c1E20J,c1F20J;
wire signed [4:0] c1021J,c1121J,c1221J,c1321J,c1421J,c1521J,c1621J,c1721J,c1821J,c1921J,c1A21J,c1B21J,c1C21J,c1D21J,c1E21J,c1F21J;
wire signed [4:0] c1022J,c1122J,c1222J,c1322J,c1422J,c1522J,c1622J,c1722J,c1822J,c1922J,c1A22J,c1B22J,c1C22J,c1D22J,c1E22J,c1F22J;
wire signed [4:0] c1000K,c1100K,c1200K,c1300K,c1400K,c1500K,c1600K,c1700K,c1800K,c1900K,c1A00K,c1B00K,c1C00K,c1D00K,c1E00K,c1F00K;
wire signed [4:0] c1001K,c1101K,c1201K,c1301K,c1401K,c1501K,c1601K,c1701K,c1801K,c1901K,c1A01K,c1B01K,c1C01K,c1D01K,c1E01K,c1F01K;
wire signed [4:0] c1002K,c1102K,c1202K,c1302K,c1402K,c1502K,c1602K,c1702K,c1802K,c1902K,c1A02K,c1B02K,c1C02K,c1D02K,c1E02K,c1F02K;
wire signed [4:0] c1010K,c1110K,c1210K,c1310K,c1410K,c1510K,c1610K,c1710K,c1810K,c1910K,c1A10K,c1B10K,c1C10K,c1D10K,c1E10K,c1F10K;
wire signed [4:0] c1011K,c1111K,c1211K,c1311K,c1411K,c1511K,c1611K,c1711K,c1811K,c1911K,c1A11K,c1B11K,c1C11K,c1D11K,c1E11K,c1F11K;
wire signed [4:0] c1012K,c1112K,c1212K,c1312K,c1412K,c1512K,c1612K,c1712K,c1812K,c1912K,c1A12K,c1B12K,c1C12K,c1D12K,c1E12K,c1F12K;
wire signed [4:0] c1020K,c1120K,c1220K,c1320K,c1420K,c1520K,c1620K,c1720K,c1820K,c1920K,c1A20K,c1B20K,c1C20K,c1D20K,c1E20K,c1F20K;
wire signed [4:0] c1021K,c1121K,c1221K,c1321K,c1421K,c1521K,c1621K,c1721K,c1821K,c1921K,c1A21K,c1B21K,c1C21K,c1D21K,c1E21K,c1F21K;
wire signed [4:0] c1022K,c1122K,c1222K,c1322K,c1422K,c1522K,c1622K,c1722K,c1822K,c1922K,c1A22K,c1B22K,c1C22K,c1D22K,c1E22K,c1F22K;
wire signed [4:0] c1000L,c1100L,c1200L,c1300L,c1400L,c1500L,c1600L,c1700L,c1800L,c1900L,c1A00L,c1B00L,c1C00L,c1D00L,c1E00L,c1F00L;
wire signed [4:0] c1001L,c1101L,c1201L,c1301L,c1401L,c1501L,c1601L,c1701L,c1801L,c1901L,c1A01L,c1B01L,c1C01L,c1D01L,c1E01L,c1F01L;
wire signed [4:0] c1002L,c1102L,c1202L,c1302L,c1402L,c1502L,c1602L,c1702L,c1802L,c1902L,c1A02L,c1B02L,c1C02L,c1D02L,c1E02L,c1F02L;
wire signed [4:0] c1010L,c1110L,c1210L,c1310L,c1410L,c1510L,c1610L,c1710L,c1810L,c1910L,c1A10L,c1B10L,c1C10L,c1D10L,c1E10L,c1F10L;
wire signed [4:0] c1011L,c1111L,c1211L,c1311L,c1411L,c1511L,c1611L,c1711L,c1811L,c1911L,c1A11L,c1B11L,c1C11L,c1D11L,c1E11L,c1F11L;
wire signed [4:0] c1012L,c1112L,c1212L,c1312L,c1412L,c1512L,c1612L,c1712L,c1812L,c1912L,c1A12L,c1B12L,c1C12L,c1D12L,c1E12L,c1F12L;
wire signed [4:0] c1020L,c1120L,c1220L,c1320L,c1420L,c1520L,c1620L,c1720L,c1820L,c1920L,c1A20L,c1B20L,c1C20L,c1D20L,c1E20L,c1F20L;
wire signed [4:0] c1021L,c1121L,c1221L,c1321L,c1421L,c1521L,c1621L,c1721L,c1821L,c1921L,c1A21L,c1B21L,c1C21L,c1D21L,c1E21L,c1F21L;
wire signed [4:0] c1022L,c1122L,c1222L,c1322L,c1422L,c1522L,c1622L,c1722L,c1822L,c1922L,c1A22L,c1B22L,c1C22L,c1D22L,c1E22L,c1F22L;
wire signed [4:0] c1000M,c1100M,c1200M,c1300M,c1400M,c1500M,c1600M,c1700M,c1800M,c1900M,c1A00M,c1B00M,c1C00M,c1D00M,c1E00M,c1F00M;
wire signed [4:0] c1001M,c1101M,c1201M,c1301M,c1401M,c1501M,c1601M,c1701M,c1801M,c1901M,c1A01M,c1B01M,c1C01M,c1D01M,c1E01M,c1F01M;
wire signed [4:0] c1002M,c1102M,c1202M,c1302M,c1402M,c1502M,c1602M,c1702M,c1802M,c1902M,c1A02M,c1B02M,c1C02M,c1D02M,c1E02M,c1F02M;
wire signed [4:0] c1010M,c1110M,c1210M,c1310M,c1410M,c1510M,c1610M,c1710M,c1810M,c1910M,c1A10M,c1B10M,c1C10M,c1D10M,c1E10M,c1F10M;
wire signed [4:0] c1011M,c1111M,c1211M,c1311M,c1411M,c1511M,c1611M,c1711M,c1811M,c1911M,c1A11M,c1B11M,c1C11M,c1D11M,c1E11M,c1F11M;
wire signed [4:0] c1012M,c1112M,c1212M,c1312M,c1412M,c1512M,c1612M,c1712M,c1812M,c1912M,c1A12M,c1B12M,c1C12M,c1D12M,c1E12M,c1F12M;
wire signed [4:0] c1020M,c1120M,c1220M,c1320M,c1420M,c1520M,c1620M,c1720M,c1820M,c1920M,c1A20M,c1B20M,c1C20M,c1D20M,c1E20M,c1F20M;
wire signed [4:0] c1021M,c1121M,c1221M,c1321M,c1421M,c1521M,c1621M,c1721M,c1821M,c1921M,c1A21M,c1B21M,c1C21M,c1D21M,c1E21M,c1F21M;
wire signed [4:0] c1022M,c1122M,c1222M,c1322M,c1422M,c1522M,c1622M,c1722M,c1822M,c1922M,c1A22M,c1B22M,c1C22M,c1D22M,c1E22M,c1F22M;
wire signed [8:0] C1000;
wire A1000;
wire signed [8:0] C1010;
wire A1010;
wire signed [8:0] C1020;
wire A1020;
wire signed [8:0] C1100;
wire A1100;
wire signed [8:0] C1110;
wire A1110;
wire signed [8:0] C1120;
wire A1120;
wire signed [8:0] C1200;
wire A1200;
wire signed [8:0] C1210;
wire A1210;
wire signed [8:0] C1220;
wire A1220;
wire signed [8:0] C1001;
wire A1001;
wire signed [8:0] C1011;
wire A1011;
wire signed [8:0] C1021;
wire A1021;
wire signed [8:0] C1101;
wire A1101;
wire signed [8:0] C1111;
wire A1111;
wire signed [8:0] C1121;
wire A1121;
wire signed [8:0] C1201;
wire A1201;
wire signed [8:0] C1211;
wire A1211;
wire signed [8:0] C1221;
wire A1221;
wire signed [8:0] C1002;
wire A1002;
wire signed [8:0] C1012;
wire A1012;
wire signed [8:0] C1022;
wire A1022;
wire signed [8:0] C1102;
wire A1102;
wire signed [8:0] C1112;
wire A1112;
wire signed [8:0] C1122;
wire A1122;
wire signed [8:0] C1202;
wire A1202;
wire signed [8:0] C1212;
wire A1212;
wire signed [8:0] C1222;
wire A1222;
wire signed [8:0] C1003;
wire A1003;
wire signed [8:0] C1013;
wire A1013;
wire signed [8:0] C1023;
wire A1023;
wire signed [8:0] C1103;
wire A1103;
wire signed [8:0] C1113;
wire A1113;
wire signed [8:0] C1123;
wire A1123;
wire signed [8:0] C1203;
wire A1203;
wire signed [8:0] C1213;
wire A1213;
wire signed [8:0] C1223;
wire A1223;
wire signed [8:0] C1004;
wire A1004;
wire signed [8:0] C1014;
wire A1014;
wire signed [8:0] C1024;
wire A1024;
wire signed [8:0] C1104;
wire A1104;
wire signed [8:0] C1114;
wire A1114;
wire signed [8:0] C1124;
wire A1124;
wire signed [8:0] C1204;
wire A1204;
wire signed [8:0] C1214;
wire A1214;
wire signed [8:0] C1224;
wire A1224;
wire signed [8:0] C1005;
wire A1005;
wire signed [8:0] C1015;
wire A1015;
wire signed [8:0] C1025;
wire A1025;
wire signed [8:0] C1105;
wire A1105;
wire signed [8:0] C1115;
wire A1115;
wire signed [8:0] C1125;
wire A1125;
wire signed [8:0] C1205;
wire A1205;
wire signed [8:0] C1215;
wire A1215;
wire signed [8:0] C1225;
wire A1225;
wire signed [8:0] C1006;
wire A1006;
wire signed [8:0] C1016;
wire A1016;
wire signed [8:0] C1026;
wire A1026;
wire signed [8:0] C1106;
wire A1106;
wire signed [8:0] C1116;
wire A1116;
wire signed [8:0] C1126;
wire A1126;
wire signed [8:0] C1206;
wire A1206;
wire signed [8:0] C1216;
wire A1216;
wire signed [8:0] C1226;
wire A1226;
wire signed [8:0] C1007;
wire A1007;
wire signed [8:0] C1017;
wire A1017;
wire signed [8:0] C1027;
wire A1027;
wire signed [8:0] C1107;
wire A1107;
wire signed [8:0] C1117;
wire A1117;
wire signed [8:0] C1127;
wire A1127;
wire signed [8:0] C1207;
wire A1207;
wire signed [8:0] C1217;
wire A1217;
wire signed [8:0] C1227;
wire A1227;
wire signed [8:0] C1008;
wire A1008;
wire signed [8:0] C1018;
wire A1018;
wire signed [8:0] C1028;
wire A1028;
wire signed [8:0] C1108;
wire A1108;
wire signed [8:0] C1118;
wire A1118;
wire signed [8:0] C1128;
wire A1128;
wire signed [8:0] C1208;
wire A1208;
wire signed [8:0] C1218;
wire A1218;
wire signed [8:0] C1228;
wire A1228;
wire signed [8:0] C1009;
wire A1009;
wire signed [8:0] C1019;
wire A1019;
wire signed [8:0] C1029;
wire A1029;
wire signed [8:0] C1109;
wire A1109;
wire signed [8:0] C1119;
wire A1119;
wire signed [8:0] C1129;
wire A1129;
wire signed [8:0] C1209;
wire A1209;
wire signed [8:0] C1219;
wire A1219;
wire signed [8:0] C1229;
wire A1229;
wire signed [8:0] C100A;
wire A100A;
wire signed [8:0] C101A;
wire A101A;
wire signed [8:0] C102A;
wire A102A;
wire signed [8:0] C110A;
wire A110A;
wire signed [8:0] C111A;
wire A111A;
wire signed [8:0] C112A;
wire A112A;
wire signed [8:0] C120A;
wire A120A;
wire signed [8:0] C121A;
wire A121A;
wire signed [8:0] C122A;
wire A122A;
wire signed [8:0] C100B;
wire A100B;
wire signed [8:0] C101B;
wire A101B;
wire signed [8:0] C102B;
wire A102B;
wire signed [8:0] C110B;
wire A110B;
wire signed [8:0] C111B;
wire A111B;
wire signed [8:0] C112B;
wire A112B;
wire signed [8:0] C120B;
wire A120B;
wire signed [8:0] C121B;
wire A121B;
wire signed [8:0] C122B;
wire A122B;
wire signed [8:0] C100C;
wire A100C;
wire signed [8:0] C101C;
wire A101C;
wire signed [8:0] C102C;
wire A102C;
wire signed [8:0] C110C;
wire A110C;
wire signed [8:0] C111C;
wire A111C;
wire signed [8:0] C112C;
wire A112C;
wire signed [8:0] C120C;
wire A120C;
wire signed [8:0] C121C;
wire A121C;
wire signed [8:0] C122C;
wire A122C;
wire signed [8:0] C100D;
wire A100D;
wire signed [8:0] C101D;
wire A101D;
wire signed [8:0] C102D;
wire A102D;
wire signed [8:0] C110D;
wire A110D;
wire signed [8:0] C111D;
wire A111D;
wire signed [8:0] C112D;
wire A112D;
wire signed [8:0] C120D;
wire A120D;
wire signed [8:0] C121D;
wire A121D;
wire signed [8:0] C122D;
wire A122D;
wire signed [8:0] C100E;
wire A100E;
wire signed [8:0] C101E;
wire A101E;
wire signed [8:0] C102E;
wire A102E;
wire signed [8:0] C110E;
wire A110E;
wire signed [8:0] C111E;
wire A111E;
wire signed [8:0] C112E;
wire A112E;
wire signed [8:0] C120E;
wire A120E;
wire signed [8:0] C121E;
wire A121E;
wire signed [8:0] C122E;
wire A122E;
wire signed [8:0] C100F;
wire A100F;
wire signed [8:0] C101F;
wire A101F;
wire signed [8:0] C102F;
wire A102F;
wire signed [8:0] C110F;
wire A110F;
wire signed [8:0] C111F;
wire A111F;
wire signed [8:0] C112F;
wire A112F;
wire signed [8:0] C120F;
wire A120F;
wire signed [8:0] C121F;
wire A121F;
wire signed [8:0] C122F;
wire A122F;
wire signed [8:0] C100G;
wire A100G;
wire signed [8:0] C101G;
wire A101G;
wire signed [8:0] C102G;
wire A102G;
wire signed [8:0] C110G;
wire A110G;
wire signed [8:0] C111G;
wire A111G;
wire signed [8:0] C112G;
wire A112G;
wire signed [8:0] C120G;
wire A120G;
wire signed [8:0] C121G;
wire A121G;
wire signed [8:0] C122G;
wire A122G;
wire signed [8:0] C100H;
wire A100H;
wire signed [8:0] C101H;
wire A101H;
wire signed [8:0] C102H;
wire A102H;
wire signed [8:0] C110H;
wire A110H;
wire signed [8:0] C111H;
wire A111H;
wire signed [8:0] C112H;
wire A112H;
wire signed [8:0] C120H;
wire A120H;
wire signed [8:0] C121H;
wire A121H;
wire signed [8:0] C122H;
wire A122H;
wire signed [8:0] C100I;
wire A100I;
wire signed [8:0] C101I;
wire A101I;
wire signed [8:0] C102I;
wire A102I;
wire signed [8:0] C110I;
wire A110I;
wire signed [8:0] C111I;
wire A111I;
wire signed [8:0] C112I;
wire A112I;
wire signed [8:0] C120I;
wire A120I;
wire signed [8:0] C121I;
wire A121I;
wire signed [8:0] C122I;
wire A122I;
wire signed [8:0] C100J;
wire A100J;
wire signed [8:0] C101J;
wire A101J;
wire signed [8:0] C102J;
wire A102J;
wire signed [8:0] C110J;
wire A110J;
wire signed [8:0] C111J;
wire A111J;
wire signed [8:0] C112J;
wire A112J;
wire signed [8:0] C120J;
wire A120J;
wire signed [8:0] C121J;
wire A121J;
wire signed [8:0] C122J;
wire A122J;
wire signed [8:0] C100K;
wire A100K;
wire signed [8:0] C101K;
wire A101K;
wire signed [8:0] C102K;
wire A102K;
wire signed [8:0] C110K;
wire A110K;
wire signed [8:0] C111K;
wire A111K;
wire signed [8:0] C112K;
wire A112K;
wire signed [8:0] C120K;
wire A120K;
wire signed [8:0] C121K;
wire A121K;
wire signed [8:0] C122K;
wire A122K;
wire signed [8:0] C100L;
wire A100L;
wire signed [8:0] C101L;
wire A101L;
wire signed [8:0] C102L;
wire A102L;
wire signed [8:0] C110L;
wire A110L;
wire signed [8:0] C111L;
wire A111L;
wire signed [8:0] C112L;
wire A112L;
wire signed [8:0] C120L;
wire A120L;
wire signed [8:0] C121L;
wire A121L;
wire signed [8:0] C122L;
wire A122L;
wire signed [8:0] C100M;
wire A100M;
wire signed [8:0] C101M;
wire A101M;
wire signed [8:0] C102M;
wire A102M;
wire signed [8:0] C110M;
wire A110M;
wire signed [8:0] C111M;
wire A111M;
wire signed [8:0] C112M;
wire A112M;
wire signed [8:0] C120M;
wire A120M;
wire signed [8:0] C121M;
wire A121M;
wire signed [8:0] C122M;
wire A122M;
DFF_save_fm DFF_W432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10000));
DFF_save_fm DFF_W433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10010));
DFF_save_fm DFF_W434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10020));
DFF_save_fm DFF_W435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10100));
DFF_save_fm DFF_W436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10110));
DFF_save_fm DFF_W437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10120));
DFF_save_fm DFF_W438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10200));
DFF_save_fm DFF_W439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10210));
DFF_save_fm DFF_W440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10220));
DFF_save_fm DFF_W441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10001));
DFF_save_fm DFF_W442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10011));
DFF_save_fm DFF_W443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10021));
DFF_save_fm DFF_W444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10101));
DFF_save_fm DFF_W445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10111));
DFF_save_fm DFF_W446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10121));
DFF_save_fm DFF_W447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10201));
DFF_save_fm DFF_W448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10211));
DFF_save_fm DFF_W449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10221));
DFF_save_fm DFF_W450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10002));
DFF_save_fm DFF_W451(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10012));
DFF_save_fm DFF_W452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10022));
DFF_save_fm DFF_W453(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10102));
DFF_save_fm DFF_W454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10112));
DFF_save_fm DFF_W455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10122));
DFF_save_fm DFF_W456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10202));
DFF_save_fm DFF_W457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10212));
DFF_save_fm DFF_W458(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10222));
DFF_save_fm DFF_W459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10003));
DFF_save_fm DFF_W460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10013));
DFF_save_fm DFF_W461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10023));
DFF_save_fm DFF_W462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10103));
DFF_save_fm DFF_W463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10113));
DFF_save_fm DFF_W464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10123));
DFF_save_fm DFF_W465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10203));
DFF_save_fm DFF_W466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10213));
DFF_save_fm DFF_W467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10223));
DFF_save_fm DFF_W468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10004));
DFF_save_fm DFF_W469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10014));
DFF_save_fm DFF_W470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10024));
DFF_save_fm DFF_W471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10104));
DFF_save_fm DFF_W472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10114));
DFF_save_fm DFF_W473(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10124));
DFF_save_fm DFF_W474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10204));
DFF_save_fm DFF_W475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10214));
DFF_save_fm DFF_W476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10224));
DFF_save_fm DFF_W477(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10005));
DFF_save_fm DFF_W478(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10015));
DFF_save_fm DFF_W479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10025));
DFF_save_fm DFF_W480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10105));
DFF_save_fm DFF_W481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10115));
DFF_save_fm DFF_W482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10125));
DFF_save_fm DFF_W483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10205));
DFF_save_fm DFF_W484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10215));
DFF_save_fm DFF_W485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10225));
DFF_save_fm DFF_W486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10006));
DFF_save_fm DFF_W487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10016));
DFF_save_fm DFF_W488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10026));
DFF_save_fm DFF_W489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10106));
DFF_save_fm DFF_W490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10116));
DFF_save_fm DFF_W491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10126));
DFF_save_fm DFF_W492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10206));
DFF_save_fm DFF_W493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10216));
DFF_save_fm DFF_W494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10226));
DFF_save_fm DFF_W495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10007));
DFF_save_fm DFF_W496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10017));
DFF_save_fm DFF_W497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10027));
DFF_save_fm DFF_W498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10107));
DFF_save_fm DFF_W499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10117));
DFF_save_fm DFF_W500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10127));
DFF_save_fm DFF_W501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10207));
DFF_save_fm DFF_W502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10217));
DFF_save_fm DFF_W503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10227));
DFF_save_fm DFF_W504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10008));
DFF_save_fm DFF_W505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10018));
DFF_save_fm DFF_W506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10028));
DFF_save_fm DFF_W507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10108));
DFF_save_fm DFF_W508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10118));
DFF_save_fm DFF_W509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10128));
DFF_save_fm DFF_W510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10208));
DFF_save_fm DFF_W511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10218));
DFF_save_fm DFF_W512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10228));
DFF_save_fm DFF_W513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10009));
DFF_save_fm DFF_W514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10019));
DFF_save_fm DFF_W515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10029));
DFF_save_fm DFF_W516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10109));
DFF_save_fm DFF_W517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10119));
DFF_save_fm DFF_W518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10129));
DFF_save_fm DFF_W519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10209));
DFF_save_fm DFF_W520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10219));
DFF_save_fm DFF_W521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10229));
DFF_save_fm DFF_W522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1000A));
DFF_save_fm DFF_W523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1001A));
DFF_save_fm DFF_W524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1002A));
DFF_save_fm DFF_W525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1010A));
DFF_save_fm DFF_W526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1011A));
DFF_save_fm DFF_W527(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1012A));
DFF_save_fm DFF_W528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1020A));
DFF_save_fm DFF_W529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1021A));
DFF_save_fm DFF_W530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1022A));
DFF_save_fm DFF_W531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1000B));
DFF_save_fm DFF_W532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1001B));
DFF_save_fm DFF_W533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1002B));
DFF_save_fm DFF_W534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1010B));
DFF_save_fm DFF_W535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1011B));
DFF_save_fm DFF_W536(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1012B));
DFF_save_fm DFF_W537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1020B));
DFF_save_fm DFF_W538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1021B));
DFF_save_fm DFF_W539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1022B));
DFF_save_fm DFF_W540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1000C));
DFF_save_fm DFF_W541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1001C));
DFF_save_fm DFF_W542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1002C));
DFF_save_fm DFF_W543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1010C));
DFF_save_fm DFF_W544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1011C));
DFF_save_fm DFF_W545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1012C));
DFF_save_fm DFF_W546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1020C));
DFF_save_fm DFF_W547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1021C));
DFF_save_fm DFF_W548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1022C));
DFF_save_fm DFF_W549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1000D));
DFF_save_fm DFF_W550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1001D));
DFF_save_fm DFF_W551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1002D));
DFF_save_fm DFF_W552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1010D));
DFF_save_fm DFF_W553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1011D));
DFF_save_fm DFF_W554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1012D));
DFF_save_fm DFF_W555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1020D));
DFF_save_fm DFF_W556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1021D));
DFF_save_fm DFF_W557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1022D));
DFF_save_fm DFF_W558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1000E));
DFF_save_fm DFF_W559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1001E));
DFF_save_fm DFF_W560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1002E));
DFF_save_fm DFF_W561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1010E));
DFF_save_fm DFF_W562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1011E));
DFF_save_fm DFF_W563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1012E));
DFF_save_fm DFF_W564(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1020E));
DFF_save_fm DFF_W565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1021E));
DFF_save_fm DFF_W566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1022E));
DFF_save_fm DFF_W567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1000F));
DFF_save_fm DFF_W568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1001F));
DFF_save_fm DFF_W569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1002F));
DFF_save_fm DFF_W570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1010F));
DFF_save_fm DFF_W571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1011F));
DFF_save_fm DFF_W572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1012F));
DFF_save_fm DFF_W573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1020F));
DFF_save_fm DFF_W574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1021F));
DFF_save_fm DFF_W575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1022F));
DFF_save_fm DFF_W576(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11000));
DFF_save_fm DFF_W577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11010));
DFF_save_fm DFF_W578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11020));
DFF_save_fm DFF_W579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11100));
DFF_save_fm DFF_W580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11110));
DFF_save_fm DFF_W581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11120));
DFF_save_fm DFF_W582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11200));
DFF_save_fm DFF_W583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11210));
DFF_save_fm DFF_W584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11220));
DFF_save_fm DFF_W585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11001));
DFF_save_fm DFF_W586(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11011));
DFF_save_fm DFF_W587(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11021));
DFF_save_fm DFF_W588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11101));
DFF_save_fm DFF_W589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11111));
DFF_save_fm DFF_W590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11121));
DFF_save_fm DFF_W591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11201));
DFF_save_fm DFF_W592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11211));
DFF_save_fm DFF_W593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11221));
DFF_save_fm DFF_W594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11002));
DFF_save_fm DFF_W595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11012));
DFF_save_fm DFF_W596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11022));
DFF_save_fm DFF_W597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11102));
DFF_save_fm DFF_W598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11112));
DFF_save_fm DFF_W599(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11122));
DFF_save_fm DFF_W600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11202));
DFF_save_fm DFF_W601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11212));
DFF_save_fm DFF_W602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11222));
DFF_save_fm DFF_W603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11003));
DFF_save_fm DFF_W604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11013));
DFF_save_fm DFF_W605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11023));
DFF_save_fm DFF_W606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11103));
DFF_save_fm DFF_W607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11113));
DFF_save_fm DFF_W608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11123));
DFF_save_fm DFF_W609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11203));
DFF_save_fm DFF_W610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11213));
DFF_save_fm DFF_W611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11223));
DFF_save_fm DFF_W612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11004));
DFF_save_fm DFF_W613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11014));
DFF_save_fm DFF_W614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11024));
DFF_save_fm DFF_W615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11104));
DFF_save_fm DFF_W616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11114));
DFF_save_fm DFF_W617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11124));
DFF_save_fm DFF_W618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11204));
DFF_save_fm DFF_W619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11214));
DFF_save_fm DFF_W620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11224));
DFF_save_fm DFF_W621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11005));
DFF_save_fm DFF_W622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11015));
DFF_save_fm DFF_W623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11025));
DFF_save_fm DFF_W624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11105));
DFF_save_fm DFF_W625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11115));
DFF_save_fm DFF_W626(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11125));
DFF_save_fm DFF_W627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11205));
DFF_save_fm DFF_W628(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11215));
DFF_save_fm DFF_W629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11225));
DFF_save_fm DFF_W630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11006));
DFF_save_fm DFF_W631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11016));
DFF_save_fm DFF_W632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11026));
DFF_save_fm DFF_W633(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11106));
DFF_save_fm DFF_W634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11116));
DFF_save_fm DFF_W635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11126));
DFF_save_fm DFF_W636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11206));
DFF_save_fm DFF_W637(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11216));
DFF_save_fm DFF_W638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11226));
DFF_save_fm DFF_W639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11007));
DFF_save_fm DFF_W640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11017));
DFF_save_fm DFF_W641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11027));
DFF_save_fm DFF_W642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11107));
DFF_save_fm DFF_W643(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11117));
DFF_save_fm DFF_W644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11127));
DFF_save_fm DFF_W645(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11207));
DFF_save_fm DFF_W646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11217));
DFF_save_fm DFF_W647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11227));
DFF_save_fm DFF_W648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11008));
DFF_save_fm DFF_W649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11018));
DFF_save_fm DFF_W650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11028));
DFF_save_fm DFF_W651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11108));
DFF_save_fm DFF_W652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11118));
DFF_save_fm DFF_W653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11128));
DFF_save_fm DFF_W654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11208));
DFF_save_fm DFF_W655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11218));
DFF_save_fm DFF_W656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11228));
DFF_save_fm DFF_W657(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11009));
DFF_save_fm DFF_W658(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11019));
DFF_save_fm DFF_W659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11029));
DFF_save_fm DFF_W660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11109));
DFF_save_fm DFF_W661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11119));
DFF_save_fm DFF_W662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11129));
DFF_save_fm DFF_W663(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11209));
DFF_save_fm DFF_W664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11219));
DFF_save_fm DFF_W665(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11229));
DFF_save_fm DFF_W666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1100A));
DFF_save_fm DFF_W667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1101A));
DFF_save_fm DFF_W668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1102A));
DFF_save_fm DFF_W669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1110A));
DFF_save_fm DFF_W670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1111A));
DFF_save_fm DFF_W671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1112A));
DFF_save_fm DFF_W672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1120A));
DFF_save_fm DFF_W673(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1121A));
DFF_save_fm DFF_W674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1122A));
DFF_save_fm DFF_W675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1100B));
DFF_save_fm DFF_W676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1101B));
DFF_save_fm DFF_W677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1102B));
DFF_save_fm DFF_W678(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1110B));
DFF_save_fm DFF_W679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1111B));
DFF_save_fm DFF_W680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1112B));
DFF_save_fm DFF_W681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1120B));
DFF_save_fm DFF_W682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1121B));
DFF_save_fm DFF_W683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1122B));
DFF_save_fm DFF_W684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1100C));
DFF_save_fm DFF_W685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1101C));
DFF_save_fm DFF_W686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1102C));
DFF_save_fm DFF_W687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1110C));
DFF_save_fm DFF_W688(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1111C));
DFF_save_fm DFF_W689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1112C));
DFF_save_fm DFF_W690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1120C));
DFF_save_fm DFF_W691(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1121C));
DFF_save_fm DFF_W692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1122C));
DFF_save_fm DFF_W693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1100D));
DFF_save_fm DFF_W694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1101D));
DFF_save_fm DFF_W695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1102D));
DFF_save_fm DFF_W696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1110D));
DFF_save_fm DFF_W697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1111D));
DFF_save_fm DFF_W698(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1112D));
DFF_save_fm DFF_W699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1120D));
DFF_save_fm DFF_W700(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1121D));
DFF_save_fm DFF_W701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1122D));
DFF_save_fm DFF_W702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1100E));
DFF_save_fm DFF_W703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1101E));
DFF_save_fm DFF_W704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1102E));
DFF_save_fm DFF_W705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1110E));
DFF_save_fm DFF_W706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1111E));
DFF_save_fm DFF_W707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1112E));
DFF_save_fm DFF_W708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1120E));
DFF_save_fm DFF_W709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1121E));
DFF_save_fm DFF_W710(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1122E));
DFF_save_fm DFF_W711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1100F));
DFF_save_fm DFF_W712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1101F));
DFF_save_fm DFF_W713(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1102F));
DFF_save_fm DFF_W714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1110F));
DFF_save_fm DFF_W715(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1111F));
DFF_save_fm DFF_W716(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1112F));
DFF_save_fm DFF_W717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1120F));
DFF_save_fm DFF_W718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1121F));
DFF_save_fm DFF_W719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1122F));
DFF_save_fm DFF_W720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12000));
DFF_save_fm DFF_W721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12010));
DFF_save_fm DFF_W722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12020));
DFF_save_fm DFF_W723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12100));
DFF_save_fm DFF_W724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12110));
DFF_save_fm DFF_W725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12120));
DFF_save_fm DFF_W726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12200));
DFF_save_fm DFF_W727(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12210));
DFF_save_fm DFF_W728(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12220));
DFF_save_fm DFF_W729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12001));
DFF_save_fm DFF_W730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12011));
DFF_save_fm DFF_W731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12021));
DFF_save_fm DFF_W732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12101));
DFF_save_fm DFF_W733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12111));
DFF_save_fm DFF_W734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12121));
DFF_save_fm DFF_W735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12201));
DFF_save_fm DFF_W736(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12211));
DFF_save_fm DFF_W737(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12221));
DFF_save_fm DFF_W738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12002));
DFF_save_fm DFF_W739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12012));
DFF_save_fm DFF_W740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12022));
DFF_save_fm DFF_W741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12102));
DFF_save_fm DFF_W742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12112));
DFF_save_fm DFF_W743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12122));
DFF_save_fm DFF_W744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12202));
DFF_save_fm DFF_W745(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12212));
DFF_save_fm DFF_W746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12222));
DFF_save_fm DFF_W747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12003));
DFF_save_fm DFF_W748(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12013));
DFF_save_fm DFF_W749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12023));
DFF_save_fm DFF_W750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12103));
DFF_save_fm DFF_W751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12113));
DFF_save_fm DFF_W752(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12123));
DFF_save_fm DFF_W753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12203));
DFF_save_fm DFF_W754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12213));
DFF_save_fm DFF_W755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12223));
DFF_save_fm DFF_W756(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12004));
DFF_save_fm DFF_W757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12014));
DFF_save_fm DFF_W758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12024));
DFF_save_fm DFF_W759(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12104));
DFF_save_fm DFF_W760(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12114));
DFF_save_fm DFF_W761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12124));
DFF_save_fm DFF_W762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12204));
DFF_save_fm DFF_W763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12214));
DFF_save_fm DFF_W764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12224));
DFF_save_fm DFF_W765(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12005));
DFF_save_fm DFF_W766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12015));
DFF_save_fm DFF_W767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12025));
DFF_save_fm DFF_W768(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12105));
DFF_save_fm DFF_W769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12115));
DFF_save_fm DFF_W770(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12125));
DFF_save_fm DFF_W771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12205));
DFF_save_fm DFF_W772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12215));
DFF_save_fm DFF_W773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12225));
DFF_save_fm DFF_W774(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12006));
DFF_save_fm DFF_W775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12016));
DFF_save_fm DFF_W776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12026));
DFF_save_fm DFF_W777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12106));
DFF_save_fm DFF_W778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12116));
DFF_save_fm DFF_W779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12126));
DFF_save_fm DFF_W780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12206));
DFF_save_fm DFF_W781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12216));
DFF_save_fm DFF_W782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12226));
DFF_save_fm DFF_W783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12007));
DFF_save_fm DFF_W784(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12017));
DFF_save_fm DFF_W785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12027));
DFF_save_fm DFF_W786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12107));
DFF_save_fm DFF_W787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12117));
DFF_save_fm DFF_W788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12127));
DFF_save_fm DFF_W789(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12207));
DFF_save_fm DFF_W790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12217));
DFF_save_fm DFF_W791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12227));
DFF_save_fm DFF_W792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12008));
DFF_save_fm DFF_W793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12018));
DFF_save_fm DFF_W794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12028));
DFF_save_fm DFF_W795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12108));
DFF_save_fm DFF_W796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12118));
DFF_save_fm DFF_W797(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12128));
DFF_save_fm DFF_W798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12208));
DFF_save_fm DFF_W799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12218));
DFF_save_fm DFF_W800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12228));
DFF_save_fm DFF_W801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12009));
DFF_save_fm DFF_W802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12019));
DFF_save_fm DFF_W803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12029));
DFF_save_fm DFF_W804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12109));
DFF_save_fm DFF_W805(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12119));
DFF_save_fm DFF_W806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12129));
DFF_save_fm DFF_W807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12209));
DFF_save_fm DFF_W808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12219));
DFF_save_fm DFF_W809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12229));
DFF_save_fm DFF_W810(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1200A));
DFF_save_fm DFF_W811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1201A));
DFF_save_fm DFF_W812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1202A));
DFF_save_fm DFF_W813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1210A));
DFF_save_fm DFF_W814(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1211A));
DFF_save_fm DFF_W815(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1212A));
DFF_save_fm DFF_W816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1220A));
DFF_save_fm DFF_W817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1221A));
DFF_save_fm DFF_W818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1222A));
DFF_save_fm DFF_W819(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1200B));
DFF_save_fm DFF_W820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1201B));
DFF_save_fm DFF_W821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1202B));
DFF_save_fm DFF_W822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1210B));
DFF_save_fm DFF_W823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1211B));
DFF_save_fm DFF_W824(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1212B));
DFF_save_fm DFF_W825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1220B));
DFF_save_fm DFF_W826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1221B));
DFF_save_fm DFF_W827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1222B));
DFF_save_fm DFF_W828(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1200C));
DFF_save_fm DFF_W829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1201C));
DFF_save_fm DFF_W830(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1202C));
DFF_save_fm DFF_W831(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1210C));
DFF_save_fm DFF_W832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1211C));
DFF_save_fm DFF_W833(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1212C));
DFF_save_fm DFF_W834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1220C));
DFF_save_fm DFF_W835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1221C));
DFF_save_fm DFF_W836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1222C));
DFF_save_fm DFF_W837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1200D));
DFF_save_fm DFF_W838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1201D));
DFF_save_fm DFF_W839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1202D));
DFF_save_fm DFF_W840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1210D));
DFF_save_fm DFF_W841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1211D));
DFF_save_fm DFF_W842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1212D));
DFF_save_fm DFF_W843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1220D));
DFF_save_fm DFF_W844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1221D));
DFF_save_fm DFF_W845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1222D));
DFF_save_fm DFF_W846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1200E));
DFF_save_fm DFF_W847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1201E));
DFF_save_fm DFF_W848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1202E));
DFF_save_fm DFF_W849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1210E));
DFF_save_fm DFF_W850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1211E));
DFF_save_fm DFF_W851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1212E));
DFF_save_fm DFF_W852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1220E));
DFF_save_fm DFF_W853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1221E));
DFF_save_fm DFF_W854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1222E));
DFF_save_fm DFF_W855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1200F));
DFF_save_fm DFF_W856(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1201F));
DFF_save_fm DFF_W857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1202F));
DFF_save_fm DFF_W858(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1210F));
DFF_save_fm DFF_W859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1211F));
DFF_save_fm DFF_W860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1212F));
DFF_save_fm DFF_W861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1220F));
DFF_save_fm DFF_W862(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1221F));
DFF_save_fm DFF_W863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1222F));
DFF_save_fm DFF_W864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13000));
DFF_save_fm DFF_W865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13010));
DFF_save_fm DFF_W866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13020));
DFF_save_fm DFF_W867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13100));
DFF_save_fm DFF_W868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13110));
DFF_save_fm DFF_W869(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13120));
DFF_save_fm DFF_W870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13200));
DFF_save_fm DFF_W871(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13210));
DFF_save_fm DFF_W872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13220));
DFF_save_fm DFF_W873(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13001));
DFF_save_fm DFF_W874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13011));
DFF_save_fm DFF_W875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13021));
DFF_save_fm DFF_W876(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13101));
DFF_save_fm DFF_W877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13111));
DFF_save_fm DFF_W878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13121));
DFF_save_fm DFF_W879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13201));
DFF_save_fm DFF_W880(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13211));
DFF_save_fm DFF_W881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13221));
DFF_save_fm DFF_W882(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13002));
DFF_save_fm DFF_W883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13012));
DFF_save_fm DFF_W884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13022));
DFF_save_fm DFF_W885(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13102));
DFF_save_fm DFF_W886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13112));
DFF_save_fm DFF_W887(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13122));
DFF_save_fm DFF_W888(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13202));
DFF_save_fm DFF_W889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13212));
DFF_save_fm DFF_W890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13222));
DFF_save_fm DFF_W891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13003));
DFF_save_fm DFF_W892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13013));
DFF_save_fm DFF_W893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13023));
DFF_save_fm DFF_W894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13103));
DFF_save_fm DFF_W895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13113));
DFF_save_fm DFF_W896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13123));
DFF_save_fm DFF_W897(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13203));
DFF_save_fm DFF_W898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13213));
DFF_save_fm DFF_W899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13223));
DFF_save_fm DFF_W900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13004));
DFF_save_fm DFF_W901(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13014));
DFF_save_fm DFF_W902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13024));
DFF_save_fm DFF_W903(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13104));
DFF_save_fm DFF_W904(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13114));
DFF_save_fm DFF_W905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13124));
DFF_save_fm DFF_W906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13204));
DFF_save_fm DFF_W907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13214));
DFF_save_fm DFF_W908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13224));
DFF_save_fm DFF_W909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13005));
DFF_save_fm DFF_W910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13015));
DFF_save_fm DFF_W911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13025));
DFF_save_fm DFF_W912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13105));
DFF_save_fm DFF_W913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13115));
DFF_save_fm DFF_W914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13125));
DFF_save_fm DFF_W915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13205));
DFF_save_fm DFF_W916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13215));
DFF_save_fm DFF_W917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13225));
DFF_save_fm DFF_W918(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13006));
DFF_save_fm DFF_W919(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13016));
DFF_save_fm DFF_W920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13026));
DFF_save_fm DFF_W921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13106));
DFF_save_fm DFF_W922(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13116));
DFF_save_fm DFF_W923(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13126));
DFF_save_fm DFF_W924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13206));
DFF_save_fm DFF_W925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13216));
DFF_save_fm DFF_W926(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13226));
DFF_save_fm DFF_W927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13007));
DFF_save_fm DFF_W928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13017));
DFF_save_fm DFF_W929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13027));
DFF_save_fm DFF_W930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13107));
DFF_save_fm DFF_W931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13117));
DFF_save_fm DFF_W932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13127));
DFF_save_fm DFF_W933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13207));
DFF_save_fm DFF_W934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13217));
DFF_save_fm DFF_W935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13227));
DFF_save_fm DFF_W936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13008));
DFF_save_fm DFF_W937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13018));
DFF_save_fm DFF_W938(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13028));
DFF_save_fm DFF_W939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13108));
DFF_save_fm DFF_W940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13118));
DFF_save_fm DFF_W941(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13128));
DFF_save_fm DFF_W942(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13208));
DFF_save_fm DFF_W943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13218));
DFF_save_fm DFF_W944(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13228));
DFF_save_fm DFF_W945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13009));
DFF_save_fm DFF_W946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13019));
DFF_save_fm DFF_W947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13029));
DFF_save_fm DFF_W948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13109));
DFF_save_fm DFF_W949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13119));
DFF_save_fm DFF_W950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13129));
DFF_save_fm DFF_W951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13209));
DFF_save_fm DFF_W952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13219));
DFF_save_fm DFF_W953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13229));
DFF_save_fm DFF_W954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1300A));
DFF_save_fm DFF_W955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1301A));
DFF_save_fm DFF_W956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1302A));
DFF_save_fm DFF_W957(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1310A));
DFF_save_fm DFF_W958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1311A));
DFF_save_fm DFF_W959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1312A));
DFF_save_fm DFF_W960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1320A));
DFF_save_fm DFF_W961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1321A));
DFF_save_fm DFF_W962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1322A));
DFF_save_fm DFF_W963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1300B));
DFF_save_fm DFF_W964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1301B));
DFF_save_fm DFF_W965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1302B));
DFF_save_fm DFF_W966(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1310B));
DFF_save_fm DFF_W967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1311B));
DFF_save_fm DFF_W968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1312B));
DFF_save_fm DFF_W969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1320B));
DFF_save_fm DFF_W970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1321B));
DFF_save_fm DFF_W971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1322B));
DFF_save_fm DFF_W972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1300C));
DFF_save_fm DFF_W973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1301C));
DFF_save_fm DFF_W974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1302C));
DFF_save_fm DFF_W975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1310C));
DFF_save_fm DFF_W976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1311C));
DFF_save_fm DFF_W977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1312C));
DFF_save_fm DFF_W978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1320C));
DFF_save_fm DFF_W979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1321C));
DFF_save_fm DFF_W980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1322C));
DFF_save_fm DFF_W981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1300D));
DFF_save_fm DFF_W982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1301D));
DFF_save_fm DFF_W983(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1302D));
DFF_save_fm DFF_W984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1310D));
DFF_save_fm DFF_W985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1311D));
DFF_save_fm DFF_W986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1312D));
DFF_save_fm DFF_W987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1320D));
DFF_save_fm DFF_W988(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1321D));
DFF_save_fm DFF_W989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1322D));
DFF_save_fm DFF_W990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1300E));
DFF_save_fm DFF_W991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1301E));
DFF_save_fm DFF_W992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1302E));
DFF_save_fm DFF_W993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1310E));
DFF_save_fm DFF_W994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1311E));
DFF_save_fm DFF_W995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1312E));
DFF_save_fm DFF_W996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1320E));
DFF_save_fm DFF_W997(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1321E));
DFF_save_fm DFF_W998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1322E));
DFF_save_fm DFF_W999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1300F));
DFF_save_fm DFF_W1000(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1301F));
DFF_save_fm DFF_W1001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1302F));
DFF_save_fm DFF_W1002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1310F));
DFF_save_fm DFF_W1003(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1311F));
DFF_save_fm DFF_W1004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1312F));
DFF_save_fm DFF_W1005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1320F));
DFF_save_fm DFF_W1006(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1321F));
DFF_save_fm DFF_W1007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1322F));
DFF_save_fm DFF_W1008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14000));
DFF_save_fm DFF_W1009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14010));
DFF_save_fm DFF_W1010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14020));
DFF_save_fm DFF_W1011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14100));
DFF_save_fm DFF_W1012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14110));
DFF_save_fm DFF_W1013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14120));
DFF_save_fm DFF_W1014(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14200));
DFF_save_fm DFF_W1015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14210));
DFF_save_fm DFF_W1016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14220));
DFF_save_fm DFF_W1017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14001));
DFF_save_fm DFF_W1018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14011));
DFF_save_fm DFF_W1019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14021));
DFF_save_fm DFF_W1020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14101));
DFF_save_fm DFF_W1021(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14111));
DFF_save_fm DFF_W1022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14121));
DFF_save_fm DFF_W1023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14201));
DFF_save_fm DFF_W1024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14211));
DFF_save_fm DFF_W1025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14221));
DFF_save_fm DFF_W1026(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14002));
DFF_save_fm DFF_W1027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14012));
DFF_save_fm DFF_W1028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14022));
DFF_save_fm DFF_W1029(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14102));
DFF_save_fm DFF_W1030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14112));
DFF_save_fm DFF_W1031(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14122));
DFF_save_fm DFF_W1032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14202));
DFF_save_fm DFF_W1033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14212));
DFF_save_fm DFF_W1034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14222));
DFF_save_fm DFF_W1035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14003));
DFF_save_fm DFF_W1036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14013));
DFF_save_fm DFF_W1037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14023));
DFF_save_fm DFF_W1038(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14103));
DFF_save_fm DFF_W1039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14113));
DFF_save_fm DFF_W1040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14123));
DFF_save_fm DFF_W1041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14203));
DFF_save_fm DFF_W1042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14213));
DFF_save_fm DFF_W1043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14223));
DFF_save_fm DFF_W1044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14004));
DFF_save_fm DFF_W1045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14014));
DFF_save_fm DFF_W1046(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14024));
DFF_save_fm DFF_W1047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14104));
DFF_save_fm DFF_W1048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14114));
DFF_save_fm DFF_W1049(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14124));
DFF_save_fm DFF_W1050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14204));
DFF_save_fm DFF_W1051(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14214));
DFF_save_fm DFF_W1052(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14224));
DFF_save_fm DFF_W1053(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14005));
DFF_save_fm DFF_W1054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14015));
DFF_save_fm DFF_W1055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14025));
DFF_save_fm DFF_W1056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14105));
DFF_save_fm DFF_W1057(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14115));
DFF_save_fm DFF_W1058(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14125));
DFF_save_fm DFF_W1059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14205));
DFF_save_fm DFF_W1060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14215));
DFF_save_fm DFF_W1061(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14225));
DFF_save_fm DFF_W1062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14006));
DFF_save_fm DFF_W1063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14016));
DFF_save_fm DFF_W1064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14026));
DFF_save_fm DFF_W1065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14106));
DFF_save_fm DFF_W1066(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14116));
DFF_save_fm DFF_W1067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14126));
DFF_save_fm DFF_W1068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14206));
DFF_save_fm DFF_W1069(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14216));
DFF_save_fm DFF_W1070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14226));
DFF_save_fm DFF_W1071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14007));
DFF_save_fm DFF_W1072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14017));
DFF_save_fm DFF_W1073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14027));
DFF_save_fm DFF_W1074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14107));
DFF_save_fm DFF_W1075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14117));
DFF_save_fm DFF_W1076(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14127));
DFF_save_fm DFF_W1077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14207));
DFF_save_fm DFF_W1078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14217));
DFF_save_fm DFF_W1079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14227));
DFF_save_fm DFF_W1080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14008));
DFF_save_fm DFF_W1081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14018));
DFF_save_fm DFF_W1082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14028));
DFF_save_fm DFF_W1083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14108));
DFF_save_fm DFF_W1084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14118));
DFF_save_fm DFF_W1085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14128));
DFF_save_fm DFF_W1086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14208));
DFF_save_fm DFF_W1087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14218));
DFF_save_fm DFF_W1088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14228));
DFF_save_fm DFF_W1089(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14009));
DFF_save_fm DFF_W1090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14019));
DFF_save_fm DFF_W1091(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14029));
DFF_save_fm DFF_W1092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14109));
DFF_save_fm DFF_W1093(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14119));
DFF_save_fm DFF_W1094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14129));
DFF_save_fm DFF_W1095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14209));
DFF_save_fm DFF_W1096(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14219));
DFF_save_fm DFF_W1097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14229));
DFF_save_fm DFF_W1098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1400A));
DFF_save_fm DFF_W1099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1401A));
DFF_save_fm DFF_W1100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1402A));
DFF_save_fm DFF_W1101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1410A));
DFF_save_fm DFF_W1102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1411A));
DFF_save_fm DFF_W1103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1412A));
DFF_save_fm DFF_W1104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1420A));
DFF_save_fm DFF_W1105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1421A));
DFF_save_fm DFF_W1106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1422A));
DFF_save_fm DFF_W1107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1400B));
DFF_save_fm DFF_W1108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1401B));
DFF_save_fm DFF_W1109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1402B));
DFF_save_fm DFF_W1110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1410B));
DFF_save_fm DFF_W1111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1411B));
DFF_save_fm DFF_W1112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1412B));
DFF_save_fm DFF_W1113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1420B));
DFF_save_fm DFF_W1114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1421B));
DFF_save_fm DFF_W1115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1422B));
DFF_save_fm DFF_W1116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1400C));
DFF_save_fm DFF_W1117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1401C));
DFF_save_fm DFF_W1118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1402C));
DFF_save_fm DFF_W1119(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1410C));
DFF_save_fm DFF_W1120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1411C));
DFF_save_fm DFF_W1121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1412C));
DFF_save_fm DFF_W1122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1420C));
DFF_save_fm DFF_W1123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1421C));
DFF_save_fm DFF_W1124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1422C));
DFF_save_fm DFF_W1125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1400D));
DFF_save_fm DFF_W1126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1401D));
DFF_save_fm DFF_W1127(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1402D));
DFF_save_fm DFF_W1128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1410D));
DFF_save_fm DFF_W1129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1411D));
DFF_save_fm DFF_W1130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1412D));
DFF_save_fm DFF_W1131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1420D));
DFF_save_fm DFF_W1132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1421D));
DFF_save_fm DFF_W1133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1422D));
DFF_save_fm DFF_W1134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1400E));
DFF_save_fm DFF_W1135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1401E));
DFF_save_fm DFF_W1136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1402E));
DFF_save_fm DFF_W1137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1410E));
DFF_save_fm DFF_W1138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1411E));
DFF_save_fm DFF_W1139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1412E));
DFF_save_fm DFF_W1140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1420E));
DFF_save_fm DFF_W1141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1421E));
DFF_save_fm DFF_W1142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1422E));
DFF_save_fm DFF_W1143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1400F));
DFF_save_fm DFF_W1144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1401F));
DFF_save_fm DFF_W1145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1402F));
DFF_save_fm DFF_W1146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1410F));
DFF_save_fm DFF_W1147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1411F));
DFF_save_fm DFF_W1148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1412F));
DFF_save_fm DFF_W1149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1420F));
DFF_save_fm DFF_W1150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1421F));
DFF_save_fm DFF_W1151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1422F));
DFF_save_fm DFF_W1152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15000));
DFF_save_fm DFF_W1153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15010));
DFF_save_fm DFF_W1154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15020));
DFF_save_fm DFF_W1155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15100));
DFF_save_fm DFF_W1156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15110));
DFF_save_fm DFF_W1157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15120));
DFF_save_fm DFF_W1158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15200));
DFF_save_fm DFF_W1159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15210));
DFF_save_fm DFF_W1160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15220));
DFF_save_fm DFF_W1161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15001));
DFF_save_fm DFF_W1162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15011));
DFF_save_fm DFF_W1163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15021));
DFF_save_fm DFF_W1164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15101));
DFF_save_fm DFF_W1165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15111));
DFF_save_fm DFF_W1166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15121));
DFF_save_fm DFF_W1167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15201));
DFF_save_fm DFF_W1168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15211));
DFF_save_fm DFF_W1169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15221));
DFF_save_fm DFF_W1170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15002));
DFF_save_fm DFF_W1171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15012));
DFF_save_fm DFF_W1172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15022));
DFF_save_fm DFF_W1173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15102));
DFF_save_fm DFF_W1174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15112));
DFF_save_fm DFF_W1175(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15122));
DFF_save_fm DFF_W1176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15202));
DFF_save_fm DFF_W1177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15212));
DFF_save_fm DFF_W1178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15222));
DFF_save_fm DFF_W1179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15003));
DFF_save_fm DFF_W1180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15013));
DFF_save_fm DFF_W1181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15023));
DFF_save_fm DFF_W1182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15103));
DFF_save_fm DFF_W1183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15113));
DFF_save_fm DFF_W1184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15123));
DFF_save_fm DFF_W1185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15203));
DFF_save_fm DFF_W1186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15213));
DFF_save_fm DFF_W1187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15223));
DFF_save_fm DFF_W1188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15004));
DFF_save_fm DFF_W1189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15014));
DFF_save_fm DFF_W1190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15024));
DFF_save_fm DFF_W1191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15104));
DFF_save_fm DFF_W1192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15114));
DFF_save_fm DFF_W1193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15124));
DFF_save_fm DFF_W1194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15204));
DFF_save_fm DFF_W1195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15214));
DFF_save_fm DFF_W1196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15224));
DFF_save_fm DFF_W1197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15005));
DFF_save_fm DFF_W1198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15015));
DFF_save_fm DFF_W1199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15025));
DFF_save_fm DFF_W1200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15105));
DFF_save_fm DFF_W1201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15115));
DFF_save_fm DFF_W1202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15125));
DFF_save_fm DFF_W1203(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15205));
DFF_save_fm DFF_W1204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15215));
DFF_save_fm DFF_W1205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15225));
DFF_save_fm DFF_W1206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15006));
DFF_save_fm DFF_W1207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15016));
DFF_save_fm DFF_W1208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15026));
DFF_save_fm DFF_W1209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15106));
DFF_save_fm DFF_W1210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15116));
DFF_save_fm DFF_W1211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15126));
DFF_save_fm DFF_W1212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15206));
DFF_save_fm DFF_W1213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15216));
DFF_save_fm DFF_W1214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15226));
DFF_save_fm DFF_W1215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15007));
DFF_save_fm DFF_W1216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15017));
DFF_save_fm DFF_W1217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15027));
DFF_save_fm DFF_W1218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15107));
DFF_save_fm DFF_W1219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15117));
DFF_save_fm DFF_W1220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15127));
DFF_save_fm DFF_W1221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15207));
DFF_save_fm DFF_W1222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15217));
DFF_save_fm DFF_W1223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15227));
DFF_save_fm DFF_W1224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15008));
DFF_save_fm DFF_W1225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15018));
DFF_save_fm DFF_W1226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15028));
DFF_save_fm DFF_W1227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15108));
DFF_save_fm DFF_W1228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15118));
DFF_save_fm DFF_W1229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15128));
DFF_save_fm DFF_W1230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15208));
DFF_save_fm DFF_W1231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15218));
DFF_save_fm DFF_W1232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15228));
DFF_save_fm DFF_W1233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15009));
DFF_save_fm DFF_W1234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15019));
DFF_save_fm DFF_W1235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15029));
DFF_save_fm DFF_W1236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15109));
DFF_save_fm DFF_W1237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15119));
DFF_save_fm DFF_W1238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15129));
DFF_save_fm DFF_W1239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15209));
DFF_save_fm DFF_W1240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15219));
DFF_save_fm DFF_W1241(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15229));
DFF_save_fm DFF_W1242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1500A));
DFF_save_fm DFF_W1243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1501A));
DFF_save_fm DFF_W1244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1502A));
DFF_save_fm DFF_W1245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1510A));
DFF_save_fm DFF_W1246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1511A));
DFF_save_fm DFF_W1247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1512A));
DFF_save_fm DFF_W1248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1520A));
DFF_save_fm DFF_W1249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1521A));
DFF_save_fm DFF_W1250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1522A));
DFF_save_fm DFF_W1251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1500B));
DFF_save_fm DFF_W1252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1501B));
DFF_save_fm DFF_W1253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1502B));
DFF_save_fm DFF_W1254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1510B));
DFF_save_fm DFF_W1255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1511B));
DFF_save_fm DFF_W1256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1512B));
DFF_save_fm DFF_W1257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1520B));
DFF_save_fm DFF_W1258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1521B));
DFF_save_fm DFF_W1259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1522B));
DFF_save_fm DFF_W1260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1500C));
DFF_save_fm DFF_W1261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1501C));
DFF_save_fm DFF_W1262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1502C));
DFF_save_fm DFF_W1263(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1510C));
DFF_save_fm DFF_W1264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1511C));
DFF_save_fm DFF_W1265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1512C));
DFF_save_fm DFF_W1266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1520C));
DFF_save_fm DFF_W1267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1521C));
DFF_save_fm DFF_W1268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1522C));
DFF_save_fm DFF_W1269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1500D));
DFF_save_fm DFF_W1270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1501D));
DFF_save_fm DFF_W1271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1502D));
DFF_save_fm DFF_W1272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1510D));
DFF_save_fm DFF_W1273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1511D));
DFF_save_fm DFF_W1274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1512D));
DFF_save_fm DFF_W1275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1520D));
DFF_save_fm DFF_W1276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1521D));
DFF_save_fm DFF_W1277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1522D));
DFF_save_fm DFF_W1278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1500E));
DFF_save_fm DFF_W1279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1501E));
DFF_save_fm DFF_W1280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1502E));
DFF_save_fm DFF_W1281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1510E));
DFF_save_fm DFF_W1282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1511E));
DFF_save_fm DFF_W1283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1512E));
DFF_save_fm DFF_W1284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1520E));
DFF_save_fm DFF_W1285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1521E));
DFF_save_fm DFF_W1286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1522E));
DFF_save_fm DFF_W1287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1500F));
DFF_save_fm DFF_W1288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1501F));
DFF_save_fm DFF_W1289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1502F));
DFF_save_fm DFF_W1290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1510F));
DFF_save_fm DFF_W1291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1511F));
DFF_save_fm DFF_W1292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1512F));
DFF_save_fm DFF_W1293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1520F));
DFF_save_fm DFF_W1294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1521F));
DFF_save_fm DFF_W1295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1522F));
DFF_save_fm DFF_W1296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16000));
DFF_save_fm DFF_W1297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16010));
DFF_save_fm DFF_W1298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16020));
DFF_save_fm DFF_W1299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16100));
DFF_save_fm DFF_W1300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16110));
DFF_save_fm DFF_W1301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16120));
DFF_save_fm DFF_W1302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16200));
DFF_save_fm DFF_W1303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16210));
DFF_save_fm DFF_W1304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16220));
DFF_save_fm DFF_W1305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16001));
DFF_save_fm DFF_W1306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16011));
DFF_save_fm DFF_W1307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16021));
DFF_save_fm DFF_W1308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16101));
DFF_save_fm DFF_W1309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16111));
DFF_save_fm DFF_W1310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16121));
DFF_save_fm DFF_W1311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16201));
DFF_save_fm DFF_W1312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16211));
DFF_save_fm DFF_W1313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16221));
DFF_save_fm DFF_W1314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16002));
DFF_save_fm DFF_W1315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16012));
DFF_save_fm DFF_W1316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16022));
DFF_save_fm DFF_W1317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16102));
DFF_save_fm DFF_W1318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16112));
DFF_save_fm DFF_W1319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16122));
DFF_save_fm DFF_W1320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16202));
DFF_save_fm DFF_W1321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16212));
DFF_save_fm DFF_W1322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16222));
DFF_save_fm DFF_W1323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16003));
DFF_save_fm DFF_W1324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16013));
DFF_save_fm DFF_W1325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16023));
DFF_save_fm DFF_W1326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16103));
DFF_save_fm DFF_W1327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16113));
DFF_save_fm DFF_W1328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16123));
DFF_save_fm DFF_W1329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16203));
DFF_save_fm DFF_W1330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16213));
DFF_save_fm DFF_W1331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16223));
DFF_save_fm DFF_W1332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16004));
DFF_save_fm DFF_W1333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16014));
DFF_save_fm DFF_W1334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16024));
DFF_save_fm DFF_W1335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16104));
DFF_save_fm DFF_W1336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16114));
DFF_save_fm DFF_W1337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16124));
DFF_save_fm DFF_W1338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16204));
DFF_save_fm DFF_W1339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16214));
DFF_save_fm DFF_W1340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16224));
DFF_save_fm DFF_W1341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16005));
DFF_save_fm DFF_W1342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16015));
DFF_save_fm DFF_W1343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16025));
DFF_save_fm DFF_W1344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16105));
DFF_save_fm DFF_W1345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16115));
DFF_save_fm DFF_W1346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16125));
DFF_save_fm DFF_W1347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16205));
DFF_save_fm DFF_W1348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16215));
DFF_save_fm DFF_W1349(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16225));
DFF_save_fm DFF_W1350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16006));
DFF_save_fm DFF_W1351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16016));
DFF_save_fm DFF_W1352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16026));
DFF_save_fm DFF_W1353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16106));
DFF_save_fm DFF_W1354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16116));
DFF_save_fm DFF_W1355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16126));
DFF_save_fm DFF_W1356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16206));
DFF_save_fm DFF_W1357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16216));
DFF_save_fm DFF_W1358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16226));
DFF_save_fm DFF_W1359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16007));
DFF_save_fm DFF_W1360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16017));
DFF_save_fm DFF_W1361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16027));
DFF_save_fm DFF_W1362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16107));
DFF_save_fm DFF_W1363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16117));
DFF_save_fm DFF_W1364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16127));
DFF_save_fm DFF_W1365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16207));
DFF_save_fm DFF_W1366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16217));
DFF_save_fm DFF_W1367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16227));
DFF_save_fm DFF_W1368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16008));
DFF_save_fm DFF_W1369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16018));
DFF_save_fm DFF_W1370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16028));
DFF_save_fm DFF_W1371(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16108));
DFF_save_fm DFF_W1372(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16118));
DFF_save_fm DFF_W1373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16128));
DFF_save_fm DFF_W1374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16208));
DFF_save_fm DFF_W1375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16218));
DFF_save_fm DFF_W1376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16228));
DFF_save_fm DFF_W1377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16009));
DFF_save_fm DFF_W1378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16019));
DFF_save_fm DFF_W1379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16029));
DFF_save_fm DFF_W1380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16109));
DFF_save_fm DFF_W1381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16119));
DFF_save_fm DFF_W1382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16129));
DFF_save_fm DFF_W1383(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16209));
DFF_save_fm DFF_W1384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16219));
DFF_save_fm DFF_W1385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16229));
DFF_save_fm DFF_W1386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1600A));
DFF_save_fm DFF_W1387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1601A));
DFF_save_fm DFF_W1388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1602A));
DFF_save_fm DFF_W1389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1610A));
DFF_save_fm DFF_W1390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1611A));
DFF_save_fm DFF_W1391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1612A));
DFF_save_fm DFF_W1392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1620A));
DFF_save_fm DFF_W1393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1621A));
DFF_save_fm DFF_W1394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1622A));
DFF_save_fm DFF_W1395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1600B));
DFF_save_fm DFF_W1396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1601B));
DFF_save_fm DFF_W1397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1602B));
DFF_save_fm DFF_W1398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1610B));
DFF_save_fm DFF_W1399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1611B));
DFF_save_fm DFF_W1400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1612B));
DFF_save_fm DFF_W1401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1620B));
DFF_save_fm DFF_W1402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1621B));
DFF_save_fm DFF_W1403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1622B));
DFF_save_fm DFF_W1404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1600C));
DFF_save_fm DFF_W1405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1601C));
DFF_save_fm DFF_W1406(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1602C));
DFF_save_fm DFF_W1407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1610C));
DFF_save_fm DFF_W1408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1611C));
DFF_save_fm DFF_W1409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1612C));
DFF_save_fm DFF_W1410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1620C));
DFF_save_fm DFF_W1411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1621C));
DFF_save_fm DFF_W1412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1622C));
DFF_save_fm DFF_W1413(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1600D));
DFF_save_fm DFF_W1414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1601D));
DFF_save_fm DFF_W1415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1602D));
DFF_save_fm DFF_W1416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1610D));
DFF_save_fm DFF_W1417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1611D));
DFF_save_fm DFF_W1418(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1612D));
DFF_save_fm DFF_W1419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1620D));
DFF_save_fm DFF_W1420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1621D));
DFF_save_fm DFF_W1421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1622D));
DFF_save_fm DFF_W1422(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1600E));
DFF_save_fm DFF_W1423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1601E));
DFF_save_fm DFF_W1424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1602E));
DFF_save_fm DFF_W1425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1610E));
DFF_save_fm DFF_W1426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1611E));
DFF_save_fm DFF_W1427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1612E));
DFF_save_fm DFF_W1428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1620E));
DFF_save_fm DFF_W1429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1621E));
DFF_save_fm DFF_W1430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1622E));
DFF_save_fm DFF_W1431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1600F));
DFF_save_fm DFF_W1432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1601F));
DFF_save_fm DFF_W1433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1602F));
DFF_save_fm DFF_W1434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1610F));
DFF_save_fm DFF_W1435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1611F));
DFF_save_fm DFF_W1436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1612F));
DFF_save_fm DFF_W1437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1620F));
DFF_save_fm DFF_W1438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1621F));
DFF_save_fm DFF_W1439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1622F));
DFF_save_fm DFF_W1440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17000));
DFF_save_fm DFF_W1441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17010));
DFF_save_fm DFF_W1442(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17020));
DFF_save_fm DFF_W1443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17100));
DFF_save_fm DFF_W1444(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17110));
DFF_save_fm DFF_W1445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17120));
DFF_save_fm DFF_W1446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17200));
DFF_save_fm DFF_W1447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17210));
DFF_save_fm DFF_W1448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17220));
DFF_save_fm DFF_W1449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17001));
DFF_save_fm DFF_W1450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17011));
DFF_save_fm DFF_W1451(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17021));
DFF_save_fm DFF_W1452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17101));
DFF_save_fm DFF_W1453(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17111));
DFF_save_fm DFF_W1454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17121));
DFF_save_fm DFF_W1455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17201));
DFF_save_fm DFF_W1456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17211));
DFF_save_fm DFF_W1457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17221));
DFF_save_fm DFF_W1458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17002));
DFF_save_fm DFF_W1459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17012));
DFF_save_fm DFF_W1460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17022));
DFF_save_fm DFF_W1461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17102));
DFF_save_fm DFF_W1462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17112));
DFF_save_fm DFF_W1463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17122));
DFF_save_fm DFF_W1464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17202));
DFF_save_fm DFF_W1465(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17212));
DFF_save_fm DFF_W1466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17222));
DFF_save_fm DFF_W1467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17003));
DFF_save_fm DFF_W1468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17013));
DFF_save_fm DFF_W1469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17023));
DFF_save_fm DFF_W1470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17103));
DFF_save_fm DFF_W1471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17113));
DFF_save_fm DFF_W1472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17123));
DFF_save_fm DFF_W1473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17203));
DFF_save_fm DFF_W1474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17213));
DFF_save_fm DFF_W1475(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17223));
DFF_save_fm DFF_W1476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17004));
DFF_save_fm DFF_W1477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17014));
DFF_save_fm DFF_W1478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17024));
DFF_save_fm DFF_W1479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17104));
DFF_save_fm DFF_W1480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17114));
DFF_save_fm DFF_W1481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17124));
DFF_save_fm DFF_W1482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17204));
DFF_save_fm DFF_W1483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17214));
DFF_save_fm DFF_W1484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17224));
DFF_save_fm DFF_W1485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17005));
DFF_save_fm DFF_W1486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17015));
DFF_save_fm DFF_W1487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17025));
DFF_save_fm DFF_W1488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17105));
DFF_save_fm DFF_W1489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17115));
DFF_save_fm DFF_W1490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17125));
DFF_save_fm DFF_W1491(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17205));
DFF_save_fm DFF_W1492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17215));
DFF_save_fm DFF_W1493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17225));
DFF_save_fm DFF_W1494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17006));
DFF_save_fm DFF_W1495(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17016));
DFF_save_fm DFF_W1496(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17026));
DFF_save_fm DFF_W1497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17106));
DFF_save_fm DFF_W1498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17116));
DFF_save_fm DFF_W1499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17126));
DFF_save_fm DFF_W1500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17206));
DFF_save_fm DFF_W1501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17216));
DFF_save_fm DFF_W1502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17226));
DFF_save_fm DFF_W1503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17007));
DFF_save_fm DFF_W1504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17017));
DFF_save_fm DFF_W1505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17027));
DFF_save_fm DFF_W1506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17107));
DFF_save_fm DFF_W1507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17117));
DFF_save_fm DFF_W1508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17127));
DFF_save_fm DFF_W1509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17207));
DFF_save_fm DFF_W1510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17217));
DFF_save_fm DFF_W1511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17227));
DFF_save_fm DFF_W1512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17008));
DFF_save_fm DFF_W1513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17018));
DFF_save_fm DFF_W1514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17028));
DFF_save_fm DFF_W1515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17108));
DFF_save_fm DFF_W1516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17118));
DFF_save_fm DFF_W1517(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17128));
DFF_save_fm DFF_W1518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17208));
DFF_save_fm DFF_W1519(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17218));
DFF_save_fm DFF_W1520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17228));
DFF_save_fm DFF_W1521(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17009));
DFF_save_fm DFF_W1522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17019));
DFF_save_fm DFF_W1523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17029));
DFF_save_fm DFF_W1524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17109));
DFF_save_fm DFF_W1525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17119));
DFF_save_fm DFF_W1526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17129));
DFF_save_fm DFF_W1527(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17209));
DFF_save_fm DFF_W1528(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17219));
DFF_save_fm DFF_W1529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17229));
DFF_save_fm DFF_W1530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1700A));
DFF_save_fm DFF_W1531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1701A));
DFF_save_fm DFF_W1532(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1702A));
DFF_save_fm DFF_W1533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1710A));
DFF_save_fm DFF_W1534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1711A));
DFF_save_fm DFF_W1535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1712A));
DFF_save_fm DFF_W1536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1720A));
DFF_save_fm DFF_W1537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1721A));
DFF_save_fm DFF_W1538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1722A));
DFF_save_fm DFF_W1539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1700B));
DFF_save_fm DFF_W1540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1701B));
DFF_save_fm DFF_W1541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1702B));
DFF_save_fm DFF_W1542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1710B));
DFF_save_fm DFF_W1543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1711B));
DFF_save_fm DFF_W1544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1712B));
DFF_save_fm DFF_W1545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1720B));
DFF_save_fm DFF_W1546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1721B));
DFF_save_fm DFF_W1547(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1722B));
DFF_save_fm DFF_W1548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1700C));
DFF_save_fm DFF_W1549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1701C));
DFF_save_fm DFF_W1550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1702C));
DFF_save_fm DFF_W1551(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1710C));
DFF_save_fm DFF_W1552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1711C));
DFF_save_fm DFF_W1553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1712C));
DFF_save_fm DFF_W1554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1720C));
DFF_save_fm DFF_W1555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1721C));
DFF_save_fm DFF_W1556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1722C));
DFF_save_fm DFF_W1557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1700D));
DFF_save_fm DFF_W1558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1701D));
DFF_save_fm DFF_W1559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1702D));
DFF_save_fm DFF_W1560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1710D));
DFF_save_fm DFF_W1561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1711D));
DFF_save_fm DFF_W1562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1712D));
DFF_save_fm DFF_W1563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1720D));
DFF_save_fm DFF_W1564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1721D));
DFF_save_fm DFF_W1565(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1722D));
DFF_save_fm DFF_W1566(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1700E));
DFF_save_fm DFF_W1567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1701E));
DFF_save_fm DFF_W1568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1702E));
DFF_save_fm DFF_W1569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1710E));
DFF_save_fm DFF_W1570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1711E));
DFF_save_fm DFF_W1571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1712E));
DFF_save_fm DFF_W1572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1720E));
DFF_save_fm DFF_W1573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1721E));
DFF_save_fm DFF_W1574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1722E));
DFF_save_fm DFF_W1575(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1700F));
DFF_save_fm DFF_W1576(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1701F));
DFF_save_fm DFF_W1577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1702F));
DFF_save_fm DFF_W1578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1710F));
DFF_save_fm DFF_W1579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1711F));
DFF_save_fm DFF_W1580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1712F));
DFF_save_fm DFF_W1581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1720F));
DFF_save_fm DFF_W1582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1721F));
DFF_save_fm DFF_W1583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1722F));
DFF_save_fm DFF_W1584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18000));
DFF_save_fm DFF_W1585(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18010));
DFF_save_fm DFF_W1586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18020));
DFF_save_fm DFF_W1587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18100));
DFF_save_fm DFF_W1588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18110));
DFF_save_fm DFF_W1589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18120));
DFF_save_fm DFF_W1590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18200));
DFF_save_fm DFF_W1591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18210));
DFF_save_fm DFF_W1592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18220));
DFF_save_fm DFF_W1593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18001));
DFF_save_fm DFF_W1594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18011));
DFF_save_fm DFF_W1595(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18021));
DFF_save_fm DFF_W1596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18101));
DFF_save_fm DFF_W1597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18111));
DFF_save_fm DFF_W1598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18121));
DFF_save_fm DFF_W1599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18201));
DFF_save_fm DFF_W1600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18211));
DFF_save_fm DFF_W1601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18221));
DFF_save_fm DFF_W1602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18002));
DFF_save_fm DFF_W1603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18012));
DFF_save_fm DFF_W1604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18022));
DFF_save_fm DFF_W1605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18102));
DFF_save_fm DFF_W1606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18112));
DFF_save_fm DFF_W1607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18122));
DFF_save_fm DFF_W1608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18202));
DFF_save_fm DFF_W1609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18212));
DFF_save_fm DFF_W1610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18222));
DFF_save_fm DFF_W1611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18003));
DFF_save_fm DFF_W1612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18013));
DFF_save_fm DFF_W1613(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18023));
DFF_save_fm DFF_W1614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18103));
DFF_save_fm DFF_W1615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18113));
DFF_save_fm DFF_W1616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18123));
DFF_save_fm DFF_W1617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18203));
DFF_save_fm DFF_W1618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18213));
DFF_save_fm DFF_W1619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18223));
DFF_save_fm DFF_W1620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18004));
DFF_save_fm DFF_W1621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18014));
DFF_save_fm DFF_W1622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18024));
DFF_save_fm DFF_W1623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18104));
DFF_save_fm DFF_W1624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18114));
DFF_save_fm DFF_W1625(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18124));
DFF_save_fm DFF_W1626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18204));
DFF_save_fm DFF_W1627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18214));
DFF_save_fm DFF_W1628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18224));
DFF_save_fm DFF_W1629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18005));
DFF_save_fm DFF_W1630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18015));
DFF_save_fm DFF_W1631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18025));
DFF_save_fm DFF_W1632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18105));
DFF_save_fm DFF_W1633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18115));
DFF_save_fm DFF_W1634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18125));
DFF_save_fm DFF_W1635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18205));
DFF_save_fm DFF_W1636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18215));
DFF_save_fm DFF_W1637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18225));
DFF_save_fm DFF_W1638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18006));
DFF_save_fm DFF_W1639(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18016));
DFF_save_fm DFF_W1640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18026));
DFF_save_fm DFF_W1641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18106));
DFF_save_fm DFF_W1642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18116));
DFF_save_fm DFF_W1643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18126));
DFF_save_fm DFF_W1644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18206));
DFF_save_fm DFF_W1645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18216));
DFF_save_fm DFF_W1646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18226));
DFF_save_fm DFF_W1647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18007));
DFF_save_fm DFF_W1648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18017));
DFF_save_fm DFF_W1649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18027));
DFF_save_fm DFF_W1650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18107));
DFF_save_fm DFF_W1651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18117));
DFF_save_fm DFF_W1652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18127));
DFF_save_fm DFF_W1653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18207));
DFF_save_fm DFF_W1654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18217));
DFF_save_fm DFF_W1655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18227));
DFF_save_fm DFF_W1656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18008));
DFF_save_fm DFF_W1657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18018));
DFF_save_fm DFF_W1658(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18028));
DFF_save_fm DFF_W1659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18108));
DFF_save_fm DFF_W1660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18118));
DFF_save_fm DFF_W1661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18128));
DFF_save_fm DFF_W1662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18208));
DFF_save_fm DFF_W1663(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18218));
DFF_save_fm DFF_W1664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18228));
DFF_save_fm DFF_W1665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18009));
DFF_save_fm DFF_W1666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18019));
DFF_save_fm DFF_W1667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18029));
DFF_save_fm DFF_W1668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18109));
DFF_save_fm DFF_W1669(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18119));
DFF_save_fm DFF_W1670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18129));
DFF_save_fm DFF_W1671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18209));
DFF_save_fm DFF_W1672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18219));
DFF_save_fm DFF_W1673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18229));
DFF_save_fm DFF_W1674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1800A));
DFF_save_fm DFF_W1675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1801A));
DFF_save_fm DFF_W1676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1802A));
DFF_save_fm DFF_W1677(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1810A));
DFF_save_fm DFF_W1678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1811A));
DFF_save_fm DFF_W1679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1812A));
DFF_save_fm DFF_W1680(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1820A));
DFF_save_fm DFF_W1681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1821A));
DFF_save_fm DFF_W1682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1822A));
DFF_save_fm DFF_W1683(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1800B));
DFF_save_fm DFF_W1684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1801B));
DFF_save_fm DFF_W1685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1802B));
DFF_save_fm DFF_W1686(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1810B));
DFF_save_fm DFF_W1687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1811B));
DFF_save_fm DFF_W1688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1812B));
DFF_save_fm DFF_W1689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1820B));
DFF_save_fm DFF_W1690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1821B));
DFF_save_fm DFF_W1691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1822B));
DFF_save_fm DFF_W1692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1800C));
DFF_save_fm DFF_W1693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1801C));
DFF_save_fm DFF_W1694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1802C));
DFF_save_fm DFF_W1695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1810C));
DFF_save_fm DFF_W1696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1811C));
DFF_save_fm DFF_W1697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1812C));
DFF_save_fm DFF_W1698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1820C));
DFF_save_fm DFF_W1699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1821C));
DFF_save_fm DFF_W1700(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1822C));
DFF_save_fm DFF_W1701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1800D));
DFF_save_fm DFF_W1702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1801D));
DFF_save_fm DFF_W1703(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1802D));
DFF_save_fm DFF_W1704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1810D));
DFF_save_fm DFF_W1705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1811D));
DFF_save_fm DFF_W1706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1812D));
DFF_save_fm DFF_W1707(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1820D));
DFF_save_fm DFF_W1708(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1821D));
DFF_save_fm DFF_W1709(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1822D));
DFF_save_fm DFF_W1710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1800E));
DFF_save_fm DFF_W1711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1801E));
DFF_save_fm DFF_W1712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1802E));
DFF_save_fm DFF_W1713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1810E));
DFF_save_fm DFF_W1714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1811E));
DFF_save_fm DFF_W1715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1812E));
DFF_save_fm DFF_W1716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1820E));
DFF_save_fm DFF_W1717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1821E));
DFF_save_fm DFF_W1718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1822E));
DFF_save_fm DFF_W1719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1800F));
DFF_save_fm DFF_W1720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1801F));
DFF_save_fm DFF_W1721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1802F));
DFF_save_fm DFF_W1722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1810F));
DFF_save_fm DFF_W1723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1811F));
DFF_save_fm DFF_W1724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1812F));
DFF_save_fm DFF_W1725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1820F));
DFF_save_fm DFF_W1726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1821F));
DFF_save_fm DFF_W1727(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1822F));
DFF_save_fm DFF_W1728(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19000));
DFF_save_fm DFF_W1729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19010));
DFF_save_fm DFF_W1730(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19020));
DFF_save_fm DFF_W1731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19100));
DFF_save_fm DFF_W1732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19110));
DFF_save_fm DFF_W1733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19120));
DFF_save_fm DFF_W1734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19200));
DFF_save_fm DFF_W1735(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19210));
DFF_save_fm DFF_W1736(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19220));
DFF_save_fm DFF_W1737(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19001));
DFF_save_fm DFF_W1738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19011));
DFF_save_fm DFF_W1739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19021));
DFF_save_fm DFF_W1740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19101));
DFF_save_fm DFF_W1741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19111));
DFF_save_fm DFF_W1742(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19121));
DFF_save_fm DFF_W1743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19201));
DFF_save_fm DFF_W1744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19211));
DFF_save_fm DFF_W1745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19221));
DFF_save_fm DFF_W1746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19002));
DFF_save_fm DFF_W1747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19012));
DFF_save_fm DFF_W1748(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19022));
DFF_save_fm DFF_W1749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19102));
DFF_save_fm DFF_W1750(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19112));
DFF_save_fm DFF_W1751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19122));
DFF_save_fm DFF_W1752(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19202));
DFF_save_fm DFF_W1753(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19212));
DFF_save_fm DFF_W1754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19222));
DFF_save_fm DFF_W1755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19003));
DFF_save_fm DFF_W1756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19013));
DFF_save_fm DFF_W1757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19023));
DFF_save_fm DFF_W1758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19103));
DFF_save_fm DFF_W1759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19113));
DFF_save_fm DFF_W1760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19123));
DFF_save_fm DFF_W1761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19203));
DFF_save_fm DFF_W1762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19213));
DFF_save_fm DFF_W1763(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19223));
DFF_save_fm DFF_W1764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19004));
DFF_save_fm DFF_W1765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19014));
DFF_save_fm DFF_W1766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19024));
DFF_save_fm DFF_W1767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19104));
DFF_save_fm DFF_W1768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19114));
DFF_save_fm DFF_W1769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19124));
DFF_save_fm DFF_W1770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19204));
DFF_save_fm DFF_W1771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19214));
DFF_save_fm DFF_W1772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19224));
DFF_save_fm DFF_W1773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19005));
DFF_save_fm DFF_W1774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19015));
DFF_save_fm DFF_W1775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19025));
DFF_save_fm DFF_W1776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19105));
DFF_save_fm DFF_W1777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19115));
DFF_save_fm DFF_W1778(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19125));
DFF_save_fm DFF_W1779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19205));
DFF_save_fm DFF_W1780(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19215));
DFF_save_fm DFF_W1781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19225));
DFF_save_fm DFF_W1782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19006));
DFF_save_fm DFF_W1783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19016));
DFF_save_fm DFF_W1784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19026));
DFF_save_fm DFF_W1785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19106));
DFF_save_fm DFF_W1786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19116));
DFF_save_fm DFF_W1787(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19126));
DFF_save_fm DFF_W1788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19206));
DFF_save_fm DFF_W1789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19216));
DFF_save_fm DFF_W1790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19226));
DFF_save_fm DFF_W1791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19007));
DFF_save_fm DFF_W1792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19017));
DFF_save_fm DFF_W1793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19027));
DFF_save_fm DFF_W1794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19107));
DFF_save_fm DFF_W1795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19117));
DFF_save_fm DFF_W1796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19127));
DFF_save_fm DFF_W1797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19207));
DFF_save_fm DFF_W1798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19217));
DFF_save_fm DFF_W1799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19227));
DFF_save_fm DFF_W1800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19008));
DFF_save_fm DFF_W1801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19018));
DFF_save_fm DFF_W1802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19028));
DFF_save_fm DFF_W1803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19108));
DFF_save_fm DFF_W1804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19118));
DFF_save_fm DFF_W1805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19128));
DFF_save_fm DFF_W1806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19208));
DFF_save_fm DFF_W1807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19218));
DFF_save_fm DFF_W1808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19228));
DFF_save_fm DFF_W1809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19009));
DFF_save_fm DFF_W1810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19019));
DFF_save_fm DFF_W1811(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19029));
DFF_save_fm DFF_W1812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19109));
DFF_save_fm DFF_W1813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19119));
DFF_save_fm DFF_W1814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19129));
DFF_save_fm DFF_W1815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19209));
DFF_save_fm DFF_W1816(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19219));
DFF_save_fm DFF_W1817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19229));
DFF_save_fm DFF_W1818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1900A));
DFF_save_fm DFF_W1819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1901A));
DFF_save_fm DFF_W1820(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1902A));
DFF_save_fm DFF_W1821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1910A));
DFF_save_fm DFF_W1822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1911A));
DFF_save_fm DFF_W1823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1912A));
DFF_save_fm DFF_W1824(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1920A));
DFF_save_fm DFF_W1825(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1921A));
DFF_save_fm DFF_W1826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1922A));
DFF_save_fm DFF_W1827(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1900B));
DFF_save_fm DFF_W1828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1901B));
DFF_save_fm DFF_W1829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1902B));
DFF_save_fm DFF_W1830(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1910B));
DFF_save_fm DFF_W1831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1911B));
DFF_save_fm DFF_W1832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1912B));
DFF_save_fm DFF_W1833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1920B));
DFF_save_fm DFF_W1834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1921B));
DFF_save_fm DFF_W1835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1922B));
DFF_save_fm DFF_W1836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1900C));
DFF_save_fm DFF_W1837(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1901C));
DFF_save_fm DFF_W1838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1902C));
DFF_save_fm DFF_W1839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1910C));
DFF_save_fm DFF_W1840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1911C));
DFF_save_fm DFF_W1841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1912C));
DFF_save_fm DFF_W1842(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1920C));
DFF_save_fm DFF_W1843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1921C));
DFF_save_fm DFF_W1844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1922C));
DFF_save_fm DFF_W1845(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1900D));
DFF_save_fm DFF_W1846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1901D));
DFF_save_fm DFF_W1847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1902D));
DFF_save_fm DFF_W1848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1910D));
DFF_save_fm DFF_W1849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1911D));
DFF_save_fm DFF_W1850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1912D));
DFF_save_fm DFF_W1851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1920D));
DFF_save_fm DFF_W1852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1921D));
DFF_save_fm DFF_W1853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1922D));
DFF_save_fm DFF_W1854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1900E));
DFF_save_fm DFF_W1855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1901E));
DFF_save_fm DFF_W1856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1902E));
DFF_save_fm DFF_W1857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1910E));
DFF_save_fm DFF_W1858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1911E));
DFF_save_fm DFF_W1859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1912E));
DFF_save_fm DFF_W1860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1920E));
DFF_save_fm DFF_W1861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1921E));
DFF_save_fm DFF_W1862(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1922E));
DFF_save_fm DFF_W1863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1900F));
DFF_save_fm DFF_W1864(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1901F));
DFF_save_fm DFF_W1865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1902F));
DFF_save_fm DFF_W1866(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1910F));
DFF_save_fm DFF_W1867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1911F));
DFF_save_fm DFF_W1868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1912F));
DFF_save_fm DFF_W1869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1920F));
DFF_save_fm DFF_W1870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1921F));
DFF_save_fm DFF_W1871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1922F));
DFF_save_fm DFF_W1872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A000));
DFF_save_fm DFF_W1873(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A010));
DFF_save_fm DFF_W1874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A020));
DFF_save_fm DFF_W1875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A100));
DFF_save_fm DFF_W1876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A110));
DFF_save_fm DFF_W1877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A120));
DFF_save_fm DFF_W1878(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A200));
DFF_save_fm DFF_W1879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A210));
DFF_save_fm DFF_W1880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A220));
DFF_save_fm DFF_W1881(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A001));
DFF_save_fm DFF_W1882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A011));
DFF_save_fm DFF_W1883(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A021));
DFF_save_fm DFF_W1884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A101));
DFF_save_fm DFF_W1885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A111));
DFF_save_fm DFF_W1886(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A121));
DFF_save_fm DFF_W1887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A201));
DFF_save_fm DFF_W1888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A211));
DFF_save_fm DFF_W1889(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A221));
DFF_save_fm DFF_W1890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A002));
DFF_save_fm DFF_W1891(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A012));
DFF_save_fm DFF_W1892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A022));
DFF_save_fm DFF_W1893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A102));
DFF_save_fm DFF_W1894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A112));
DFF_save_fm DFF_W1895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A122));
DFF_save_fm DFF_W1896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A202));
DFF_save_fm DFF_W1897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A212));
DFF_save_fm DFF_W1898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A222));
DFF_save_fm DFF_W1899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A003));
DFF_save_fm DFF_W1900(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A013));
DFF_save_fm DFF_W1901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A023));
DFF_save_fm DFF_W1902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A103));
DFF_save_fm DFF_W1903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A113));
DFF_save_fm DFF_W1904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A123));
DFF_save_fm DFF_W1905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A203));
DFF_save_fm DFF_W1906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A213));
DFF_save_fm DFF_W1907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A223));
DFF_save_fm DFF_W1908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A004));
DFF_save_fm DFF_W1909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A014));
DFF_save_fm DFF_W1910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A024));
DFF_save_fm DFF_W1911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A104));
DFF_save_fm DFF_W1912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A114));
DFF_save_fm DFF_W1913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A124));
DFF_save_fm DFF_W1914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A204));
DFF_save_fm DFF_W1915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A214));
DFF_save_fm DFF_W1916(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A224));
DFF_save_fm DFF_W1917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A005));
DFF_save_fm DFF_W1918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A015));
DFF_save_fm DFF_W1919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A025));
DFF_save_fm DFF_W1920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A105));
DFF_save_fm DFF_W1921(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A115));
DFF_save_fm DFF_W1922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A125));
DFF_save_fm DFF_W1923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A205));
DFF_save_fm DFF_W1924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A215));
DFF_save_fm DFF_W1925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A225));
DFF_save_fm DFF_W1926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A006));
DFF_save_fm DFF_W1927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A016));
DFF_save_fm DFF_W1928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A026));
DFF_save_fm DFF_W1929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A106));
DFF_save_fm DFF_W1930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A116));
DFF_save_fm DFF_W1931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A126));
DFF_save_fm DFF_W1932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A206));
DFF_save_fm DFF_W1933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A216));
DFF_save_fm DFF_W1934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A226));
DFF_save_fm DFF_W1935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A007));
DFF_save_fm DFF_W1936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A017));
DFF_save_fm DFF_W1937(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A027));
DFF_save_fm DFF_W1938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A107));
DFF_save_fm DFF_W1939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A117));
DFF_save_fm DFF_W1940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A127));
DFF_save_fm DFF_W1941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A207));
DFF_save_fm DFF_W1942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A217));
DFF_save_fm DFF_W1943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A227));
DFF_save_fm DFF_W1944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A008));
DFF_save_fm DFF_W1945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A018));
DFF_save_fm DFF_W1946(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A028));
DFF_save_fm DFF_W1947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A108));
DFF_save_fm DFF_W1948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A118));
DFF_save_fm DFF_W1949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A128));
DFF_save_fm DFF_W1950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A208));
DFF_save_fm DFF_W1951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A218));
DFF_save_fm DFF_W1952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A228));
DFF_save_fm DFF_W1953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A009));
DFF_save_fm DFF_W1954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A019));
DFF_save_fm DFF_W1955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A029));
DFF_save_fm DFF_W1956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A109));
DFF_save_fm DFF_W1957(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A119));
DFF_save_fm DFF_W1958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A129));
DFF_save_fm DFF_W1959(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A209));
DFF_save_fm DFF_W1960(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A219));
DFF_save_fm DFF_W1961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A229));
DFF_save_fm DFF_W1962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A00A));
DFF_save_fm DFF_W1963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A01A));
DFF_save_fm DFF_W1964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A02A));
DFF_save_fm DFF_W1965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A10A));
DFF_save_fm DFF_W1966(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A11A));
DFF_save_fm DFF_W1967(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A12A));
DFF_save_fm DFF_W1968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A20A));
DFF_save_fm DFF_W1969(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A21A));
DFF_save_fm DFF_W1970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A22A));
DFF_save_fm DFF_W1971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A00B));
DFF_save_fm DFF_W1972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A01B));
DFF_save_fm DFF_W1973(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A02B));
DFF_save_fm DFF_W1974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A10B));
DFF_save_fm DFF_W1975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A11B));
DFF_save_fm DFF_W1976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A12B));
DFF_save_fm DFF_W1977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A20B));
DFF_save_fm DFF_W1978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A21B));
DFF_save_fm DFF_W1979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A22B));
DFF_save_fm DFF_W1980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A00C));
DFF_save_fm DFF_W1981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A01C));
DFF_save_fm DFF_W1982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A02C));
DFF_save_fm DFF_W1983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A10C));
DFF_save_fm DFF_W1984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A11C));
DFF_save_fm DFF_W1985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A12C));
DFF_save_fm DFF_W1986(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A20C));
DFF_save_fm DFF_W1987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A21C));
DFF_save_fm DFF_W1988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A22C));
DFF_save_fm DFF_W1989(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A00D));
DFF_save_fm DFF_W1990(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A01D));
DFF_save_fm DFF_W1991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A02D));
DFF_save_fm DFF_W1992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A10D));
DFF_save_fm DFF_W1993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A11D));
DFF_save_fm DFF_W1994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A12D));
DFF_save_fm DFF_W1995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A20D));
DFF_save_fm DFF_W1996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A21D));
DFF_save_fm DFF_W1997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A22D));
DFF_save_fm DFF_W1998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A00E));
DFF_save_fm DFF_W1999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A01E));
DFF_save_fm DFF_W2000(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A02E));
DFF_save_fm DFF_W2001(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A10E));
DFF_save_fm DFF_W2002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A11E));
DFF_save_fm DFF_W2003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A12E));
DFF_save_fm DFF_W2004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A20E));
DFF_save_fm DFF_W2005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A21E));
DFF_save_fm DFF_W2006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A22E));
DFF_save_fm DFF_W2007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A00F));
DFF_save_fm DFF_W2008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A01F));
DFF_save_fm DFF_W2009(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A02F));
DFF_save_fm DFF_W2010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A10F));
DFF_save_fm DFF_W2011(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A11F));
DFF_save_fm DFF_W2012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A12F));
DFF_save_fm DFF_W2013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A20F));
DFF_save_fm DFF_W2014(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A21F));
DFF_save_fm DFF_W2015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A22F));
DFF_save_fm DFF_W2016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B000));
DFF_save_fm DFF_W2017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B010));
DFF_save_fm DFF_W2018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B020));
DFF_save_fm DFF_W2019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B100));
DFF_save_fm DFF_W2020(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B110));
DFF_save_fm DFF_W2021(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B120));
DFF_save_fm DFF_W2022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B200));
DFF_save_fm DFF_W2023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B210));
DFF_save_fm DFF_W2024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B220));
DFF_save_fm DFF_W2025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B001));
DFF_save_fm DFF_W2026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B011));
DFF_save_fm DFF_W2027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B021));
DFF_save_fm DFF_W2028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B101));
DFF_save_fm DFF_W2029(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B111));
DFF_save_fm DFF_W2030(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B121));
DFF_save_fm DFF_W2031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B201));
DFF_save_fm DFF_W2032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B211));
DFF_save_fm DFF_W2033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B221));
DFF_save_fm DFF_W2034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B002));
DFF_save_fm DFF_W2035(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B012));
DFF_save_fm DFF_W2036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B022));
DFF_save_fm DFF_W2037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B102));
DFF_save_fm DFF_W2038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B112));
DFF_save_fm DFF_W2039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B122));
DFF_save_fm DFF_W2040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B202));
DFF_save_fm DFF_W2041(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B212));
DFF_save_fm DFF_W2042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B222));
DFF_save_fm DFF_W2043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B003));
DFF_save_fm DFF_W2044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B013));
DFF_save_fm DFF_W2045(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B023));
DFF_save_fm DFF_W2046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B103));
DFF_save_fm DFF_W2047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B113));
DFF_save_fm DFF_W2048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B123));
DFF_save_fm DFF_W2049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B203));
DFF_save_fm DFF_W2050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B213));
DFF_save_fm DFF_W2051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B223));
DFF_save_fm DFF_W2052(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B004));
DFF_save_fm DFF_W2053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B014));
DFF_save_fm DFF_W2054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B024));
DFF_save_fm DFF_W2055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B104));
DFF_save_fm DFF_W2056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B114));
DFF_save_fm DFF_W2057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B124));
DFF_save_fm DFF_W2058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B204));
DFF_save_fm DFF_W2059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B214));
DFF_save_fm DFF_W2060(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B224));
DFF_save_fm DFF_W2061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B005));
DFF_save_fm DFF_W2062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B015));
DFF_save_fm DFF_W2063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B025));
DFF_save_fm DFF_W2064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B105));
DFF_save_fm DFF_W2065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B115));
DFF_save_fm DFF_W2066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B125));
DFF_save_fm DFF_W2067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B205));
DFF_save_fm DFF_W2068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B215));
DFF_save_fm DFF_W2069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B225));
DFF_save_fm DFF_W2070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B006));
DFF_save_fm DFF_W2071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B016));
DFF_save_fm DFF_W2072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B026));
DFF_save_fm DFF_W2073(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B106));
DFF_save_fm DFF_W2074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B116));
DFF_save_fm DFF_W2075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B126));
DFF_save_fm DFF_W2076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B206));
DFF_save_fm DFF_W2077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B216));
DFF_save_fm DFF_W2078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B226));
DFF_save_fm DFF_W2079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B007));
DFF_save_fm DFF_W2080(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B017));
DFF_save_fm DFF_W2081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B027));
DFF_save_fm DFF_W2082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B107));
DFF_save_fm DFF_W2083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B117));
DFF_save_fm DFF_W2084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B127));
DFF_save_fm DFF_W2085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B207));
DFF_save_fm DFF_W2086(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B217));
DFF_save_fm DFF_W2087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B227));
DFF_save_fm DFF_W2088(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B008));
DFF_save_fm DFF_W2089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B018));
DFF_save_fm DFF_W2090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B028));
DFF_save_fm DFF_W2091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B108));
DFF_save_fm DFF_W2092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B118));
DFF_save_fm DFF_W2093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B128));
DFF_save_fm DFF_W2094(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B208));
DFF_save_fm DFF_W2095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B218));
DFF_save_fm DFF_W2096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B228));
DFF_save_fm DFF_W2097(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B009));
DFF_save_fm DFF_W2098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B019));
DFF_save_fm DFF_W2099(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B029));
DFF_save_fm DFF_W2100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B109));
DFF_save_fm DFF_W2101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B119));
DFF_save_fm DFF_W2102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B129));
DFF_save_fm DFF_W2103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B209));
DFF_save_fm DFF_W2104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B219));
DFF_save_fm DFF_W2105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B229));
DFF_save_fm DFF_W2106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B00A));
DFF_save_fm DFF_W2107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B01A));
DFF_save_fm DFF_W2108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B02A));
DFF_save_fm DFF_W2109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B10A));
DFF_save_fm DFF_W2110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B11A));
DFF_save_fm DFF_W2111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B12A));
DFF_save_fm DFF_W2112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B20A));
DFF_save_fm DFF_W2113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B21A));
DFF_save_fm DFF_W2114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B22A));
DFF_save_fm DFF_W2115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B00B));
DFF_save_fm DFF_W2116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B01B));
DFF_save_fm DFF_W2117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B02B));
DFF_save_fm DFF_W2118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B10B));
DFF_save_fm DFF_W2119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B11B));
DFF_save_fm DFF_W2120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B12B));
DFF_save_fm DFF_W2121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B20B));
DFF_save_fm DFF_W2122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B21B));
DFF_save_fm DFF_W2123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B22B));
DFF_save_fm DFF_W2124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B00C));
DFF_save_fm DFF_W2125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B01C));
DFF_save_fm DFF_W2126(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B02C));
DFF_save_fm DFF_W2127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B10C));
DFF_save_fm DFF_W2128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B11C));
DFF_save_fm DFF_W2129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B12C));
DFF_save_fm DFF_W2130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B20C));
DFF_save_fm DFF_W2131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B21C));
DFF_save_fm DFF_W2132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B22C));
DFF_save_fm DFF_W2133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B00D));
DFF_save_fm DFF_W2134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B01D));
DFF_save_fm DFF_W2135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B02D));
DFF_save_fm DFF_W2136(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B10D));
DFF_save_fm DFF_W2137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B11D));
DFF_save_fm DFF_W2138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B12D));
DFF_save_fm DFF_W2139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B20D));
DFF_save_fm DFF_W2140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B21D));
DFF_save_fm DFF_W2141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B22D));
DFF_save_fm DFF_W2142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B00E));
DFF_save_fm DFF_W2143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B01E));
DFF_save_fm DFF_W2144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B02E));
DFF_save_fm DFF_W2145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B10E));
DFF_save_fm DFF_W2146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B11E));
DFF_save_fm DFF_W2147(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B12E));
DFF_save_fm DFF_W2148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B20E));
DFF_save_fm DFF_W2149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B21E));
DFF_save_fm DFF_W2150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B22E));
DFF_save_fm DFF_W2151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B00F));
DFF_save_fm DFF_W2152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B01F));
DFF_save_fm DFF_W2153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B02F));
DFF_save_fm DFF_W2154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B10F));
DFF_save_fm DFF_W2155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B11F));
DFF_save_fm DFF_W2156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B12F));
DFF_save_fm DFF_W2157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B20F));
DFF_save_fm DFF_W2158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B21F));
DFF_save_fm DFF_W2159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B22F));
DFF_save_fm DFF_W2160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C000));
DFF_save_fm DFF_W2161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C010));
DFF_save_fm DFF_W2162(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C020));
DFF_save_fm DFF_W2163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C100));
DFF_save_fm DFF_W2164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C110));
DFF_save_fm DFF_W2165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C120));
DFF_save_fm DFF_W2166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C200));
DFF_save_fm DFF_W2167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C210));
DFF_save_fm DFF_W2168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C220));
DFF_save_fm DFF_W2169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C001));
DFF_save_fm DFF_W2170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C011));
DFF_save_fm DFF_W2171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C021));
DFF_save_fm DFF_W2172(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C101));
DFF_save_fm DFF_W2173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C111));
DFF_save_fm DFF_W2174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C121));
DFF_save_fm DFF_W2175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C201));
DFF_save_fm DFF_W2176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C211));
DFF_save_fm DFF_W2177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C221));
DFF_save_fm DFF_W2178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C002));
DFF_save_fm DFF_W2179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C012));
DFF_save_fm DFF_W2180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C022));
DFF_save_fm DFF_W2181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C102));
DFF_save_fm DFF_W2182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C112));
DFF_save_fm DFF_W2183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C122));
DFF_save_fm DFF_W2184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C202));
DFF_save_fm DFF_W2185(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C212));
DFF_save_fm DFF_W2186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C222));
DFF_save_fm DFF_W2187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C003));
DFF_save_fm DFF_W2188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C013));
DFF_save_fm DFF_W2189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C023));
DFF_save_fm DFF_W2190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C103));
DFF_save_fm DFF_W2191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C113));
DFF_save_fm DFF_W2192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C123));
DFF_save_fm DFF_W2193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C203));
DFF_save_fm DFF_W2194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C213));
DFF_save_fm DFF_W2195(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C223));
DFF_save_fm DFF_W2196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C004));
DFF_save_fm DFF_W2197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C014));
DFF_save_fm DFF_W2198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C024));
DFF_save_fm DFF_W2199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C104));
DFF_save_fm DFF_W2200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C114));
DFF_save_fm DFF_W2201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C124));
DFF_save_fm DFF_W2202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C204));
DFF_save_fm DFF_W2203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C214));
DFF_save_fm DFF_W2204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C224));
DFF_save_fm DFF_W2205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C005));
DFF_save_fm DFF_W2206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C015));
DFF_save_fm DFF_W2207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C025));
DFF_save_fm DFF_W2208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C105));
DFF_save_fm DFF_W2209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C115));
DFF_save_fm DFF_W2210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C125));
DFF_save_fm DFF_W2211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C205));
DFF_save_fm DFF_W2212(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C215));
DFF_save_fm DFF_W2213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C225));
DFF_save_fm DFF_W2214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C006));
DFF_save_fm DFF_W2215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C016));
DFF_save_fm DFF_W2216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C026));
DFF_save_fm DFF_W2217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C106));
DFF_save_fm DFF_W2218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C116));
DFF_save_fm DFF_W2219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C126));
DFF_save_fm DFF_W2220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C206));
DFF_save_fm DFF_W2221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C216));
DFF_save_fm DFF_W2222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C226));
DFF_save_fm DFF_W2223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C007));
DFF_save_fm DFF_W2224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C017));
DFF_save_fm DFF_W2225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C027));
DFF_save_fm DFF_W2226(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C107));
DFF_save_fm DFF_W2227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C117));
DFF_save_fm DFF_W2228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C127));
DFF_save_fm DFF_W2229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C207));
DFF_save_fm DFF_W2230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C217));
DFF_save_fm DFF_W2231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C227));
DFF_save_fm DFF_W2232(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C008));
DFF_save_fm DFF_W2233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C018));
DFF_save_fm DFF_W2234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C028));
DFF_save_fm DFF_W2235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C108));
DFF_save_fm DFF_W2236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C118));
DFF_save_fm DFF_W2237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C128));
DFF_save_fm DFF_W2238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C208));
DFF_save_fm DFF_W2239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C218));
DFF_save_fm DFF_W2240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C228));
DFF_save_fm DFF_W2241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C009));
DFF_save_fm DFF_W2242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C019));
DFF_save_fm DFF_W2243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C029));
DFF_save_fm DFF_W2244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C109));
DFF_save_fm DFF_W2245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C119));
DFF_save_fm DFF_W2246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C129));
DFF_save_fm DFF_W2247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C209));
DFF_save_fm DFF_W2248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C219));
DFF_save_fm DFF_W2249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C229));
DFF_save_fm DFF_W2250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C00A));
DFF_save_fm DFF_W2251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C01A));
DFF_save_fm DFF_W2252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C02A));
DFF_save_fm DFF_W2253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C10A));
DFF_save_fm DFF_W2254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C11A));
DFF_save_fm DFF_W2255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C12A));
DFF_save_fm DFF_W2256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C20A));
DFF_save_fm DFF_W2257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C21A));
DFF_save_fm DFF_W2258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C22A));
DFF_save_fm DFF_W2259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C00B));
DFF_save_fm DFF_W2260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C01B));
DFF_save_fm DFF_W2261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C02B));
DFF_save_fm DFF_W2262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C10B));
DFF_save_fm DFF_W2263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C11B));
DFF_save_fm DFF_W2264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C12B));
DFF_save_fm DFF_W2265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C20B));
DFF_save_fm DFF_W2266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C21B));
DFF_save_fm DFF_W2267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C22B));
DFF_save_fm DFF_W2268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C00C));
DFF_save_fm DFF_W2269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C01C));
DFF_save_fm DFF_W2270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C02C));
DFF_save_fm DFF_W2271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C10C));
DFF_save_fm DFF_W2272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C11C));
DFF_save_fm DFF_W2273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C12C));
DFF_save_fm DFF_W2274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C20C));
DFF_save_fm DFF_W2275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C21C));
DFF_save_fm DFF_W2276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C22C));
DFF_save_fm DFF_W2277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C00D));
DFF_save_fm DFF_W2278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C01D));
DFF_save_fm DFF_W2279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C02D));
DFF_save_fm DFF_W2280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C10D));
DFF_save_fm DFF_W2281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C11D));
DFF_save_fm DFF_W2282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C12D));
DFF_save_fm DFF_W2283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C20D));
DFF_save_fm DFF_W2284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C21D));
DFF_save_fm DFF_W2285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C22D));
DFF_save_fm DFF_W2286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C00E));
DFF_save_fm DFF_W2287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C01E));
DFF_save_fm DFF_W2288(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C02E));
DFF_save_fm DFF_W2289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C10E));
DFF_save_fm DFF_W2290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C11E));
DFF_save_fm DFF_W2291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C12E));
DFF_save_fm DFF_W2292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C20E));
DFF_save_fm DFF_W2293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C21E));
DFF_save_fm DFF_W2294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C22E));
DFF_save_fm DFF_W2295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C00F));
DFF_save_fm DFF_W2296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C01F));
DFF_save_fm DFF_W2297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C02F));
DFF_save_fm DFF_W2298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C10F));
DFF_save_fm DFF_W2299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C11F));
DFF_save_fm DFF_W2300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C12F));
DFF_save_fm DFF_W2301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C20F));
DFF_save_fm DFF_W2302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C21F));
DFF_save_fm DFF_W2303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C22F));
DFF_save_fm DFF_W2304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D000));
DFF_save_fm DFF_W2305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D010));
DFF_save_fm DFF_W2306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D020));
DFF_save_fm DFF_W2307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D100));
DFF_save_fm DFF_W2308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D110));
DFF_save_fm DFF_W2309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D120));
DFF_save_fm DFF_W2310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D200));
DFF_save_fm DFF_W2311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D210));
DFF_save_fm DFF_W2312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D220));
DFF_save_fm DFF_W2313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D001));
DFF_save_fm DFF_W2314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D011));
DFF_save_fm DFF_W2315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D021));
DFF_save_fm DFF_W2316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D101));
DFF_save_fm DFF_W2317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D111));
DFF_save_fm DFF_W2318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D121));
DFF_save_fm DFF_W2319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D201));
DFF_save_fm DFF_W2320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D211));
DFF_save_fm DFF_W2321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D221));
DFF_save_fm DFF_W2322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D002));
DFF_save_fm DFF_W2323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D012));
DFF_save_fm DFF_W2324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D022));
DFF_save_fm DFF_W2325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D102));
DFF_save_fm DFF_W2326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D112));
DFF_save_fm DFF_W2327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D122));
DFF_save_fm DFF_W2328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D202));
DFF_save_fm DFF_W2329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D212));
DFF_save_fm DFF_W2330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D222));
DFF_save_fm DFF_W2331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D003));
DFF_save_fm DFF_W2332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D013));
DFF_save_fm DFF_W2333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D023));
DFF_save_fm DFF_W2334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D103));
DFF_save_fm DFF_W2335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D113));
DFF_save_fm DFF_W2336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D123));
DFF_save_fm DFF_W2337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D203));
DFF_save_fm DFF_W2338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D213));
DFF_save_fm DFF_W2339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D223));
DFF_save_fm DFF_W2340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D004));
DFF_save_fm DFF_W2341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D014));
DFF_save_fm DFF_W2342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D024));
DFF_save_fm DFF_W2343(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D104));
DFF_save_fm DFF_W2344(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D114));
DFF_save_fm DFF_W2345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D124));
DFF_save_fm DFF_W2346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D204));
DFF_save_fm DFF_W2347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D214));
DFF_save_fm DFF_W2348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D224));
DFF_save_fm DFF_W2349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D005));
DFF_save_fm DFF_W2350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D015));
DFF_save_fm DFF_W2351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D025));
DFF_save_fm DFF_W2352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D105));
DFF_save_fm DFF_W2353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D115));
DFF_save_fm DFF_W2354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D125));
DFF_save_fm DFF_W2355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D205));
DFF_save_fm DFF_W2356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D215));
DFF_save_fm DFF_W2357(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D225));
DFF_save_fm DFF_W2358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D006));
DFF_save_fm DFF_W2359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D016));
DFF_save_fm DFF_W2360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D026));
DFF_save_fm DFF_W2361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D106));
DFF_save_fm DFF_W2362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D116));
DFF_save_fm DFF_W2363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D126));
DFF_save_fm DFF_W2364(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D206));
DFF_save_fm DFF_W2365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D216));
DFF_save_fm DFF_W2366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D226));
DFF_save_fm DFF_W2367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D007));
DFF_save_fm DFF_W2368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D017));
DFF_save_fm DFF_W2369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D027));
DFF_save_fm DFF_W2370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D107));
DFF_save_fm DFF_W2371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D117));
DFF_save_fm DFF_W2372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D127));
DFF_save_fm DFF_W2373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D207));
DFF_save_fm DFF_W2374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D217));
DFF_save_fm DFF_W2375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D227));
DFF_save_fm DFF_W2376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D008));
DFF_save_fm DFF_W2377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D018));
DFF_save_fm DFF_W2378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D028));
DFF_save_fm DFF_W2379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D108));
DFF_save_fm DFF_W2380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D118));
DFF_save_fm DFF_W2381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D128));
DFF_save_fm DFF_W2382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D208));
DFF_save_fm DFF_W2383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D218));
DFF_save_fm DFF_W2384(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D228));
DFF_save_fm DFF_W2385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D009));
DFF_save_fm DFF_W2386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D019));
DFF_save_fm DFF_W2387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D029));
DFF_save_fm DFF_W2388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D109));
DFF_save_fm DFF_W2389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D119));
DFF_save_fm DFF_W2390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D129));
DFF_save_fm DFF_W2391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D209));
DFF_save_fm DFF_W2392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D219));
DFF_save_fm DFF_W2393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D229));
DFF_save_fm DFF_W2394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D00A));
DFF_save_fm DFF_W2395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D01A));
DFF_save_fm DFF_W2396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D02A));
DFF_save_fm DFF_W2397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D10A));
DFF_save_fm DFF_W2398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D11A));
DFF_save_fm DFF_W2399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D12A));
DFF_save_fm DFF_W2400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D20A));
DFF_save_fm DFF_W2401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D21A));
DFF_save_fm DFF_W2402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D22A));
DFF_save_fm DFF_W2403(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D00B));
DFF_save_fm DFF_W2404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D01B));
DFF_save_fm DFF_W2405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D02B));
DFF_save_fm DFF_W2406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D10B));
DFF_save_fm DFF_W2407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D11B));
DFF_save_fm DFF_W2408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D12B));
DFF_save_fm DFF_W2409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D20B));
DFF_save_fm DFF_W2410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D21B));
DFF_save_fm DFF_W2411(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D22B));
DFF_save_fm DFF_W2412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D00C));
DFF_save_fm DFF_W2413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D01C));
DFF_save_fm DFF_W2414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D02C));
DFF_save_fm DFF_W2415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D10C));
DFF_save_fm DFF_W2416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D11C));
DFF_save_fm DFF_W2417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D12C));
DFF_save_fm DFF_W2418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D20C));
DFF_save_fm DFF_W2419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D21C));
DFF_save_fm DFF_W2420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D22C));
DFF_save_fm DFF_W2421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D00D));
DFF_save_fm DFF_W2422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D01D));
DFF_save_fm DFF_W2423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D02D));
DFF_save_fm DFF_W2424(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D10D));
DFF_save_fm DFF_W2425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D11D));
DFF_save_fm DFF_W2426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D12D));
DFF_save_fm DFF_W2427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D20D));
DFF_save_fm DFF_W2428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D21D));
DFF_save_fm DFF_W2429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D22D));
DFF_save_fm DFF_W2430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D00E));
DFF_save_fm DFF_W2431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D01E));
DFF_save_fm DFF_W2432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D02E));
DFF_save_fm DFF_W2433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D10E));
DFF_save_fm DFF_W2434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D11E));
DFF_save_fm DFF_W2435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D12E));
DFF_save_fm DFF_W2436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D20E));
DFF_save_fm DFF_W2437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D21E));
DFF_save_fm DFF_W2438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D22E));
DFF_save_fm DFF_W2439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D00F));
DFF_save_fm DFF_W2440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D01F));
DFF_save_fm DFF_W2441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D02F));
DFF_save_fm DFF_W2442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D10F));
DFF_save_fm DFF_W2443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D11F));
DFF_save_fm DFF_W2444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D12F));
DFF_save_fm DFF_W2445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D20F));
DFF_save_fm DFF_W2446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D21F));
DFF_save_fm DFF_W2447(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D22F));
DFF_save_fm DFF_W2448(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E000));
DFF_save_fm DFF_W2449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E010));
DFF_save_fm DFF_W2450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E020));
DFF_save_fm DFF_W2451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E100));
DFF_save_fm DFF_W2452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E110));
DFF_save_fm DFF_W2453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E120));
DFF_save_fm DFF_W2454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E200));
DFF_save_fm DFF_W2455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E210));
DFF_save_fm DFF_W2456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E220));
DFF_save_fm DFF_W2457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E001));
DFF_save_fm DFF_W2458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E011));
DFF_save_fm DFF_W2459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E021));
DFF_save_fm DFF_W2460(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E101));
DFF_save_fm DFF_W2461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E111));
DFF_save_fm DFF_W2462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E121));
DFF_save_fm DFF_W2463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E201));
DFF_save_fm DFF_W2464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E211));
DFF_save_fm DFF_W2465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E221));
DFF_save_fm DFF_W2466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E002));
DFF_save_fm DFF_W2467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E012));
DFF_save_fm DFF_W2468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E022));
DFF_save_fm DFF_W2469(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E102));
DFF_save_fm DFF_W2470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E112));
DFF_save_fm DFF_W2471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E122));
DFF_save_fm DFF_W2472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E202));
DFF_save_fm DFF_W2473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E212));
DFF_save_fm DFF_W2474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E222));
DFF_save_fm DFF_W2475(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E003));
DFF_save_fm DFF_W2476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E013));
DFF_save_fm DFF_W2477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E023));
DFF_save_fm DFF_W2478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E103));
DFF_save_fm DFF_W2479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E113));
DFF_save_fm DFF_W2480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E123));
DFF_save_fm DFF_W2481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E203));
DFF_save_fm DFF_W2482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E213));
DFF_save_fm DFF_W2483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E223));
DFF_save_fm DFF_W2484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E004));
DFF_save_fm DFF_W2485(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E014));
DFF_save_fm DFF_W2486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E024));
DFF_save_fm DFF_W2487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E104));
DFF_save_fm DFF_W2488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E114));
DFF_save_fm DFF_W2489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E124));
DFF_save_fm DFF_W2490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E204));
DFF_save_fm DFF_W2491(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E214));
DFF_save_fm DFF_W2492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E224));
DFF_save_fm DFF_W2493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E005));
DFF_save_fm DFF_W2494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E015));
DFF_save_fm DFF_W2495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E025));
DFF_save_fm DFF_W2496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E105));
DFF_save_fm DFF_W2497(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E115));
DFF_save_fm DFF_W2498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E125));
DFF_save_fm DFF_W2499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E205));
DFF_save_fm DFF_W2500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E215));
DFF_save_fm DFF_W2501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E225));
DFF_save_fm DFF_W2502(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E006));
DFF_save_fm DFF_W2503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E016));
DFF_save_fm DFF_W2504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E026));
DFF_save_fm DFF_W2505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E106));
DFF_save_fm DFF_W2506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E116));
DFF_save_fm DFF_W2507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E126));
DFF_save_fm DFF_W2508(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E206));
DFF_save_fm DFF_W2509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E216));
DFF_save_fm DFF_W2510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E226));
DFF_save_fm DFF_W2511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E007));
DFF_save_fm DFF_W2512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E017));
DFF_save_fm DFF_W2513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E027));
DFF_save_fm DFF_W2514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E107));
DFF_save_fm DFF_W2515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E117));
DFF_save_fm DFF_W2516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E127));
DFF_save_fm DFF_W2517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E207));
DFF_save_fm DFF_W2518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E217));
DFF_save_fm DFF_W2519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E227));
DFF_save_fm DFF_W2520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E008));
DFF_save_fm DFF_W2521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E018));
DFF_save_fm DFF_W2522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E028));
DFF_save_fm DFF_W2523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E108));
DFF_save_fm DFF_W2524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E118));
DFF_save_fm DFF_W2525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E128));
DFF_save_fm DFF_W2526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E208));
DFF_save_fm DFF_W2527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E218));
DFF_save_fm DFF_W2528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E228));
DFF_save_fm DFF_W2529(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E009));
DFF_save_fm DFF_W2530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E019));
DFF_save_fm DFF_W2531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E029));
DFF_save_fm DFF_W2532(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E109));
DFF_save_fm DFF_W2533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E119));
DFF_save_fm DFF_W2534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E129));
DFF_save_fm DFF_W2535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E209));
DFF_save_fm DFF_W2536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E219));
DFF_save_fm DFF_W2537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E229));
DFF_save_fm DFF_W2538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E00A));
DFF_save_fm DFF_W2539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E01A));
DFF_save_fm DFF_W2540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E02A));
DFF_save_fm DFF_W2541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E10A));
DFF_save_fm DFF_W2542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E11A));
DFF_save_fm DFF_W2543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E12A));
DFF_save_fm DFF_W2544(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E20A));
DFF_save_fm DFF_W2545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E21A));
DFF_save_fm DFF_W2546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E22A));
DFF_save_fm DFF_W2547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E00B));
DFF_save_fm DFF_W2548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E01B));
DFF_save_fm DFF_W2549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E02B));
DFF_save_fm DFF_W2550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E10B));
DFF_save_fm DFF_W2551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E11B));
DFF_save_fm DFF_W2552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E12B));
DFF_save_fm DFF_W2553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E20B));
DFF_save_fm DFF_W2554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E21B));
DFF_save_fm DFF_W2555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E22B));
DFF_save_fm DFF_W2556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E00C));
DFF_save_fm DFF_W2557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E01C));
DFF_save_fm DFF_W2558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E02C));
DFF_save_fm DFF_W2559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E10C));
DFF_save_fm DFF_W2560(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E11C));
DFF_save_fm DFF_W2561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E12C));
DFF_save_fm DFF_W2562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E20C));
DFF_save_fm DFF_W2563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E21C));
DFF_save_fm DFF_W2564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E22C));
DFF_save_fm DFF_W2565(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E00D));
DFF_save_fm DFF_W2566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E01D));
DFF_save_fm DFF_W2567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E02D));
DFF_save_fm DFF_W2568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E10D));
DFF_save_fm DFF_W2569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E11D));
DFF_save_fm DFF_W2570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E12D));
DFF_save_fm DFF_W2571(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E20D));
DFF_save_fm DFF_W2572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E21D));
DFF_save_fm DFF_W2573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E22D));
DFF_save_fm DFF_W2574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E00E));
DFF_save_fm DFF_W2575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E01E));
DFF_save_fm DFF_W2576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E02E));
DFF_save_fm DFF_W2577(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E10E));
DFF_save_fm DFF_W2578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E11E));
DFF_save_fm DFF_W2579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E12E));
DFF_save_fm DFF_W2580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E20E));
DFF_save_fm DFF_W2581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E21E));
DFF_save_fm DFF_W2582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E22E));
DFF_save_fm DFF_W2583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E00F));
DFF_save_fm DFF_W2584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E01F));
DFF_save_fm DFF_W2585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E02F));
DFF_save_fm DFF_W2586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E10F));
DFF_save_fm DFF_W2587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E11F));
DFF_save_fm DFF_W2588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E12F));
DFF_save_fm DFF_W2589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E20F));
DFF_save_fm DFF_W2590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E21F));
DFF_save_fm DFF_W2591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E22F));
DFF_save_fm DFF_W2592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F000));
DFF_save_fm DFF_W2593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F010));
DFF_save_fm DFF_W2594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F020));
DFF_save_fm DFF_W2595(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F100));
DFF_save_fm DFF_W2596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F110));
DFF_save_fm DFF_W2597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F120));
DFF_save_fm DFF_W2598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F200));
DFF_save_fm DFF_W2599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F210));
DFF_save_fm DFF_W2600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F220));
DFF_save_fm DFF_W2601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F001));
DFF_save_fm DFF_W2602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F011));
DFF_save_fm DFF_W2603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F021));
DFF_save_fm DFF_W2604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F101));
DFF_save_fm DFF_W2605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F111));
DFF_save_fm DFF_W2606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F121));
DFF_save_fm DFF_W2607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F201));
DFF_save_fm DFF_W2608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F211));
DFF_save_fm DFF_W2609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F221));
DFF_save_fm DFF_W2610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F002));
DFF_save_fm DFF_W2611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F012));
DFF_save_fm DFF_W2612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F022));
DFF_save_fm DFF_W2613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F102));
DFF_save_fm DFF_W2614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F112));
DFF_save_fm DFF_W2615(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F122));
DFF_save_fm DFF_W2616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F202));
DFF_save_fm DFF_W2617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F212));
DFF_save_fm DFF_W2618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F222));
DFF_save_fm DFF_W2619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F003));
DFF_save_fm DFF_W2620(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F013));
DFF_save_fm DFF_W2621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F023));
DFF_save_fm DFF_W2622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F103));
DFF_save_fm DFF_W2623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F113));
DFF_save_fm DFF_W2624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F123));
DFF_save_fm DFF_W2625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F203));
DFF_save_fm DFF_W2626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F213));
DFF_save_fm DFF_W2627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F223));
DFF_save_fm DFF_W2628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F004));
DFF_save_fm DFF_W2629(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F014));
DFF_save_fm DFF_W2630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F024));
DFF_save_fm DFF_W2631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F104));
DFF_save_fm DFF_W2632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F114));
DFF_save_fm DFF_W2633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F124));
DFF_save_fm DFF_W2634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F204));
DFF_save_fm DFF_W2635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F214));
DFF_save_fm DFF_W2636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F224));
DFF_save_fm DFF_W2637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F005));
DFF_save_fm DFF_W2638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F015));
DFF_save_fm DFF_W2639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F025));
DFF_save_fm DFF_W2640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F105));
DFF_save_fm DFF_W2641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F115));
DFF_save_fm DFF_W2642(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F125));
DFF_save_fm DFF_W2643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F205));
DFF_save_fm DFF_W2644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F215));
DFF_save_fm DFF_W2645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F225));
DFF_save_fm DFF_W2646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F006));
DFF_save_fm DFF_W2647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F016));
DFF_save_fm DFF_W2648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F026));
DFF_save_fm DFF_W2649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F106));
DFF_save_fm DFF_W2650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F116));
DFF_save_fm DFF_W2651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F126));
DFF_save_fm DFF_W2652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F206));
DFF_save_fm DFF_W2653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F216));
DFF_save_fm DFF_W2654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F226));
DFF_save_fm DFF_W2655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F007));
DFF_save_fm DFF_W2656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F017));
DFF_save_fm DFF_W2657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F027));
DFF_save_fm DFF_W2658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F107));
DFF_save_fm DFF_W2659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F117));
DFF_save_fm DFF_W2660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F127));
DFF_save_fm DFF_W2661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F207));
DFF_save_fm DFF_W2662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F217));
DFF_save_fm DFF_W2663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F227));
DFF_save_fm DFF_W2664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F008));
DFF_save_fm DFF_W2665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F018));
DFF_save_fm DFF_W2666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F028));
DFF_save_fm DFF_W2667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F108));
DFF_save_fm DFF_W2668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F118));
DFF_save_fm DFF_W2669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F128));
DFF_save_fm DFF_W2670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F208));
DFF_save_fm DFF_W2671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F218));
DFF_save_fm DFF_W2672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F228));
DFF_save_fm DFF_W2673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F009));
DFF_save_fm DFF_W2674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F019));
DFF_save_fm DFF_W2675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F029));
DFF_save_fm DFF_W2676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F109));
DFF_save_fm DFF_W2677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F119));
DFF_save_fm DFF_W2678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F129));
DFF_save_fm DFF_W2679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F209));
DFF_save_fm DFF_W2680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F219));
DFF_save_fm DFF_W2681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F229));
DFF_save_fm DFF_W2682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F00A));
DFF_save_fm DFF_W2683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F01A));
DFF_save_fm DFF_W2684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F02A));
DFF_save_fm DFF_W2685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F10A));
DFF_save_fm DFF_W2686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F11A));
DFF_save_fm DFF_W2687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F12A));
DFF_save_fm DFF_W2688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F20A));
DFF_save_fm DFF_W2689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F21A));
DFF_save_fm DFF_W2690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F22A));
DFF_save_fm DFF_W2691(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F00B));
DFF_save_fm DFF_W2692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F01B));
DFF_save_fm DFF_W2693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F02B));
DFF_save_fm DFF_W2694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F10B));
DFF_save_fm DFF_W2695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F11B));
DFF_save_fm DFF_W2696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F12B));
DFF_save_fm DFF_W2697(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F20B));
DFF_save_fm DFF_W2698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F21B));
DFF_save_fm DFF_W2699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F22B));
DFF_save_fm DFF_W2700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F00C));
DFF_save_fm DFF_W2701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F01C));
DFF_save_fm DFF_W2702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F02C));
DFF_save_fm DFF_W2703(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F10C));
DFF_save_fm DFF_W2704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F11C));
DFF_save_fm DFF_W2705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F12C));
DFF_save_fm DFF_W2706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F20C));
DFF_save_fm DFF_W2707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F21C));
DFF_save_fm DFF_W2708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F22C));
DFF_save_fm DFF_W2709(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F00D));
DFF_save_fm DFF_W2710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F01D));
DFF_save_fm DFF_W2711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F02D));
DFF_save_fm DFF_W2712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F10D));
DFF_save_fm DFF_W2713(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F11D));
DFF_save_fm DFF_W2714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F12D));
DFF_save_fm DFF_W2715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F20D));
DFF_save_fm DFF_W2716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F21D));
DFF_save_fm DFF_W2717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F22D));
DFF_save_fm DFF_W2718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F00E));
DFF_save_fm DFF_W2719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F01E));
DFF_save_fm DFF_W2720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F02E));
DFF_save_fm DFF_W2721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F10E));
DFF_save_fm DFF_W2722(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F11E));
DFF_save_fm DFF_W2723(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F12E));
DFF_save_fm DFF_W2724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F20E));
DFF_save_fm DFF_W2725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F21E));
DFF_save_fm DFF_W2726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F22E));
DFF_save_fm DFF_W2727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F00F));
DFF_save_fm DFF_W2728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F01F));
DFF_save_fm DFF_W2729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F02F));
DFF_save_fm DFF_W2730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F10F));
DFF_save_fm DFF_W2731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F11F));
DFF_save_fm DFF_W2732(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F12F));
DFF_save_fm DFF_W2733(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F20F));
DFF_save_fm DFF_W2734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F21F));
DFF_save_fm DFF_W2735(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F22F));
DFF_save_fm DFF_W2736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G000));
DFF_save_fm DFF_W2737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G010));
DFF_save_fm DFF_W2738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G020));
DFF_save_fm DFF_W2739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G100));
DFF_save_fm DFF_W2740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G110));
DFF_save_fm DFF_W2741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G120));
DFF_save_fm DFF_W2742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G200));
DFF_save_fm DFF_W2743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G210));
DFF_save_fm DFF_W2744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G220));
DFF_save_fm DFF_W2745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G001));
DFF_save_fm DFF_W2746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G011));
DFF_save_fm DFF_W2747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G021));
DFF_save_fm DFF_W2748(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G101));
DFF_save_fm DFF_W2749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G111));
DFF_save_fm DFF_W2750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G121));
DFF_save_fm DFF_W2751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G201));
DFF_save_fm DFF_W2752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G211));
DFF_save_fm DFF_W2753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G221));
DFF_save_fm DFF_W2754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G002));
DFF_save_fm DFF_W2755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G012));
DFF_save_fm DFF_W2756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G022));
DFF_save_fm DFF_W2757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G102));
DFF_save_fm DFF_W2758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G112));
DFF_save_fm DFF_W2759(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G122));
DFF_save_fm DFF_W2760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G202));
DFF_save_fm DFF_W2761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G212));
DFF_save_fm DFF_W2762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G222));
DFF_save_fm DFF_W2763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G003));
DFF_save_fm DFF_W2764(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G013));
DFF_save_fm DFF_W2765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G023));
DFF_save_fm DFF_W2766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G103));
DFF_save_fm DFF_W2767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G113));
DFF_save_fm DFF_W2768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G123));
DFF_save_fm DFF_W2769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G203));
DFF_save_fm DFF_W2770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G213));
DFF_save_fm DFF_W2771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G223));
DFF_save_fm DFF_W2772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G004));
DFF_save_fm DFF_W2773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G014));
DFF_save_fm DFF_W2774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G024));
DFF_save_fm DFF_W2775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G104));
DFF_save_fm DFF_W2776(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G114));
DFF_save_fm DFF_W2777(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G124));
DFF_save_fm DFF_W2778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G204));
DFF_save_fm DFF_W2779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G214));
DFF_save_fm DFF_W2780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G224));
DFF_save_fm DFF_W2781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G005));
DFF_save_fm DFF_W2782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G015));
DFF_save_fm DFF_W2783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G025));
DFF_save_fm DFF_W2784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G105));
DFF_save_fm DFF_W2785(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G115));
DFF_save_fm DFF_W2786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G125));
DFF_save_fm DFF_W2787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G205));
DFF_save_fm DFF_W2788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G215));
DFF_save_fm DFF_W2789(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G225));
DFF_save_fm DFF_W2790(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G006));
DFF_save_fm DFF_W2791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G016));
DFF_save_fm DFF_W2792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G026));
DFF_save_fm DFF_W2793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G106));
DFF_save_fm DFF_W2794(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G116));
DFF_save_fm DFF_W2795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G126));
DFF_save_fm DFF_W2796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G206));
DFF_save_fm DFF_W2797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G216));
DFF_save_fm DFF_W2798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G226));
DFF_save_fm DFF_W2799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G007));
DFF_save_fm DFF_W2800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G017));
DFF_save_fm DFF_W2801(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G027));
DFF_save_fm DFF_W2802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G107));
DFF_save_fm DFF_W2803(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G117));
DFF_save_fm DFF_W2804(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G127));
DFF_save_fm DFF_W2805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G207));
DFF_save_fm DFF_W2806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G217));
DFF_save_fm DFF_W2807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G227));
DFF_save_fm DFF_W2808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G008));
DFF_save_fm DFF_W2809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G018));
DFF_save_fm DFF_W2810(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G028));
DFF_save_fm DFF_W2811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G108));
DFF_save_fm DFF_W2812(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G118));
DFF_save_fm DFF_W2813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G128));
DFF_save_fm DFF_W2814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G208));
DFF_save_fm DFF_W2815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G218));
DFF_save_fm DFF_W2816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G228));
DFF_save_fm DFF_W2817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G009));
DFF_save_fm DFF_W2818(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G019));
DFF_save_fm DFF_W2819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G029));
DFF_save_fm DFF_W2820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G109));
DFF_save_fm DFF_W2821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G119));
DFF_save_fm DFF_W2822(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G129));
DFF_save_fm DFF_W2823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G209));
DFF_save_fm DFF_W2824(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G219));
DFF_save_fm DFF_W2825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G229));
DFF_save_fm DFF_W2826(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G00A));
DFF_save_fm DFF_W2827(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G01A));
DFF_save_fm DFF_W2828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G02A));
DFF_save_fm DFF_W2829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G10A));
DFF_save_fm DFF_W2830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G11A));
DFF_save_fm DFF_W2831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G12A));
DFF_save_fm DFF_W2832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G20A));
DFF_save_fm DFF_W2833(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G21A));
DFF_save_fm DFF_W2834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G22A));
DFF_save_fm DFF_W2835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G00B));
DFF_save_fm DFF_W2836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G01B));
DFF_save_fm DFF_W2837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G02B));
DFF_save_fm DFF_W2838(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G10B));
DFF_save_fm DFF_W2839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G11B));
DFF_save_fm DFF_W2840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G12B));
DFF_save_fm DFF_W2841(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G20B));
DFF_save_fm DFF_W2842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G21B));
DFF_save_fm DFF_W2843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G22B));
DFF_save_fm DFF_W2844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G00C));
DFF_save_fm DFF_W2845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G01C));
DFF_save_fm DFF_W2846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G02C));
DFF_save_fm DFF_W2847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G10C));
DFF_save_fm DFF_W2848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G11C));
DFF_save_fm DFF_W2849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G12C));
DFF_save_fm DFF_W2850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G20C));
DFF_save_fm DFF_W2851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G21C));
DFF_save_fm DFF_W2852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G22C));
DFF_save_fm DFF_W2853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G00D));
DFF_save_fm DFF_W2854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G01D));
DFF_save_fm DFF_W2855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G02D));
DFF_save_fm DFF_W2856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G10D));
DFF_save_fm DFF_W2857(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G11D));
DFF_save_fm DFF_W2858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G12D));
DFF_save_fm DFF_W2859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G20D));
DFF_save_fm DFF_W2860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G21D));
DFF_save_fm DFF_W2861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G22D));
DFF_save_fm DFF_W2862(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G00E));
DFF_save_fm DFF_W2863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G01E));
DFF_save_fm DFF_W2864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G02E));
DFF_save_fm DFF_W2865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G10E));
DFF_save_fm DFF_W2866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G11E));
DFF_save_fm DFF_W2867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G12E));
DFF_save_fm DFF_W2868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G20E));
DFF_save_fm DFF_W2869(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G21E));
DFF_save_fm DFF_W2870(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G22E));
DFF_save_fm DFF_W2871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G00F));
DFF_save_fm DFF_W2872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G01F));
DFF_save_fm DFF_W2873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G02F));
DFF_save_fm DFF_W2874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G10F));
DFF_save_fm DFF_W2875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G11F));
DFF_save_fm DFF_W2876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G12F));
DFF_save_fm DFF_W2877(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1G20F));
DFF_save_fm DFF_W2878(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G21F));
DFF_save_fm DFF_W2879(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1G22F));
DFF_save_fm DFF_W2880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H000));
DFF_save_fm DFF_W2881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H010));
DFF_save_fm DFF_W2882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H020));
DFF_save_fm DFF_W2883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H100));
DFF_save_fm DFF_W2884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H110));
DFF_save_fm DFF_W2885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H120));
DFF_save_fm DFF_W2886(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H200));
DFF_save_fm DFF_W2887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H210));
DFF_save_fm DFF_W2888(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H220));
DFF_save_fm DFF_W2889(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H001));
DFF_save_fm DFF_W2890(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H011));
DFF_save_fm DFF_W2891(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H021));
DFF_save_fm DFF_W2892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H101));
DFF_save_fm DFF_W2893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H111));
DFF_save_fm DFF_W2894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H121));
DFF_save_fm DFF_W2895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H201));
DFF_save_fm DFF_W2896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H211));
DFF_save_fm DFF_W2897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H221));
DFF_save_fm DFF_W2898(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H002));
DFF_save_fm DFF_W2899(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H012));
DFF_save_fm DFF_W2900(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H022));
DFF_save_fm DFF_W2901(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H102));
DFF_save_fm DFF_W2902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H112));
DFF_save_fm DFF_W2903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H122));
DFF_save_fm DFF_W2904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H202));
DFF_save_fm DFF_W2905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H212));
DFF_save_fm DFF_W2906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H222));
DFF_save_fm DFF_W2907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H003));
DFF_save_fm DFF_W2908(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H013));
DFF_save_fm DFF_W2909(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H023));
DFF_save_fm DFF_W2910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H103));
DFF_save_fm DFF_W2911(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H113));
DFF_save_fm DFF_W2912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H123));
DFF_save_fm DFF_W2913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H203));
DFF_save_fm DFF_W2914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H213));
DFF_save_fm DFF_W2915(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H223));
DFF_save_fm DFF_W2916(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H004));
DFF_save_fm DFF_W2917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H014));
DFF_save_fm DFF_W2918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H024));
DFF_save_fm DFF_W2919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H104));
DFF_save_fm DFF_W2920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H114));
DFF_save_fm DFF_W2921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H124));
DFF_save_fm DFF_W2922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H204));
DFF_save_fm DFF_W2923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H214));
DFF_save_fm DFF_W2924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H224));
DFF_save_fm DFF_W2925(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H005));
DFF_save_fm DFF_W2926(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H015));
DFF_save_fm DFF_W2927(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H025));
DFF_save_fm DFF_W2928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H105));
DFF_save_fm DFF_W2929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H115));
DFF_save_fm DFF_W2930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H125));
DFF_save_fm DFF_W2931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H205));
DFF_save_fm DFF_W2932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H215));
DFF_save_fm DFF_W2933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H225));
DFF_save_fm DFF_W2934(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H006));
DFF_save_fm DFF_W2935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H016));
DFF_save_fm DFF_W2936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H026));
DFF_save_fm DFF_W2937(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H106));
DFF_save_fm DFF_W2938(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H116));
DFF_save_fm DFF_W2939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H126));
DFF_save_fm DFF_W2940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H206));
DFF_save_fm DFF_W2941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H216));
DFF_save_fm DFF_W2942(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H226));
DFF_save_fm DFF_W2943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H007));
DFF_save_fm DFF_W2944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H017));
DFF_save_fm DFF_W2945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H027));
DFF_save_fm DFF_W2946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H107));
DFF_save_fm DFF_W2947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H117));
DFF_save_fm DFF_W2948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H127));
DFF_save_fm DFF_W2949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H207));
DFF_save_fm DFF_W2950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H217));
DFF_save_fm DFF_W2951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H227));
DFF_save_fm DFF_W2952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H008));
DFF_save_fm DFF_W2953(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H018));
DFF_save_fm DFF_W2954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H028));
DFF_save_fm DFF_W2955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H108));
DFF_save_fm DFF_W2956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H118));
DFF_save_fm DFF_W2957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H128));
DFF_save_fm DFF_W2958(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H208));
DFF_save_fm DFF_W2959(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H218));
DFF_save_fm DFF_W2960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H228));
DFF_save_fm DFF_W2961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H009));
DFF_save_fm DFF_W2962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H019));
DFF_save_fm DFF_W2963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H029));
DFF_save_fm DFF_W2964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H109));
DFF_save_fm DFF_W2965(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H119));
DFF_save_fm DFF_W2966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H129));
DFF_save_fm DFF_W2967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H209));
DFF_save_fm DFF_W2968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H219));
DFF_save_fm DFF_W2969(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H229));
DFF_save_fm DFF_W2970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H00A));
DFF_save_fm DFF_W2971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H01A));
DFF_save_fm DFF_W2972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H02A));
DFF_save_fm DFF_W2973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H10A));
DFF_save_fm DFF_W2974(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H11A));
DFF_save_fm DFF_W2975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H12A));
DFF_save_fm DFF_W2976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H20A));
DFF_save_fm DFF_W2977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H21A));
DFF_save_fm DFF_W2978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H22A));
DFF_save_fm DFF_W2979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H00B));
DFF_save_fm DFF_W2980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H01B));
DFF_save_fm DFF_W2981(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H02B));
DFF_save_fm DFF_W2982(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H10B));
DFF_save_fm DFF_W2983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H11B));
DFF_save_fm DFF_W2984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H12B));
DFF_save_fm DFF_W2985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H20B));
DFF_save_fm DFF_W2986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H21B));
DFF_save_fm DFF_W2987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H22B));
DFF_save_fm DFF_W2988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H00C));
DFF_save_fm DFF_W2989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H01C));
DFF_save_fm DFF_W2990(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H02C));
DFF_save_fm DFF_W2991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H10C));
DFF_save_fm DFF_W2992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H11C));
DFF_save_fm DFF_W2993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H12C));
DFF_save_fm DFF_W2994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H20C));
DFF_save_fm DFF_W2995(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H21C));
DFF_save_fm DFF_W2996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H22C));
DFF_save_fm DFF_W2997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H00D));
DFF_save_fm DFF_W2998(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H01D));
DFF_save_fm DFF_W2999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H02D));
DFF_save_fm DFF_W3000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H10D));
DFF_save_fm DFF_W3001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H11D));
DFF_save_fm DFF_W3002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H12D));
DFF_save_fm DFF_W3003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H20D));
DFF_save_fm DFF_W3004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H21D));
DFF_save_fm DFF_W3005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H22D));
DFF_save_fm DFF_W3006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H00E));
DFF_save_fm DFF_W3007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H01E));
DFF_save_fm DFF_W3008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H02E));
DFF_save_fm DFF_W3009(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H10E));
DFF_save_fm DFF_W3010(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H11E));
DFF_save_fm DFF_W3011(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H12E));
DFF_save_fm DFF_W3012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H20E));
DFF_save_fm DFF_W3013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H21E));
DFF_save_fm DFF_W3014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H22E));
DFF_save_fm DFF_W3015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H00F));
DFF_save_fm DFF_W3016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H01F));
DFF_save_fm DFF_W3017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H02F));
DFF_save_fm DFF_W3018(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H10F));
DFF_save_fm DFF_W3019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H11F));
DFF_save_fm DFF_W3020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H12F));
DFF_save_fm DFF_W3021(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1H20F));
DFF_save_fm DFF_W3022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H21F));
DFF_save_fm DFF_W3023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1H22F));
DFF_save_fm DFF_W3024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I000));
DFF_save_fm DFF_W3025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I010));
DFF_save_fm DFF_W3026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I020));
DFF_save_fm DFF_W3027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I100));
DFF_save_fm DFF_W3028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I110));
DFF_save_fm DFF_W3029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I120));
DFF_save_fm DFF_W3030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I200));
DFF_save_fm DFF_W3031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I210));
DFF_save_fm DFF_W3032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I220));
DFF_save_fm DFF_W3033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I001));
DFF_save_fm DFF_W3034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I011));
DFF_save_fm DFF_W3035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I021));
DFF_save_fm DFF_W3036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I101));
DFF_save_fm DFF_W3037(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I111));
DFF_save_fm DFF_W3038(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I121));
DFF_save_fm DFF_W3039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I201));
DFF_save_fm DFF_W3040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I211));
DFF_save_fm DFF_W3041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I221));
DFF_save_fm DFF_W3042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I002));
DFF_save_fm DFF_W3043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I012));
DFF_save_fm DFF_W3044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I022));
DFF_save_fm DFF_W3045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I102));
DFF_save_fm DFF_W3046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I112));
DFF_save_fm DFF_W3047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I122));
DFF_save_fm DFF_W3048(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I202));
DFF_save_fm DFF_W3049(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I212));
DFF_save_fm DFF_W3050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I222));
DFF_save_fm DFF_W3051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I003));
DFF_save_fm DFF_W3052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I013));
DFF_save_fm DFF_W3053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I023));
DFF_save_fm DFF_W3054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I103));
DFF_save_fm DFF_W3055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I113));
DFF_save_fm DFF_W3056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I123));
DFF_save_fm DFF_W3057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I203));
DFF_save_fm DFF_W3058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I213));
DFF_save_fm DFF_W3059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I223));
DFF_save_fm DFF_W3060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I004));
DFF_save_fm DFF_W3061(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I014));
DFF_save_fm DFF_W3062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I024));
DFF_save_fm DFF_W3063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I104));
DFF_save_fm DFF_W3064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I114));
DFF_save_fm DFF_W3065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I124));
DFF_save_fm DFF_W3066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I204));
DFF_save_fm DFF_W3067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I214));
DFF_save_fm DFF_W3068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I224));
DFF_save_fm DFF_W3069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I005));
DFF_save_fm DFF_W3070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I015));
DFF_save_fm DFF_W3071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I025));
DFF_save_fm DFF_W3072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I105));
DFF_save_fm DFF_W3073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I115));
DFF_save_fm DFF_W3074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I125));
DFF_save_fm DFF_W3075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I205));
DFF_save_fm DFF_W3076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I215));
DFF_save_fm DFF_W3077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I225));
DFF_save_fm DFF_W3078(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I006));
DFF_save_fm DFF_W3079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I016));
DFF_save_fm DFF_W3080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I026));
DFF_save_fm DFF_W3081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I106));
DFF_save_fm DFF_W3082(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I116));
DFF_save_fm DFF_W3083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I126));
DFF_save_fm DFF_W3084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I206));
DFF_save_fm DFF_W3085(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I216));
DFF_save_fm DFF_W3086(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I226));
DFF_save_fm DFF_W3087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I007));
DFF_save_fm DFF_W3088(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I017));
DFF_save_fm DFF_W3089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I027));
DFF_save_fm DFF_W3090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I107));
DFF_save_fm DFF_W3091(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I117));
DFF_save_fm DFF_W3092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I127));
DFF_save_fm DFF_W3093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I207));
DFF_save_fm DFF_W3094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I217));
DFF_save_fm DFF_W3095(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I227));
DFF_save_fm DFF_W3096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I008));
DFF_save_fm DFF_W3097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I018));
DFF_save_fm DFF_W3098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I028));
DFF_save_fm DFF_W3099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I108));
DFF_save_fm DFF_W3100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I118));
DFF_save_fm DFF_W3101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I128));
DFF_save_fm DFF_W3102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I208));
DFF_save_fm DFF_W3103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I218));
DFF_save_fm DFF_W3104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I228));
DFF_save_fm DFF_W3105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I009));
DFF_save_fm DFF_W3106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I019));
DFF_save_fm DFF_W3107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I029));
DFF_save_fm DFF_W3108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I109));
DFF_save_fm DFF_W3109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I119));
DFF_save_fm DFF_W3110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I129));
DFF_save_fm DFF_W3111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I209));
DFF_save_fm DFF_W3112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I219));
DFF_save_fm DFF_W3113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I229));
DFF_save_fm DFF_W3114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I00A));
DFF_save_fm DFF_W3115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I01A));
DFF_save_fm DFF_W3116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I02A));
DFF_save_fm DFF_W3117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I10A));
DFF_save_fm DFF_W3118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I11A));
DFF_save_fm DFF_W3119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I12A));
DFF_save_fm DFF_W3120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I20A));
DFF_save_fm DFF_W3121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I21A));
DFF_save_fm DFF_W3122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I22A));
DFF_save_fm DFF_W3123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I00B));
DFF_save_fm DFF_W3124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I01B));
DFF_save_fm DFF_W3125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I02B));
DFF_save_fm DFF_W3126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I10B));
DFF_save_fm DFF_W3127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I11B));
DFF_save_fm DFF_W3128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I12B));
DFF_save_fm DFF_W3129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I20B));
DFF_save_fm DFF_W3130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I21B));
DFF_save_fm DFF_W3131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I22B));
DFF_save_fm DFF_W3132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I00C));
DFF_save_fm DFF_W3133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I01C));
DFF_save_fm DFF_W3134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I02C));
DFF_save_fm DFF_W3135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I10C));
DFF_save_fm DFF_W3136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I11C));
DFF_save_fm DFF_W3137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I12C));
DFF_save_fm DFF_W3138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I20C));
DFF_save_fm DFF_W3139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I21C));
DFF_save_fm DFF_W3140(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I22C));
DFF_save_fm DFF_W3141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I00D));
DFF_save_fm DFF_W3142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I01D));
DFF_save_fm DFF_W3143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I02D));
DFF_save_fm DFF_W3144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I10D));
DFF_save_fm DFF_W3145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I11D));
DFF_save_fm DFF_W3146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I12D));
DFF_save_fm DFF_W3147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I20D));
DFF_save_fm DFF_W3148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I21D));
DFF_save_fm DFF_W3149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I22D));
DFF_save_fm DFF_W3150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I00E));
DFF_save_fm DFF_W3151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I01E));
DFF_save_fm DFF_W3152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I02E));
DFF_save_fm DFF_W3153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I10E));
DFF_save_fm DFF_W3154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I11E));
DFF_save_fm DFF_W3155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I12E));
DFF_save_fm DFF_W3156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I20E));
DFF_save_fm DFF_W3157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I21E));
DFF_save_fm DFF_W3158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I22E));
DFF_save_fm DFF_W3159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I00F));
DFF_save_fm DFF_W3160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I01F));
DFF_save_fm DFF_W3161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I02F));
DFF_save_fm DFF_W3162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I10F));
DFF_save_fm DFF_W3163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I11F));
DFF_save_fm DFF_W3164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I12F));
DFF_save_fm DFF_W3165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1I20F));
DFF_save_fm DFF_W3166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I21F));
DFF_save_fm DFF_W3167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1I22F));
DFF_save_fm DFF_W3168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J000));
DFF_save_fm DFF_W3169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J010));
DFF_save_fm DFF_W3170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J020));
DFF_save_fm DFF_W3171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J100));
DFF_save_fm DFF_W3172(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J110));
DFF_save_fm DFF_W3173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J120));
DFF_save_fm DFF_W3174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J200));
DFF_save_fm DFF_W3175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J210));
DFF_save_fm DFF_W3176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J220));
DFF_save_fm DFF_W3177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J001));
DFF_save_fm DFF_W3178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J011));
DFF_save_fm DFF_W3179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J021));
DFF_save_fm DFF_W3180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J101));
DFF_save_fm DFF_W3181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J111));
DFF_save_fm DFF_W3182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J121));
DFF_save_fm DFF_W3183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J201));
DFF_save_fm DFF_W3184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J211));
DFF_save_fm DFF_W3185(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J221));
DFF_save_fm DFF_W3186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J002));
DFF_save_fm DFF_W3187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J012));
DFF_save_fm DFF_W3188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J022));
DFF_save_fm DFF_W3189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J102));
DFF_save_fm DFF_W3190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J112));
DFF_save_fm DFF_W3191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J122));
DFF_save_fm DFF_W3192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J202));
DFF_save_fm DFF_W3193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J212));
DFF_save_fm DFF_W3194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J222));
DFF_save_fm DFF_W3195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J003));
DFF_save_fm DFF_W3196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J013));
DFF_save_fm DFF_W3197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J023));
DFF_save_fm DFF_W3198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J103));
DFF_save_fm DFF_W3199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J113));
DFF_save_fm DFF_W3200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J123));
DFF_save_fm DFF_W3201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J203));
DFF_save_fm DFF_W3202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J213));
DFF_save_fm DFF_W3203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J223));
DFF_save_fm DFF_W3204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J004));
DFF_save_fm DFF_W3205(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J014));
DFF_save_fm DFF_W3206(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J024));
DFF_save_fm DFF_W3207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J104));
DFF_save_fm DFF_W3208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J114));
DFF_save_fm DFF_W3209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J124));
DFF_save_fm DFF_W3210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J204));
DFF_save_fm DFF_W3211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J214));
DFF_save_fm DFF_W3212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J224));
DFF_save_fm DFF_W3213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J005));
DFF_save_fm DFF_W3214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J015));
DFF_save_fm DFF_W3215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J025));
DFF_save_fm DFF_W3216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J105));
DFF_save_fm DFF_W3217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J115));
DFF_save_fm DFF_W3218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J125));
DFF_save_fm DFF_W3219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J205));
DFF_save_fm DFF_W3220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J215));
DFF_save_fm DFF_W3221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J225));
DFF_save_fm DFF_W3222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J006));
DFF_save_fm DFF_W3223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J016));
DFF_save_fm DFF_W3224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J026));
DFF_save_fm DFF_W3225(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J106));
DFF_save_fm DFF_W3226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J116));
DFF_save_fm DFF_W3227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J126));
DFF_save_fm DFF_W3228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J206));
DFF_save_fm DFF_W3229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J216));
DFF_save_fm DFF_W3230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J226));
DFF_save_fm DFF_W3231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J007));
DFF_save_fm DFF_W3232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J017));
DFF_save_fm DFF_W3233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J027));
DFF_save_fm DFF_W3234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J107));
DFF_save_fm DFF_W3235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J117));
DFF_save_fm DFF_W3236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J127));
DFF_save_fm DFF_W3237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J207));
DFF_save_fm DFF_W3238(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J217));
DFF_save_fm DFF_W3239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J227));
DFF_save_fm DFF_W3240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J008));
DFF_save_fm DFF_W3241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J018));
DFF_save_fm DFF_W3242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J028));
DFF_save_fm DFF_W3243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J108));
DFF_save_fm DFF_W3244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J118));
DFF_save_fm DFF_W3245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J128));
DFF_save_fm DFF_W3246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J208));
DFF_save_fm DFF_W3247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J218));
DFF_save_fm DFF_W3248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J228));
DFF_save_fm DFF_W3249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J009));
DFF_save_fm DFF_W3250(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J019));
DFF_save_fm DFF_W3251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J029));
DFF_save_fm DFF_W3252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J109));
DFF_save_fm DFF_W3253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J119));
DFF_save_fm DFF_W3254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J129));
DFF_save_fm DFF_W3255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J209));
DFF_save_fm DFF_W3256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J219));
DFF_save_fm DFF_W3257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J229));
DFF_save_fm DFF_W3258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J00A));
DFF_save_fm DFF_W3259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J01A));
DFF_save_fm DFF_W3260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J02A));
DFF_save_fm DFF_W3261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J10A));
DFF_save_fm DFF_W3262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J11A));
DFF_save_fm DFF_W3263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J12A));
DFF_save_fm DFF_W3264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J20A));
DFF_save_fm DFF_W3265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J21A));
DFF_save_fm DFF_W3266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J22A));
DFF_save_fm DFF_W3267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J00B));
DFF_save_fm DFF_W3268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J01B));
DFF_save_fm DFF_W3269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J02B));
DFF_save_fm DFF_W3270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J10B));
DFF_save_fm DFF_W3271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J11B));
DFF_save_fm DFF_W3272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J12B));
DFF_save_fm DFF_W3273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J20B));
DFF_save_fm DFF_W3274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J21B));
DFF_save_fm DFF_W3275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J22B));
DFF_save_fm DFF_W3276(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J00C));
DFF_save_fm DFF_W3277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J01C));
DFF_save_fm DFF_W3278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J02C));
DFF_save_fm DFF_W3279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J10C));
DFF_save_fm DFF_W3280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J11C));
DFF_save_fm DFF_W3281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J12C));
DFF_save_fm DFF_W3282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J20C));
DFF_save_fm DFF_W3283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J21C));
DFF_save_fm DFF_W3284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J22C));
DFF_save_fm DFF_W3285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J00D));
DFF_save_fm DFF_W3286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J01D));
DFF_save_fm DFF_W3287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J02D));
DFF_save_fm DFF_W3288(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J10D));
DFF_save_fm DFF_W3289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J11D));
DFF_save_fm DFF_W3290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J12D));
DFF_save_fm DFF_W3291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J20D));
DFF_save_fm DFF_W3292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J21D));
DFF_save_fm DFF_W3293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J22D));
DFF_save_fm DFF_W3294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J00E));
DFF_save_fm DFF_W3295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J01E));
DFF_save_fm DFF_W3296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J02E));
DFF_save_fm DFF_W3297(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J10E));
DFF_save_fm DFF_W3298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J11E));
DFF_save_fm DFF_W3299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J12E));
DFF_save_fm DFF_W3300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J20E));
DFF_save_fm DFF_W3301(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J21E));
DFF_save_fm DFF_W3302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J22E));
DFF_save_fm DFF_W3303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J00F));
DFF_save_fm DFF_W3304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J01F));
DFF_save_fm DFF_W3305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J02F));
DFF_save_fm DFF_W3306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J10F));
DFF_save_fm DFF_W3307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J11F));
DFF_save_fm DFF_W3308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J12F));
DFF_save_fm DFF_W3309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J20F));
DFF_save_fm DFF_W3310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1J21F));
DFF_save_fm DFF_W3311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1J22F));
DFF_save_fm DFF_W3312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K000));
DFF_save_fm DFF_W3313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K010));
DFF_save_fm DFF_W3314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K020));
DFF_save_fm DFF_W3315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K100));
DFF_save_fm DFF_W3316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K110));
DFF_save_fm DFF_W3317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K120));
DFF_save_fm DFF_W3318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K200));
DFF_save_fm DFF_W3319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K210));
DFF_save_fm DFF_W3320(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K220));
DFF_save_fm DFF_W3321(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K001));
DFF_save_fm DFF_W3322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K011));
DFF_save_fm DFF_W3323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K021));
DFF_save_fm DFF_W3324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K101));
DFF_save_fm DFF_W3325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K111));
DFF_save_fm DFF_W3326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K121));
DFF_save_fm DFF_W3327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K201));
DFF_save_fm DFF_W3328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K211));
DFF_save_fm DFF_W3329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K221));
DFF_save_fm DFF_W3330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K002));
DFF_save_fm DFF_W3331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K012));
DFF_save_fm DFF_W3332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K022));
DFF_save_fm DFF_W3333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K102));
DFF_save_fm DFF_W3334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K112));
DFF_save_fm DFF_W3335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K122));
DFF_save_fm DFF_W3336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K202));
DFF_save_fm DFF_W3337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K212));
DFF_save_fm DFF_W3338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K222));
DFF_save_fm DFF_W3339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K003));
DFF_save_fm DFF_W3340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K013));
DFF_save_fm DFF_W3341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K023));
DFF_save_fm DFF_W3342(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K103));
DFF_save_fm DFF_W3343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K113));
DFF_save_fm DFF_W3344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K123));
DFF_save_fm DFF_W3345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K203));
DFF_save_fm DFF_W3346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K213));
DFF_save_fm DFF_W3347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K223));
DFF_save_fm DFF_W3348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K004));
DFF_save_fm DFF_W3349(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K014));
DFF_save_fm DFF_W3350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K024));
DFF_save_fm DFF_W3351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K104));
DFF_save_fm DFF_W3352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K114));
DFF_save_fm DFF_W3353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K124));
DFF_save_fm DFF_W3354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K204));
DFF_save_fm DFF_W3355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K214));
DFF_save_fm DFF_W3356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K224));
DFF_save_fm DFF_W3357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K005));
DFF_save_fm DFF_W3358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K015));
DFF_save_fm DFF_W3359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K025));
DFF_save_fm DFF_W3360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K105));
DFF_save_fm DFF_W3361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K115));
DFF_save_fm DFF_W3362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K125));
DFF_save_fm DFF_W3363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K205));
DFF_save_fm DFF_W3364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K215));
DFF_save_fm DFF_W3365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K225));
DFF_save_fm DFF_W3366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K006));
DFF_save_fm DFF_W3367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K016));
DFF_save_fm DFF_W3368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K026));
DFF_save_fm DFF_W3369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K106));
DFF_save_fm DFF_W3370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K116));
DFF_save_fm DFF_W3371(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K126));
DFF_save_fm DFF_W3372(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K206));
DFF_save_fm DFF_W3373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K216));
DFF_save_fm DFF_W3374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K226));
DFF_save_fm DFF_W3375(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K007));
DFF_save_fm DFF_W3376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K017));
DFF_save_fm DFF_W3377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K027));
DFF_save_fm DFF_W3378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K107));
DFF_save_fm DFF_W3379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K117));
DFF_save_fm DFF_W3380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K127));
DFF_save_fm DFF_W3381(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K207));
DFF_save_fm DFF_W3382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K217));
DFF_save_fm DFF_W3383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K227));
DFF_save_fm DFF_W3384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K008));
DFF_save_fm DFF_W3385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K018));
DFF_save_fm DFF_W3386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K028));
DFF_save_fm DFF_W3387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K108));
DFF_save_fm DFF_W3388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K118));
DFF_save_fm DFF_W3389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K128));
DFF_save_fm DFF_W3390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K208));
DFF_save_fm DFF_W3391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K218));
DFF_save_fm DFF_W3392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K228));
DFF_save_fm DFF_W3393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K009));
DFF_save_fm DFF_W3394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K019));
DFF_save_fm DFF_W3395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K029));
DFF_save_fm DFF_W3396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K109));
DFF_save_fm DFF_W3397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K119));
DFF_save_fm DFF_W3398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K129));
DFF_save_fm DFF_W3399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K209));
DFF_save_fm DFF_W3400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K219));
DFF_save_fm DFF_W3401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K229));
DFF_save_fm DFF_W3402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K00A));
DFF_save_fm DFF_W3403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K01A));
DFF_save_fm DFF_W3404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K02A));
DFF_save_fm DFF_W3405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K10A));
DFF_save_fm DFF_W3406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K11A));
DFF_save_fm DFF_W3407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K12A));
DFF_save_fm DFF_W3408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K20A));
DFF_save_fm DFF_W3409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K21A));
DFF_save_fm DFF_W3410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K22A));
DFF_save_fm DFF_W3411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K00B));
DFF_save_fm DFF_W3412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K01B));
DFF_save_fm DFF_W3413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K02B));
DFF_save_fm DFF_W3414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K10B));
DFF_save_fm DFF_W3415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K11B));
DFF_save_fm DFF_W3416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K12B));
DFF_save_fm DFF_W3417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K20B));
DFF_save_fm DFF_W3418(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K21B));
DFF_save_fm DFF_W3419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K22B));
DFF_save_fm DFF_W3420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K00C));
DFF_save_fm DFF_W3421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K01C));
DFF_save_fm DFF_W3422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K02C));
DFF_save_fm DFF_W3423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K10C));
DFF_save_fm DFF_W3424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K11C));
DFF_save_fm DFF_W3425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K12C));
DFF_save_fm DFF_W3426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K20C));
DFF_save_fm DFF_W3427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K21C));
DFF_save_fm DFF_W3428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K22C));
DFF_save_fm DFF_W3429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K00D));
DFF_save_fm DFF_W3430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K01D));
DFF_save_fm DFF_W3431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K02D));
DFF_save_fm DFF_W3432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K10D));
DFF_save_fm DFF_W3433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K11D));
DFF_save_fm DFF_W3434(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K12D));
DFF_save_fm DFF_W3435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K20D));
DFF_save_fm DFF_W3436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K21D));
DFF_save_fm DFF_W3437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K22D));
DFF_save_fm DFF_W3438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K00E));
DFF_save_fm DFF_W3439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K01E));
DFF_save_fm DFF_W3440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K02E));
DFF_save_fm DFF_W3441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K10E));
DFF_save_fm DFF_W3442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K11E));
DFF_save_fm DFF_W3443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K12E));
DFF_save_fm DFF_W3444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K20E));
DFF_save_fm DFF_W3445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K21E));
DFF_save_fm DFF_W3446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K22E));
DFF_save_fm DFF_W3447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K00F));
DFF_save_fm DFF_W3448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K01F));
DFF_save_fm DFF_W3449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K02F));
DFF_save_fm DFF_W3450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K10F));
DFF_save_fm DFF_W3451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K11F));
DFF_save_fm DFF_W3452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K12F));
DFF_save_fm DFF_W3453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K20F));
DFF_save_fm DFF_W3454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1K21F));
DFF_save_fm DFF_W3455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1K22F));
DFF_save_fm DFF_W3456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L000));
DFF_save_fm DFF_W3457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L010));
DFF_save_fm DFF_W3458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L020));
DFF_save_fm DFF_W3459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L100));
DFF_save_fm DFF_W3460(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L110));
DFF_save_fm DFF_W3461(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L120));
DFF_save_fm DFF_W3462(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L200));
DFF_save_fm DFF_W3463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L210));
DFF_save_fm DFF_W3464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L220));
DFF_save_fm DFF_W3465(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L001));
DFF_save_fm DFF_W3466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L011));
DFF_save_fm DFF_W3467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L021));
DFF_save_fm DFF_W3468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L101));
DFF_save_fm DFF_W3469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L111));
DFF_save_fm DFF_W3470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L121));
DFF_save_fm DFF_W3471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L201));
DFF_save_fm DFF_W3472(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L211));
DFF_save_fm DFF_W3473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L221));
DFF_save_fm DFF_W3474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L002));
DFF_save_fm DFF_W3475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L012));
DFF_save_fm DFF_W3476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L022));
DFF_save_fm DFF_W3477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L102));
DFF_save_fm DFF_W3478(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L112));
DFF_save_fm DFF_W3479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L122));
DFF_save_fm DFF_W3480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L202));
DFF_save_fm DFF_W3481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L212));
DFF_save_fm DFF_W3482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L222));
DFF_save_fm DFF_W3483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L003));
DFF_save_fm DFF_W3484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L013));
DFF_save_fm DFF_W3485(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L023));
DFF_save_fm DFF_W3486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L103));
DFF_save_fm DFF_W3487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L113));
DFF_save_fm DFF_W3488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L123));
DFF_save_fm DFF_W3489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L203));
DFF_save_fm DFF_W3490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L213));
DFF_save_fm DFF_W3491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L223));
DFF_save_fm DFF_W3492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L004));
DFF_save_fm DFF_W3493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L014));
DFF_save_fm DFF_W3494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L024));
DFF_save_fm DFF_W3495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L104));
DFF_save_fm DFF_W3496(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L114));
DFF_save_fm DFF_W3497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L124));
DFF_save_fm DFF_W3498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L204));
DFF_save_fm DFF_W3499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L214));
DFF_save_fm DFF_W3500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L224));
DFF_save_fm DFF_W3501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L005));
DFF_save_fm DFF_W3502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L015));
DFF_save_fm DFF_W3503(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L025));
DFF_save_fm DFF_W3504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L105));
DFF_save_fm DFF_W3505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L115));
DFF_save_fm DFF_W3506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L125));
DFF_save_fm DFF_W3507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L205));
DFF_save_fm DFF_W3508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L215));
DFF_save_fm DFF_W3509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L225));
DFF_save_fm DFF_W3510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L006));
DFF_save_fm DFF_W3511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L016));
DFF_save_fm DFF_W3512(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L026));
DFF_save_fm DFF_W3513(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L106));
DFF_save_fm DFF_W3514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L116));
DFF_save_fm DFF_W3515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L126));
DFF_save_fm DFF_W3516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L206));
DFF_save_fm DFF_W3517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L216));
DFF_save_fm DFF_W3518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L226));
DFF_save_fm DFF_W3519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L007));
DFF_save_fm DFF_W3520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L017));
DFF_save_fm DFF_W3521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L027));
DFF_save_fm DFF_W3522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L107));
DFF_save_fm DFF_W3523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L117));
DFF_save_fm DFF_W3524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L127));
DFF_save_fm DFF_W3525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L207));
DFF_save_fm DFF_W3526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L217));
DFF_save_fm DFF_W3527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L227));
DFF_save_fm DFF_W3528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L008));
DFF_save_fm DFF_W3529(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L018));
DFF_save_fm DFF_W3530(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L028));
DFF_save_fm DFF_W3531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L108));
DFF_save_fm DFF_W3532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L118));
DFF_save_fm DFF_W3533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L128));
DFF_save_fm DFF_W3534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L208));
DFF_save_fm DFF_W3535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L218));
DFF_save_fm DFF_W3536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L228));
DFF_save_fm DFF_W3537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L009));
DFF_save_fm DFF_W3538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L019));
DFF_save_fm DFF_W3539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L029));
DFF_save_fm DFF_W3540(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L109));
DFF_save_fm DFF_W3541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L119));
DFF_save_fm DFF_W3542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L129));
DFF_save_fm DFF_W3543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L209));
DFF_save_fm DFF_W3544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L219));
DFF_save_fm DFF_W3545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L229));
DFF_save_fm DFF_W3546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L00A));
DFF_save_fm DFF_W3547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L01A));
DFF_save_fm DFF_W3548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L02A));
DFF_save_fm DFF_W3549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L10A));
DFF_save_fm DFF_W3550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L11A));
DFF_save_fm DFF_W3551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L12A));
DFF_save_fm DFF_W3552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L20A));
DFF_save_fm DFF_W3553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L21A));
DFF_save_fm DFF_W3554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L22A));
DFF_save_fm DFF_W3555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L00B));
DFF_save_fm DFF_W3556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L01B));
DFF_save_fm DFF_W3557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L02B));
DFF_save_fm DFF_W3558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L10B));
DFF_save_fm DFF_W3559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L11B));
DFF_save_fm DFF_W3560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L12B));
DFF_save_fm DFF_W3561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L20B));
DFF_save_fm DFF_W3562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L21B));
DFF_save_fm DFF_W3563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L22B));
DFF_save_fm DFF_W3564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L00C));
DFF_save_fm DFF_W3565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L01C));
DFF_save_fm DFF_W3566(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L02C));
DFF_save_fm DFF_W3567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L10C));
DFF_save_fm DFF_W3568(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L11C));
DFF_save_fm DFF_W3569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L12C));
DFF_save_fm DFF_W3570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L20C));
DFF_save_fm DFF_W3571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L21C));
DFF_save_fm DFF_W3572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L22C));
DFF_save_fm DFF_W3573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L00D));
DFF_save_fm DFF_W3574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L01D));
DFF_save_fm DFF_W3575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L02D));
DFF_save_fm DFF_W3576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L10D));
DFF_save_fm DFF_W3577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L11D));
DFF_save_fm DFF_W3578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L12D));
DFF_save_fm DFF_W3579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L20D));
DFF_save_fm DFF_W3580(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L21D));
DFF_save_fm DFF_W3581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L22D));
DFF_save_fm DFF_W3582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L00E));
DFF_save_fm DFF_W3583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L01E));
DFF_save_fm DFF_W3584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L02E));
DFF_save_fm DFF_W3585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L10E));
DFF_save_fm DFF_W3586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L11E));
DFF_save_fm DFF_W3587(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L12E));
DFF_save_fm DFF_W3588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L20E));
DFF_save_fm DFF_W3589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L21E));
DFF_save_fm DFF_W3590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L22E));
DFF_save_fm DFF_W3591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L00F));
DFF_save_fm DFF_W3592(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L01F));
DFF_save_fm DFF_W3593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L02F));
DFF_save_fm DFF_W3594(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L10F));
DFF_save_fm DFF_W3595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L11F));
DFF_save_fm DFF_W3596(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L12F));
DFF_save_fm DFF_W3597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L20F));
DFF_save_fm DFF_W3598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1L21F));
DFF_save_fm DFF_W3599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1L22F));
DFF_save_fm DFF_W3600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M000));
DFF_save_fm DFF_W3601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M010));
DFF_save_fm DFF_W3602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M020));
DFF_save_fm DFF_W3603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M100));
DFF_save_fm DFF_W3604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M110));
DFF_save_fm DFF_W3605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M120));
DFF_save_fm DFF_W3606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M200));
DFF_save_fm DFF_W3607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M210));
DFF_save_fm DFF_W3608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M220));
DFF_save_fm DFF_W3609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M001));
DFF_save_fm DFF_W3610(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M011));
DFF_save_fm DFF_W3611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M021));
DFF_save_fm DFF_W3612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M101));
DFF_save_fm DFF_W3613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M111));
DFF_save_fm DFF_W3614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M121));
DFF_save_fm DFF_W3615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M201));
DFF_save_fm DFF_W3616(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M211));
DFF_save_fm DFF_W3617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M221));
DFF_save_fm DFF_W3618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M002));
DFF_save_fm DFF_W3619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M012));
DFF_save_fm DFF_W3620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M022));
DFF_save_fm DFF_W3621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M102));
DFF_save_fm DFF_W3622(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M112));
DFF_save_fm DFF_W3623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M122));
DFF_save_fm DFF_W3624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M202));
DFF_save_fm DFF_W3625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M212));
DFF_save_fm DFF_W3626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M222));
DFF_save_fm DFF_W3627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M003));
DFF_save_fm DFF_W3628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M013));
DFF_save_fm DFF_W3629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M023));
DFF_save_fm DFF_W3630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M103));
DFF_save_fm DFF_W3631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M113));
DFF_save_fm DFF_W3632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M123));
DFF_save_fm DFF_W3633(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M203));
DFF_save_fm DFF_W3634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M213));
DFF_save_fm DFF_W3635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M223));
DFF_save_fm DFF_W3636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M004));
DFF_save_fm DFF_W3637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M014));
DFF_save_fm DFF_W3638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M024));
DFF_save_fm DFF_W3639(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M104));
DFF_save_fm DFF_W3640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M114));
DFF_save_fm DFF_W3641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M124));
DFF_save_fm DFF_W3642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M204));
DFF_save_fm DFF_W3643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M214));
DFF_save_fm DFF_W3644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M224));
DFF_save_fm DFF_W3645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M005));
DFF_save_fm DFF_W3646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M015));
DFF_save_fm DFF_W3647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M025));
DFF_save_fm DFF_W3648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M105));
DFF_save_fm DFF_W3649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M115));
DFF_save_fm DFF_W3650(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M125));
DFF_save_fm DFF_W3651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M205));
DFF_save_fm DFF_W3652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M215));
DFF_save_fm DFF_W3653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M225));
DFF_save_fm DFF_W3654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M006));
DFF_save_fm DFF_W3655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M016));
DFF_save_fm DFF_W3656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M026));
DFF_save_fm DFF_W3657(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M106));
DFF_save_fm DFF_W3658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M116));
DFF_save_fm DFF_W3659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M126));
DFF_save_fm DFF_W3660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M206));
DFF_save_fm DFF_W3661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M216));
DFF_save_fm DFF_W3662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M226));
DFF_save_fm DFF_W3663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M007));
DFF_save_fm DFF_W3664(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M017));
DFF_save_fm DFF_W3665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M027));
DFF_save_fm DFF_W3666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M107));
DFF_save_fm DFF_W3667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M117));
DFF_save_fm DFF_W3668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M127));
DFF_save_fm DFF_W3669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M207));
DFF_save_fm DFF_W3670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M217));
DFF_save_fm DFF_W3671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M227));
DFF_save_fm DFF_W3672(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M008));
DFF_save_fm DFF_W3673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M018));
DFF_save_fm DFF_W3674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M028));
DFF_save_fm DFF_W3675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M108));
DFF_save_fm DFF_W3676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M118));
DFF_save_fm DFF_W3677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M128));
DFF_save_fm DFF_W3678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M208));
DFF_save_fm DFF_W3679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M218));
DFF_save_fm DFF_W3680(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M228));
DFF_save_fm DFF_W3681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M009));
DFF_save_fm DFF_W3682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M019));
DFF_save_fm DFF_W3683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M029));
DFF_save_fm DFF_W3684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M109));
DFF_save_fm DFF_W3685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M119));
DFF_save_fm DFF_W3686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M129));
DFF_save_fm DFF_W3687(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M209));
DFF_save_fm DFF_W3688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M219));
DFF_save_fm DFF_W3689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M229));
DFF_save_fm DFF_W3690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M00A));
DFF_save_fm DFF_W3691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M01A));
DFF_save_fm DFF_W3692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M02A));
DFF_save_fm DFF_W3693(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M10A));
DFF_save_fm DFF_W3694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M11A));
DFF_save_fm DFF_W3695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M12A));
DFF_save_fm DFF_W3696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M20A));
DFF_save_fm DFF_W3697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M21A));
DFF_save_fm DFF_W3698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M22A));
DFF_save_fm DFF_W3699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M00B));
DFF_save_fm DFF_W3700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M01B));
DFF_save_fm DFF_W3701(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M02B));
DFF_save_fm DFF_W3702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M10B));
DFF_save_fm DFF_W3703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M11B));
DFF_save_fm DFF_W3704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M12B));
DFF_save_fm DFF_W3705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M20B));
DFF_save_fm DFF_W3706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M21B));
DFF_save_fm DFF_W3707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M22B));
DFF_save_fm DFF_W3708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M00C));
DFF_save_fm DFF_W3709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M01C));
DFF_save_fm DFF_W3710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M02C));
DFF_save_fm DFF_W3711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M10C));
DFF_save_fm DFF_W3712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M11C));
DFF_save_fm DFF_W3713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M12C));
DFF_save_fm DFF_W3714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M20C));
DFF_save_fm DFF_W3715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M21C));
DFF_save_fm DFF_W3716(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M22C));
DFF_save_fm DFF_W3717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M00D));
DFF_save_fm DFF_W3718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M01D));
DFF_save_fm DFF_W3719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M02D));
DFF_save_fm DFF_W3720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M10D));
DFF_save_fm DFF_W3721(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M11D));
DFF_save_fm DFF_W3722(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M12D));
DFF_save_fm DFF_W3723(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M20D));
DFF_save_fm DFF_W3724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M21D));
DFF_save_fm DFF_W3725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M22D));
DFF_save_fm DFF_W3726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M00E));
DFF_save_fm DFF_W3727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M01E));
DFF_save_fm DFF_W3728(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M02E));
DFF_save_fm DFF_W3729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M10E));
DFF_save_fm DFF_W3730(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M11E));
DFF_save_fm DFF_W3731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M12E));
DFF_save_fm DFF_W3732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M20E));
DFF_save_fm DFF_W3733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M21E));
DFF_save_fm DFF_W3734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M22E));
DFF_save_fm DFF_W3735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M00F));
DFF_save_fm DFF_W3736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M01F));
DFF_save_fm DFF_W3737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M02F));
DFF_save_fm DFF_W3738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M10F));
DFF_save_fm DFF_W3739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M11F));
DFF_save_fm DFF_W3740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M12F));
DFF_save_fm DFF_W3741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1M20F));
DFF_save_fm DFF_W3742(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M21F));
DFF_save_fm DFF_W3743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1M22F));
ninexnine_unit ninexnine_unit_1200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10000)
);

ninexnine_unit ninexnine_unit_1201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11000)
);

ninexnine_unit ninexnine_unit_1202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12000)
);

ninexnine_unit ninexnine_unit_1203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13000)
);

ninexnine_unit ninexnine_unit_1204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14000)
);

ninexnine_unit ninexnine_unit_1205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15000)
);

ninexnine_unit ninexnine_unit_1206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16000)
);

ninexnine_unit ninexnine_unit_1207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17000)
);

ninexnine_unit ninexnine_unit_1208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18000)
);

ninexnine_unit ninexnine_unit_1209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19000)
);

ninexnine_unit ninexnine_unit_1210(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A000)
);

ninexnine_unit ninexnine_unit_1211(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B000)
);

ninexnine_unit ninexnine_unit_1212(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C000)
);

ninexnine_unit ninexnine_unit_1213(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D000)
);

ninexnine_unit ninexnine_unit_1214(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E000)
);

ninexnine_unit ninexnine_unit_1215(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F000)
);

assign C1000=c10000+c11000+c12000+c13000+c14000+c15000+c16000+c17000+c18000+c19000+c1A000+c1B000+c1C000+c1D000+c1E000+c1F000;
assign A1000=(C1000>=0)?1:0;

assign P2000=A1000;

ninexnine_unit ninexnine_unit_1216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10010)
);

ninexnine_unit ninexnine_unit_1217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11010)
);

ninexnine_unit ninexnine_unit_1218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12010)
);

ninexnine_unit ninexnine_unit_1219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13010)
);

ninexnine_unit ninexnine_unit_1220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14010)
);

ninexnine_unit ninexnine_unit_1221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15010)
);

ninexnine_unit ninexnine_unit_1222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16010)
);

ninexnine_unit ninexnine_unit_1223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17010)
);

ninexnine_unit ninexnine_unit_1224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18010)
);

ninexnine_unit ninexnine_unit_1225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19010)
);

ninexnine_unit ninexnine_unit_1226(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A010)
);

ninexnine_unit ninexnine_unit_1227(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B010)
);

ninexnine_unit ninexnine_unit_1228(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C010)
);

ninexnine_unit ninexnine_unit_1229(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D010)
);

ninexnine_unit ninexnine_unit_1230(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E010)
);

ninexnine_unit ninexnine_unit_1231(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F010)
);

assign C1010=c10010+c11010+c12010+c13010+c14010+c15010+c16010+c17010+c18010+c19010+c1A010+c1B010+c1C010+c1D010+c1E010+c1F010;
assign A1010=(C1010>=0)?1:0;

assign P2010=A1010;

ninexnine_unit ninexnine_unit_1232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10020)
);

ninexnine_unit ninexnine_unit_1233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11020)
);

ninexnine_unit ninexnine_unit_1234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12020)
);

ninexnine_unit ninexnine_unit_1235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13020)
);

ninexnine_unit ninexnine_unit_1236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14020)
);

ninexnine_unit ninexnine_unit_1237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15020)
);

ninexnine_unit ninexnine_unit_1238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16020)
);

ninexnine_unit ninexnine_unit_1239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17020)
);

ninexnine_unit ninexnine_unit_1240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18020)
);

ninexnine_unit ninexnine_unit_1241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19020)
);

ninexnine_unit ninexnine_unit_1242(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A020)
);

ninexnine_unit ninexnine_unit_1243(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B020)
);

ninexnine_unit ninexnine_unit_1244(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C020)
);

ninexnine_unit ninexnine_unit_1245(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D020)
);

ninexnine_unit ninexnine_unit_1246(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E020)
);

ninexnine_unit ninexnine_unit_1247(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F020)
);

assign C1020=c10020+c11020+c12020+c13020+c14020+c15020+c16020+c17020+c18020+c19020+c1A020+c1B020+c1C020+c1D020+c1E020+c1F020;
assign A1020=(C1020>=0)?1:0;

assign P2020=A1020;

ninexnine_unit ninexnine_unit_1248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10100)
);

ninexnine_unit ninexnine_unit_1249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11100)
);

ninexnine_unit ninexnine_unit_1250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12100)
);

ninexnine_unit ninexnine_unit_1251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13100)
);

ninexnine_unit ninexnine_unit_1252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14100)
);

ninexnine_unit ninexnine_unit_1253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15100)
);

ninexnine_unit ninexnine_unit_1254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16100)
);

ninexnine_unit ninexnine_unit_1255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17100)
);

ninexnine_unit ninexnine_unit_1256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18100)
);

ninexnine_unit ninexnine_unit_1257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19100)
);

ninexnine_unit ninexnine_unit_1258(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A100)
);

ninexnine_unit ninexnine_unit_1259(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B100)
);

ninexnine_unit ninexnine_unit_1260(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C100)
);

ninexnine_unit ninexnine_unit_1261(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D100)
);

ninexnine_unit ninexnine_unit_1262(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E100)
);

ninexnine_unit ninexnine_unit_1263(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F100)
);

assign C1100=c10100+c11100+c12100+c13100+c14100+c15100+c16100+c17100+c18100+c19100+c1A100+c1B100+c1C100+c1D100+c1E100+c1F100;
assign A1100=(C1100>=0)?1:0;

assign P2100=A1100;

ninexnine_unit ninexnine_unit_1264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10110)
);

ninexnine_unit ninexnine_unit_1265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11110)
);

ninexnine_unit ninexnine_unit_1266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12110)
);

ninexnine_unit ninexnine_unit_1267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13110)
);

ninexnine_unit ninexnine_unit_1268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14110)
);

ninexnine_unit ninexnine_unit_1269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15110)
);

ninexnine_unit ninexnine_unit_1270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16110)
);

ninexnine_unit ninexnine_unit_1271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17110)
);

ninexnine_unit ninexnine_unit_1272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18110)
);

ninexnine_unit ninexnine_unit_1273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19110)
);

ninexnine_unit ninexnine_unit_1274(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A110)
);

ninexnine_unit ninexnine_unit_1275(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B110)
);

ninexnine_unit ninexnine_unit_1276(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C110)
);

ninexnine_unit ninexnine_unit_1277(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D110)
);

ninexnine_unit ninexnine_unit_1278(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E110)
);

ninexnine_unit ninexnine_unit_1279(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F110)
);

assign C1110=c10110+c11110+c12110+c13110+c14110+c15110+c16110+c17110+c18110+c19110+c1A110+c1B110+c1C110+c1D110+c1E110+c1F110;
assign A1110=(C1110>=0)?1:0;

assign P2110=A1110;

ninexnine_unit ninexnine_unit_1280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10120)
);

ninexnine_unit ninexnine_unit_1281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11120)
);

ninexnine_unit ninexnine_unit_1282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12120)
);

ninexnine_unit ninexnine_unit_1283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13120)
);

ninexnine_unit ninexnine_unit_1284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14120)
);

ninexnine_unit ninexnine_unit_1285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15120)
);

ninexnine_unit ninexnine_unit_1286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16120)
);

ninexnine_unit ninexnine_unit_1287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17120)
);

ninexnine_unit ninexnine_unit_1288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18120)
);

ninexnine_unit ninexnine_unit_1289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19120)
);

ninexnine_unit ninexnine_unit_1290(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A120)
);

ninexnine_unit ninexnine_unit_1291(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B120)
);

ninexnine_unit ninexnine_unit_1292(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C120)
);

ninexnine_unit ninexnine_unit_1293(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D120)
);

ninexnine_unit ninexnine_unit_1294(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E120)
);

ninexnine_unit ninexnine_unit_1295(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F120)
);

assign C1120=c10120+c11120+c12120+c13120+c14120+c15120+c16120+c17120+c18120+c19120+c1A120+c1B120+c1C120+c1D120+c1E120+c1F120;
assign A1120=(C1120>=0)?1:0;

assign P2120=A1120;

ninexnine_unit ninexnine_unit_1296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10200)
);

ninexnine_unit ninexnine_unit_1297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11200)
);

ninexnine_unit ninexnine_unit_1298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12200)
);

ninexnine_unit ninexnine_unit_1299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13200)
);

ninexnine_unit ninexnine_unit_1300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14200)
);

ninexnine_unit ninexnine_unit_1301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15200)
);

ninexnine_unit ninexnine_unit_1302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16200)
);

ninexnine_unit ninexnine_unit_1303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17200)
);

ninexnine_unit ninexnine_unit_1304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18200)
);

ninexnine_unit ninexnine_unit_1305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19200)
);

ninexnine_unit ninexnine_unit_1306(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A200)
);

ninexnine_unit ninexnine_unit_1307(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B200)
);

ninexnine_unit ninexnine_unit_1308(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C200)
);

ninexnine_unit ninexnine_unit_1309(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D200)
);

ninexnine_unit ninexnine_unit_1310(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E200)
);

ninexnine_unit ninexnine_unit_1311(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F200)
);

assign C1200=c10200+c11200+c12200+c13200+c14200+c15200+c16200+c17200+c18200+c19200+c1A200+c1B200+c1C200+c1D200+c1E200+c1F200;
assign A1200=(C1200>=0)?1:0;

assign P2200=A1200;

ninexnine_unit ninexnine_unit_1312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10210)
);

ninexnine_unit ninexnine_unit_1313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11210)
);

ninexnine_unit ninexnine_unit_1314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12210)
);

ninexnine_unit ninexnine_unit_1315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13210)
);

ninexnine_unit ninexnine_unit_1316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14210)
);

ninexnine_unit ninexnine_unit_1317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15210)
);

ninexnine_unit ninexnine_unit_1318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16210)
);

ninexnine_unit ninexnine_unit_1319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17210)
);

ninexnine_unit ninexnine_unit_1320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18210)
);

ninexnine_unit ninexnine_unit_1321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19210)
);

ninexnine_unit ninexnine_unit_1322(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A210)
);

ninexnine_unit ninexnine_unit_1323(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B210)
);

ninexnine_unit ninexnine_unit_1324(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C210)
);

ninexnine_unit ninexnine_unit_1325(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D210)
);

ninexnine_unit ninexnine_unit_1326(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E210)
);

ninexnine_unit ninexnine_unit_1327(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F210)
);

assign C1210=c10210+c11210+c12210+c13210+c14210+c15210+c16210+c17210+c18210+c19210+c1A210+c1B210+c1C210+c1D210+c1E210+c1F210;
assign A1210=(C1210>=0)?1:0;

assign P2210=A1210;

ninexnine_unit ninexnine_unit_1328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10220)
);

ninexnine_unit ninexnine_unit_1329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11220)
);

ninexnine_unit ninexnine_unit_1330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12220)
);

ninexnine_unit ninexnine_unit_1331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13220)
);

ninexnine_unit ninexnine_unit_1332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W10004),
				.b1(W10014),
				.b2(W10024),
				.b3(W10104),
				.b4(W10114),
				.b5(W10124),
				.b6(W10204),
				.b7(W10214),
				.b8(W10224),
				.c(c14220)
);

ninexnine_unit ninexnine_unit_1333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W10005),
				.b1(W10015),
				.b2(W10025),
				.b3(W10105),
				.b4(W10115),
				.b5(W10125),
				.b6(W10205),
				.b7(W10215),
				.b8(W10225),
				.c(c15220)
);

ninexnine_unit ninexnine_unit_1334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W10006),
				.b1(W10016),
				.b2(W10026),
				.b3(W10106),
				.b4(W10116),
				.b5(W10126),
				.b6(W10206),
				.b7(W10216),
				.b8(W10226),
				.c(c16220)
);

ninexnine_unit ninexnine_unit_1335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W10007),
				.b1(W10017),
				.b2(W10027),
				.b3(W10107),
				.b4(W10117),
				.b5(W10127),
				.b6(W10207),
				.b7(W10217),
				.b8(W10227),
				.c(c17220)
);

ninexnine_unit ninexnine_unit_1336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W10008),
				.b1(W10018),
				.b2(W10028),
				.b3(W10108),
				.b4(W10118),
				.b5(W10128),
				.b6(W10208),
				.b7(W10218),
				.b8(W10228),
				.c(c18220)
);

ninexnine_unit ninexnine_unit_1337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W10009),
				.b1(W10019),
				.b2(W10029),
				.b3(W10109),
				.b4(W10119),
				.b5(W10129),
				.b6(W10209),
				.b7(W10219),
				.b8(W10229),
				.c(c19220)
);

ninexnine_unit ninexnine_unit_1338(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1000A),
				.b1(W1001A),
				.b2(W1002A),
				.b3(W1010A),
				.b4(W1011A),
				.b5(W1012A),
				.b6(W1020A),
				.b7(W1021A),
				.b8(W1022A),
				.c(c1A220)
);

ninexnine_unit ninexnine_unit_1339(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1000B),
				.b1(W1001B),
				.b2(W1002B),
				.b3(W1010B),
				.b4(W1011B),
				.b5(W1012B),
				.b6(W1020B),
				.b7(W1021B),
				.b8(W1022B),
				.c(c1B220)
);

ninexnine_unit ninexnine_unit_1340(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1000C),
				.b1(W1001C),
				.b2(W1002C),
				.b3(W1010C),
				.b4(W1011C),
				.b5(W1012C),
				.b6(W1020C),
				.b7(W1021C),
				.b8(W1022C),
				.c(c1C220)
);

ninexnine_unit ninexnine_unit_1341(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1000D),
				.b1(W1001D),
				.b2(W1002D),
				.b3(W1010D),
				.b4(W1011D),
				.b5(W1012D),
				.b6(W1020D),
				.b7(W1021D),
				.b8(W1022D),
				.c(c1D220)
);

ninexnine_unit ninexnine_unit_1342(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1000E),
				.b1(W1001E),
				.b2(W1002E),
				.b3(W1010E),
				.b4(W1011E),
				.b5(W1012E),
				.b6(W1020E),
				.b7(W1021E),
				.b8(W1022E),
				.c(c1E220)
);

ninexnine_unit ninexnine_unit_1343(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1000F),
				.b1(W1001F),
				.b2(W1002F),
				.b3(W1010F),
				.b4(W1011F),
				.b5(W1012F),
				.b6(W1020F),
				.b7(W1021F),
				.b8(W1022F),
				.c(c1F220)
);

assign C1220=c10220+c11220+c12220+c13220+c14220+c15220+c16220+c17220+c18220+c19220+c1A220+c1B220+c1C220+c1D220+c1E220+c1F220;
assign A1220=(C1220>=0)?1:0;

assign P2220=A1220;

ninexnine_unit ninexnine_unit_1344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10001)
);

ninexnine_unit ninexnine_unit_1345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11001)
);

ninexnine_unit ninexnine_unit_1346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12001)
);

ninexnine_unit ninexnine_unit_1347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13001)
);

ninexnine_unit ninexnine_unit_1348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14001)
);

ninexnine_unit ninexnine_unit_1349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15001)
);

ninexnine_unit ninexnine_unit_1350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16001)
);

ninexnine_unit ninexnine_unit_1351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17001)
);

ninexnine_unit ninexnine_unit_1352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18001)
);

ninexnine_unit ninexnine_unit_1353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19001)
);

ninexnine_unit ninexnine_unit_1354(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A001)
);

ninexnine_unit ninexnine_unit_1355(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B001)
);

ninexnine_unit ninexnine_unit_1356(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C001)
);

ninexnine_unit ninexnine_unit_1357(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D001)
);

ninexnine_unit ninexnine_unit_1358(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E001)
);

ninexnine_unit ninexnine_unit_1359(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F001)
);

assign C1001=c10001+c11001+c12001+c13001+c14001+c15001+c16001+c17001+c18001+c19001+c1A001+c1B001+c1C001+c1D001+c1E001+c1F001;
assign A1001=(C1001>=0)?1:0;

assign P2001=A1001;

ninexnine_unit ninexnine_unit_1360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10011)
);

ninexnine_unit ninexnine_unit_1361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11011)
);

ninexnine_unit ninexnine_unit_1362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12011)
);

ninexnine_unit ninexnine_unit_1363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13011)
);

ninexnine_unit ninexnine_unit_1364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14011)
);

ninexnine_unit ninexnine_unit_1365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15011)
);

ninexnine_unit ninexnine_unit_1366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16011)
);

ninexnine_unit ninexnine_unit_1367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17011)
);

ninexnine_unit ninexnine_unit_1368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18011)
);

ninexnine_unit ninexnine_unit_1369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19011)
);

ninexnine_unit ninexnine_unit_1370(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A011)
);

ninexnine_unit ninexnine_unit_1371(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B011)
);

ninexnine_unit ninexnine_unit_1372(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C011)
);

ninexnine_unit ninexnine_unit_1373(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D011)
);

ninexnine_unit ninexnine_unit_1374(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E011)
);

ninexnine_unit ninexnine_unit_1375(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F011)
);

assign C1011=c10011+c11011+c12011+c13011+c14011+c15011+c16011+c17011+c18011+c19011+c1A011+c1B011+c1C011+c1D011+c1E011+c1F011;
assign A1011=(C1011>=0)?1:0;

assign P2011=A1011;

ninexnine_unit ninexnine_unit_1376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10021)
);

ninexnine_unit ninexnine_unit_1377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11021)
);

ninexnine_unit ninexnine_unit_1378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12021)
);

ninexnine_unit ninexnine_unit_1379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13021)
);

ninexnine_unit ninexnine_unit_1380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14021)
);

ninexnine_unit ninexnine_unit_1381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15021)
);

ninexnine_unit ninexnine_unit_1382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16021)
);

ninexnine_unit ninexnine_unit_1383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17021)
);

ninexnine_unit ninexnine_unit_1384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18021)
);

ninexnine_unit ninexnine_unit_1385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19021)
);

ninexnine_unit ninexnine_unit_1386(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A021)
);

ninexnine_unit ninexnine_unit_1387(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B021)
);

ninexnine_unit ninexnine_unit_1388(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C021)
);

ninexnine_unit ninexnine_unit_1389(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D021)
);

ninexnine_unit ninexnine_unit_1390(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E021)
);

ninexnine_unit ninexnine_unit_1391(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F021)
);

assign C1021=c10021+c11021+c12021+c13021+c14021+c15021+c16021+c17021+c18021+c19021+c1A021+c1B021+c1C021+c1D021+c1E021+c1F021;
assign A1021=(C1021>=0)?1:0;

assign P2021=A1021;

ninexnine_unit ninexnine_unit_1392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10101)
);

ninexnine_unit ninexnine_unit_1393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11101)
);

ninexnine_unit ninexnine_unit_1394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12101)
);

ninexnine_unit ninexnine_unit_1395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13101)
);

ninexnine_unit ninexnine_unit_1396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14101)
);

ninexnine_unit ninexnine_unit_1397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15101)
);

ninexnine_unit ninexnine_unit_1398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16101)
);

ninexnine_unit ninexnine_unit_1399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17101)
);

ninexnine_unit ninexnine_unit_1400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18101)
);

ninexnine_unit ninexnine_unit_1401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19101)
);

ninexnine_unit ninexnine_unit_1402(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A101)
);

ninexnine_unit ninexnine_unit_1403(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B101)
);

ninexnine_unit ninexnine_unit_1404(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C101)
);

ninexnine_unit ninexnine_unit_1405(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D101)
);

ninexnine_unit ninexnine_unit_1406(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E101)
);

ninexnine_unit ninexnine_unit_1407(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F101)
);

assign C1101=c10101+c11101+c12101+c13101+c14101+c15101+c16101+c17101+c18101+c19101+c1A101+c1B101+c1C101+c1D101+c1E101+c1F101;
assign A1101=(C1101>=0)?1:0;

assign P2101=A1101;

ninexnine_unit ninexnine_unit_1408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10111)
);

ninexnine_unit ninexnine_unit_1409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11111)
);

ninexnine_unit ninexnine_unit_1410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12111)
);

ninexnine_unit ninexnine_unit_1411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13111)
);

ninexnine_unit ninexnine_unit_1412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14111)
);

ninexnine_unit ninexnine_unit_1413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15111)
);

ninexnine_unit ninexnine_unit_1414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16111)
);

ninexnine_unit ninexnine_unit_1415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17111)
);

ninexnine_unit ninexnine_unit_1416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18111)
);

ninexnine_unit ninexnine_unit_1417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19111)
);

ninexnine_unit ninexnine_unit_1418(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A111)
);

ninexnine_unit ninexnine_unit_1419(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B111)
);

ninexnine_unit ninexnine_unit_1420(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C111)
);

ninexnine_unit ninexnine_unit_1421(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D111)
);

ninexnine_unit ninexnine_unit_1422(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E111)
);

ninexnine_unit ninexnine_unit_1423(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F111)
);

assign C1111=c10111+c11111+c12111+c13111+c14111+c15111+c16111+c17111+c18111+c19111+c1A111+c1B111+c1C111+c1D111+c1E111+c1F111;
assign A1111=(C1111>=0)?1:0;

assign P2111=A1111;

ninexnine_unit ninexnine_unit_1424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10121)
);

ninexnine_unit ninexnine_unit_1425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11121)
);

ninexnine_unit ninexnine_unit_1426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12121)
);

ninexnine_unit ninexnine_unit_1427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13121)
);

ninexnine_unit ninexnine_unit_1428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14121)
);

ninexnine_unit ninexnine_unit_1429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15121)
);

ninexnine_unit ninexnine_unit_1430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16121)
);

ninexnine_unit ninexnine_unit_1431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17121)
);

ninexnine_unit ninexnine_unit_1432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18121)
);

ninexnine_unit ninexnine_unit_1433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19121)
);

ninexnine_unit ninexnine_unit_1434(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A121)
);

ninexnine_unit ninexnine_unit_1435(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B121)
);

ninexnine_unit ninexnine_unit_1436(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C121)
);

ninexnine_unit ninexnine_unit_1437(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D121)
);

ninexnine_unit ninexnine_unit_1438(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E121)
);

ninexnine_unit ninexnine_unit_1439(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F121)
);

assign C1121=c10121+c11121+c12121+c13121+c14121+c15121+c16121+c17121+c18121+c19121+c1A121+c1B121+c1C121+c1D121+c1E121+c1F121;
assign A1121=(C1121>=0)?1:0;

assign P2121=A1121;

ninexnine_unit ninexnine_unit_1440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10201)
);

ninexnine_unit ninexnine_unit_1441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11201)
);

ninexnine_unit ninexnine_unit_1442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12201)
);

ninexnine_unit ninexnine_unit_1443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13201)
);

ninexnine_unit ninexnine_unit_1444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14201)
);

ninexnine_unit ninexnine_unit_1445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15201)
);

ninexnine_unit ninexnine_unit_1446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16201)
);

ninexnine_unit ninexnine_unit_1447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17201)
);

ninexnine_unit ninexnine_unit_1448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18201)
);

ninexnine_unit ninexnine_unit_1449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19201)
);

ninexnine_unit ninexnine_unit_1450(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A201)
);

ninexnine_unit ninexnine_unit_1451(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B201)
);

ninexnine_unit ninexnine_unit_1452(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C201)
);

ninexnine_unit ninexnine_unit_1453(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D201)
);

ninexnine_unit ninexnine_unit_1454(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E201)
);

ninexnine_unit ninexnine_unit_1455(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F201)
);

assign C1201=c10201+c11201+c12201+c13201+c14201+c15201+c16201+c17201+c18201+c19201+c1A201+c1B201+c1C201+c1D201+c1E201+c1F201;
assign A1201=(C1201>=0)?1:0;

assign P2201=A1201;

ninexnine_unit ninexnine_unit_1456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10211)
);

ninexnine_unit ninexnine_unit_1457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11211)
);

ninexnine_unit ninexnine_unit_1458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12211)
);

ninexnine_unit ninexnine_unit_1459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13211)
);

ninexnine_unit ninexnine_unit_1460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14211)
);

ninexnine_unit ninexnine_unit_1461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15211)
);

ninexnine_unit ninexnine_unit_1462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16211)
);

ninexnine_unit ninexnine_unit_1463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17211)
);

ninexnine_unit ninexnine_unit_1464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18211)
);

ninexnine_unit ninexnine_unit_1465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19211)
);

ninexnine_unit ninexnine_unit_1466(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A211)
);

ninexnine_unit ninexnine_unit_1467(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B211)
);

ninexnine_unit ninexnine_unit_1468(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C211)
);

ninexnine_unit ninexnine_unit_1469(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D211)
);

ninexnine_unit ninexnine_unit_1470(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E211)
);

ninexnine_unit ninexnine_unit_1471(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F211)
);

assign C1211=c10211+c11211+c12211+c13211+c14211+c15211+c16211+c17211+c18211+c19211+c1A211+c1B211+c1C211+c1D211+c1E211+c1F211;
assign A1211=(C1211>=0)?1:0;

assign P2211=A1211;

ninexnine_unit ninexnine_unit_1472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10221)
);

ninexnine_unit ninexnine_unit_1473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11221)
);

ninexnine_unit ninexnine_unit_1474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12221)
);

ninexnine_unit ninexnine_unit_1475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W11003),
				.b1(W11013),
				.b2(W11023),
				.b3(W11103),
				.b4(W11113),
				.b5(W11123),
				.b6(W11203),
				.b7(W11213),
				.b8(W11223),
				.c(c13221)
);

ninexnine_unit ninexnine_unit_1476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W11004),
				.b1(W11014),
				.b2(W11024),
				.b3(W11104),
				.b4(W11114),
				.b5(W11124),
				.b6(W11204),
				.b7(W11214),
				.b8(W11224),
				.c(c14221)
);

ninexnine_unit ninexnine_unit_1477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W11005),
				.b1(W11015),
				.b2(W11025),
				.b3(W11105),
				.b4(W11115),
				.b5(W11125),
				.b6(W11205),
				.b7(W11215),
				.b8(W11225),
				.c(c15221)
);

ninexnine_unit ninexnine_unit_1478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W11006),
				.b1(W11016),
				.b2(W11026),
				.b3(W11106),
				.b4(W11116),
				.b5(W11126),
				.b6(W11206),
				.b7(W11216),
				.b8(W11226),
				.c(c16221)
);

ninexnine_unit ninexnine_unit_1479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W11007),
				.b1(W11017),
				.b2(W11027),
				.b3(W11107),
				.b4(W11117),
				.b5(W11127),
				.b6(W11207),
				.b7(W11217),
				.b8(W11227),
				.c(c17221)
);

ninexnine_unit ninexnine_unit_1480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W11008),
				.b1(W11018),
				.b2(W11028),
				.b3(W11108),
				.b4(W11118),
				.b5(W11128),
				.b6(W11208),
				.b7(W11218),
				.b8(W11228),
				.c(c18221)
);

ninexnine_unit ninexnine_unit_1481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W11009),
				.b1(W11019),
				.b2(W11029),
				.b3(W11109),
				.b4(W11119),
				.b5(W11129),
				.b6(W11209),
				.b7(W11219),
				.b8(W11229),
				.c(c19221)
);

ninexnine_unit ninexnine_unit_1482(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1100A),
				.b1(W1101A),
				.b2(W1102A),
				.b3(W1110A),
				.b4(W1111A),
				.b5(W1112A),
				.b6(W1120A),
				.b7(W1121A),
				.b8(W1122A),
				.c(c1A221)
);

ninexnine_unit ninexnine_unit_1483(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1100B),
				.b1(W1101B),
				.b2(W1102B),
				.b3(W1110B),
				.b4(W1111B),
				.b5(W1112B),
				.b6(W1120B),
				.b7(W1121B),
				.b8(W1122B),
				.c(c1B221)
);

ninexnine_unit ninexnine_unit_1484(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1100C),
				.b1(W1101C),
				.b2(W1102C),
				.b3(W1110C),
				.b4(W1111C),
				.b5(W1112C),
				.b6(W1120C),
				.b7(W1121C),
				.b8(W1122C),
				.c(c1C221)
);

ninexnine_unit ninexnine_unit_1485(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1100D),
				.b1(W1101D),
				.b2(W1102D),
				.b3(W1110D),
				.b4(W1111D),
				.b5(W1112D),
				.b6(W1120D),
				.b7(W1121D),
				.b8(W1122D),
				.c(c1D221)
);

ninexnine_unit ninexnine_unit_1486(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1100E),
				.b1(W1101E),
				.b2(W1102E),
				.b3(W1110E),
				.b4(W1111E),
				.b5(W1112E),
				.b6(W1120E),
				.b7(W1121E),
				.b8(W1122E),
				.c(c1E221)
);

ninexnine_unit ninexnine_unit_1487(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1100F),
				.b1(W1101F),
				.b2(W1102F),
				.b3(W1110F),
				.b4(W1111F),
				.b5(W1112F),
				.b6(W1120F),
				.b7(W1121F),
				.b8(W1122F),
				.c(c1F221)
);

assign C1221=c10221+c11221+c12221+c13221+c14221+c15221+c16221+c17221+c18221+c19221+c1A221+c1B221+c1C221+c1D221+c1E221+c1F221;
assign A1221=(C1221>=0)?1:0;

assign P2221=A1221;

ninexnine_unit ninexnine_unit_1488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10002)
);

ninexnine_unit ninexnine_unit_1489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11002)
);

ninexnine_unit ninexnine_unit_1490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12002)
);

ninexnine_unit ninexnine_unit_1491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13002)
);

ninexnine_unit ninexnine_unit_1492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14002)
);

ninexnine_unit ninexnine_unit_1493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15002)
);

ninexnine_unit ninexnine_unit_1494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16002)
);

ninexnine_unit ninexnine_unit_1495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17002)
);

ninexnine_unit ninexnine_unit_1496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18002)
);

ninexnine_unit ninexnine_unit_1497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19002)
);

ninexnine_unit ninexnine_unit_1498(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A002)
);

ninexnine_unit ninexnine_unit_1499(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B002)
);

ninexnine_unit ninexnine_unit_1500(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C002)
);

ninexnine_unit ninexnine_unit_1501(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D002)
);

ninexnine_unit ninexnine_unit_1502(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E002)
);

ninexnine_unit ninexnine_unit_1503(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F002)
);

assign C1002=c10002+c11002+c12002+c13002+c14002+c15002+c16002+c17002+c18002+c19002+c1A002+c1B002+c1C002+c1D002+c1E002+c1F002;
assign A1002=(C1002>=0)?1:0;

assign P2002=A1002;

ninexnine_unit ninexnine_unit_1504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10012)
);

ninexnine_unit ninexnine_unit_1505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11012)
);

ninexnine_unit ninexnine_unit_1506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12012)
);

ninexnine_unit ninexnine_unit_1507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13012)
);

ninexnine_unit ninexnine_unit_1508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14012)
);

ninexnine_unit ninexnine_unit_1509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15012)
);

ninexnine_unit ninexnine_unit_1510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16012)
);

ninexnine_unit ninexnine_unit_1511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17012)
);

ninexnine_unit ninexnine_unit_1512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18012)
);

ninexnine_unit ninexnine_unit_1513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19012)
);

ninexnine_unit ninexnine_unit_1514(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A012)
);

ninexnine_unit ninexnine_unit_1515(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B012)
);

ninexnine_unit ninexnine_unit_1516(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C012)
);

ninexnine_unit ninexnine_unit_1517(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D012)
);

ninexnine_unit ninexnine_unit_1518(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E012)
);

ninexnine_unit ninexnine_unit_1519(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F012)
);

assign C1012=c10012+c11012+c12012+c13012+c14012+c15012+c16012+c17012+c18012+c19012+c1A012+c1B012+c1C012+c1D012+c1E012+c1F012;
assign A1012=(C1012>=0)?1:0;

assign P2012=A1012;

ninexnine_unit ninexnine_unit_1520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10022)
);

ninexnine_unit ninexnine_unit_1521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11022)
);

ninexnine_unit ninexnine_unit_1522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12022)
);

ninexnine_unit ninexnine_unit_1523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13022)
);

ninexnine_unit ninexnine_unit_1524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14022)
);

ninexnine_unit ninexnine_unit_1525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15022)
);

ninexnine_unit ninexnine_unit_1526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16022)
);

ninexnine_unit ninexnine_unit_1527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17022)
);

ninexnine_unit ninexnine_unit_1528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18022)
);

ninexnine_unit ninexnine_unit_1529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19022)
);

ninexnine_unit ninexnine_unit_1530(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A022)
);

ninexnine_unit ninexnine_unit_1531(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B022)
);

ninexnine_unit ninexnine_unit_1532(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C022)
);

ninexnine_unit ninexnine_unit_1533(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D022)
);

ninexnine_unit ninexnine_unit_1534(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E022)
);

ninexnine_unit ninexnine_unit_1535(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F022)
);

assign C1022=c10022+c11022+c12022+c13022+c14022+c15022+c16022+c17022+c18022+c19022+c1A022+c1B022+c1C022+c1D022+c1E022+c1F022;
assign A1022=(C1022>=0)?1:0;

assign P2022=A1022;

ninexnine_unit ninexnine_unit_1536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10102)
);

ninexnine_unit ninexnine_unit_1537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11102)
);

ninexnine_unit ninexnine_unit_1538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12102)
);

ninexnine_unit ninexnine_unit_1539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13102)
);

ninexnine_unit ninexnine_unit_1540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14102)
);

ninexnine_unit ninexnine_unit_1541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15102)
);

ninexnine_unit ninexnine_unit_1542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16102)
);

ninexnine_unit ninexnine_unit_1543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17102)
);

ninexnine_unit ninexnine_unit_1544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18102)
);

ninexnine_unit ninexnine_unit_1545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19102)
);

ninexnine_unit ninexnine_unit_1546(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A102)
);

ninexnine_unit ninexnine_unit_1547(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B102)
);

ninexnine_unit ninexnine_unit_1548(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C102)
);

ninexnine_unit ninexnine_unit_1549(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D102)
);

ninexnine_unit ninexnine_unit_1550(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E102)
);

ninexnine_unit ninexnine_unit_1551(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F102)
);

assign C1102=c10102+c11102+c12102+c13102+c14102+c15102+c16102+c17102+c18102+c19102+c1A102+c1B102+c1C102+c1D102+c1E102+c1F102;
assign A1102=(C1102>=0)?1:0;

assign P2102=A1102;

ninexnine_unit ninexnine_unit_1552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10112)
);

ninexnine_unit ninexnine_unit_1553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11112)
);

ninexnine_unit ninexnine_unit_1554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12112)
);

ninexnine_unit ninexnine_unit_1555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13112)
);

ninexnine_unit ninexnine_unit_1556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14112)
);

ninexnine_unit ninexnine_unit_1557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15112)
);

ninexnine_unit ninexnine_unit_1558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16112)
);

ninexnine_unit ninexnine_unit_1559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17112)
);

ninexnine_unit ninexnine_unit_1560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18112)
);

ninexnine_unit ninexnine_unit_1561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19112)
);

ninexnine_unit ninexnine_unit_1562(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A112)
);

ninexnine_unit ninexnine_unit_1563(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B112)
);

ninexnine_unit ninexnine_unit_1564(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C112)
);

ninexnine_unit ninexnine_unit_1565(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D112)
);

ninexnine_unit ninexnine_unit_1566(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E112)
);

ninexnine_unit ninexnine_unit_1567(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F112)
);

assign C1112=c10112+c11112+c12112+c13112+c14112+c15112+c16112+c17112+c18112+c19112+c1A112+c1B112+c1C112+c1D112+c1E112+c1F112;
assign A1112=(C1112>=0)?1:0;

assign P2112=A1112;

ninexnine_unit ninexnine_unit_1568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10122)
);

ninexnine_unit ninexnine_unit_1569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11122)
);

ninexnine_unit ninexnine_unit_1570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12122)
);

ninexnine_unit ninexnine_unit_1571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13122)
);

ninexnine_unit ninexnine_unit_1572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14122)
);

ninexnine_unit ninexnine_unit_1573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15122)
);

ninexnine_unit ninexnine_unit_1574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16122)
);

ninexnine_unit ninexnine_unit_1575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17122)
);

ninexnine_unit ninexnine_unit_1576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18122)
);

ninexnine_unit ninexnine_unit_1577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19122)
);

ninexnine_unit ninexnine_unit_1578(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A122)
);

ninexnine_unit ninexnine_unit_1579(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B122)
);

ninexnine_unit ninexnine_unit_1580(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C122)
);

ninexnine_unit ninexnine_unit_1581(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D122)
);

ninexnine_unit ninexnine_unit_1582(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E122)
);

ninexnine_unit ninexnine_unit_1583(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F122)
);

assign C1122=c10122+c11122+c12122+c13122+c14122+c15122+c16122+c17122+c18122+c19122+c1A122+c1B122+c1C122+c1D122+c1E122+c1F122;
assign A1122=(C1122>=0)?1:0;

assign P2122=A1122;

ninexnine_unit ninexnine_unit_1584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10202)
);

ninexnine_unit ninexnine_unit_1585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11202)
);

ninexnine_unit ninexnine_unit_1586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12202)
);

ninexnine_unit ninexnine_unit_1587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13202)
);

ninexnine_unit ninexnine_unit_1588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14202)
);

ninexnine_unit ninexnine_unit_1589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15202)
);

ninexnine_unit ninexnine_unit_1590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16202)
);

ninexnine_unit ninexnine_unit_1591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17202)
);

ninexnine_unit ninexnine_unit_1592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18202)
);

ninexnine_unit ninexnine_unit_1593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19202)
);

ninexnine_unit ninexnine_unit_1594(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A202)
);

ninexnine_unit ninexnine_unit_1595(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B202)
);

ninexnine_unit ninexnine_unit_1596(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C202)
);

ninexnine_unit ninexnine_unit_1597(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D202)
);

ninexnine_unit ninexnine_unit_1598(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E202)
);

ninexnine_unit ninexnine_unit_1599(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F202)
);

assign C1202=c10202+c11202+c12202+c13202+c14202+c15202+c16202+c17202+c18202+c19202+c1A202+c1B202+c1C202+c1D202+c1E202+c1F202;
assign A1202=(C1202>=0)?1:0;

assign P2202=A1202;

ninexnine_unit ninexnine_unit_1600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10212)
);

ninexnine_unit ninexnine_unit_1601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11212)
);

ninexnine_unit ninexnine_unit_1602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12212)
);

ninexnine_unit ninexnine_unit_1603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13212)
);

ninexnine_unit ninexnine_unit_1604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14212)
);

ninexnine_unit ninexnine_unit_1605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15212)
);

ninexnine_unit ninexnine_unit_1606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16212)
);

ninexnine_unit ninexnine_unit_1607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17212)
);

ninexnine_unit ninexnine_unit_1608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18212)
);

ninexnine_unit ninexnine_unit_1609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19212)
);

ninexnine_unit ninexnine_unit_1610(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A212)
);

ninexnine_unit ninexnine_unit_1611(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B212)
);

ninexnine_unit ninexnine_unit_1612(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C212)
);

ninexnine_unit ninexnine_unit_1613(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D212)
);

ninexnine_unit ninexnine_unit_1614(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E212)
);

ninexnine_unit ninexnine_unit_1615(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F212)
);

assign C1212=c10212+c11212+c12212+c13212+c14212+c15212+c16212+c17212+c18212+c19212+c1A212+c1B212+c1C212+c1D212+c1E212+c1F212;
assign A1212=(C1212>=0)?1:0;

assign P2212=A1212;

ninexnine_unit ninexnine_unit_1616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10222)
);

ninexnine_unit ninexnine_unit_1617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11222)
);

ninexnine_unit ninexnine_unit_1618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12222)
);

ninexnine_unit ninexnine_unit_1619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W12003),
				.b1(W12013),
				.b2(W12023),
				.b3(W12103),
				.b4(W12113),
				.b5(W12123),
				.b6(W12203),
				.b7(W12213),
				.b8(W12223),
				.c(c13222)
);

ninexnine_unit ninexnine_unit_1620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W12004),
				.b1(W12014),
				.b2(W12024),
				.b3(W12104),
				.b4(W12114),
				.b5(W12124),
				.b6(W12204),
				.b7(W12214),
				.b8(W12224),
				.c(c14222)
);

ninexnine_unit ninexnine_unit_1621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W12005),
				.b1(W12015),
				.b2(W12025),
				.b3(W12105),
				.b4(W12115),
				.b5(W12125),
				.b6(W12205),
				.b7(W12215),
				.b8(W12225),
				.c(c15222)
);

ninexnine_unit ninexnine_unit_1622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W12006),
				.b1(W12016),
				.b2(W12026),
				.b3(W12106),
				.b4(W12116),
				.b5(W12126),
				.b6(W12206),
				.b7(W12216),
				.b8(W12226),
				.c(c16222)
);

ninexnine_unit ninexnine_unit_1623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W12007),
				.b1(W12017),
				.b2(W12027),
				.b3(W12107),
				.b4(W12117),
				.b5(W12127),
				.b6(W12207),
				.b7(W12217),
				.b8(W12227),
				.c(c17222)
);

ninexnine_unit ninexnine_unit_1624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W12008),
				.b1(W12018),
				.b2(W12028),
				.b3(W12108),
				.b4(W12118),
				.b5(W12128),
				.b6(W12208),
				.b7(W12218),
				.b8(W12228),
				.c(c18222)
);

ninexnine_unit ninexnine_unit_1625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W12009),
				.b1(W12019),
				.b2(W12029),
				.b3(W12109),
				.b4(W12119),
				.b5(W12129),
				.b6(W12209),
				.b7(W12219),
				.b8(W12229),
				.c(c19222)
);

ninexnine_unit ninexnine_unit_1626(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1200A),
				.b1(W1201A),
				.b2(W1202A),
				.b3(W1210A),
				.b4(W1211A),
				.b5(W1212A),
				.b6(W1220A),
				.b7(W1221A),
				.b8(W1222A),
				.c(c1A222)
);

ninexnine_unit ninexnine_unit_1627(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1200B),
				.b1(W1201B),
				.b2(W1202B),
				.b3(W1210B),
				.b4(W1211B),
				.b5(W1212B),
				.b6(W1220B),
				.b7(W1221B),
				.b8(W1222B),
				.c(c1B222)
);

ninexnine_unit ninexnine_unit_1628(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1200C),
				.b1(W1201C),
				.b2(W1202C),
				.b3(W1210C),
				.b4(W1211C),
				.b5(W1212C),
				.b6(W1220C),
				.b7(W1221C),
				.b8(W1222C),
				.c(c1C222)
);

ninexnine_unit ninexnine_unit_1629(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1200D),
				.b1(W1201D),
				.b2(W1202D),
				.b3(W1210D),
				.b4(W1211D),
				.b5(W1212D),
				.b6(W1220D),
				.b7(W1221D),
				.b8(W1222D),
				.c(c1D222)
);

ninexnine_unit ninexnine_unit_1630(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1200E),
				.b1(W1201E),
				.b2(W1202E),
				.b3(W1210E),
				.b4(W1211E),
				.b5(W1212E),
				.b6(W1220E),
				.b7(W1221E),
				.b8(W1222E),
				.c(c1E222)
);

ninexnine_unit ninexnine_unit_1631(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1200F),
				.b1(W1201F),
				.b2(W1202F),
				.b3(W1210F),
				.b4(W1211F),
				.b5(W1212F),
				.b6(W1220F),
				.b7(W1221F),
				.b8(W1222F),
				.c(c1F222)
);

assign C1222=c10222+c11222+c12222+c13222+c14222+c15222+c16222+c17222+c18222+c19222+c1A222+c1B222+c1C222+c1D222+c1E222+c1F222;
assign A1222=(C1222>=0)?1:0;

assign P2222=A1222;

ninexnine_unit ninexnine_unit_1632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10003)
);

ninexnine_unit ninexnine_unit_1633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11003)
);

ninexnine_unit ninexnine_unit_1634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12003)
);

ninexnine_unit ninexnine_unit_1635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13003)
);

ninexnine_unit ninexnine_unit_1636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14003)
);

ninexnine_unit ninexnine_unit_1637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15003)
);

ninexnine_unit ninexnine_unit_1638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16003)
);

ninexnine_unit ninexnine_unit_1639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17003)
);

ninexnine_unit ninexnine_unit_1640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18003)
);

ninexnine_unit ninexnine_unit_1641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19003)
);

ninexnine_unit ninexnine_unit_1642(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A003)
);

ninexnine_unit ninexnine_unit_1643(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B003)
);

ninexnine_unit ninexnine_unit_1644(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C003)
);

ninexnine_unit ninexnine_unit_1645(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D003)
);

ninexnine_unit ninexnine_unit_1646(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E003)
);

ninexnine_unit ninexnine_unit_1647(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F003)
);

assign C1003=c10003+c11003+c12003+c13003+c14003+c15003+c16003+c17003+c18003+c19003+c1A003+c1B003+c1C003+c1D003+c1E003+c1F003;
assign A1003=(C1003>=0)?1:0;

assign P2003=A1003;

ninexnine_unit ninexnine_unit_1648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10013)
);

ninexnine_unit ninexnine_unit_1649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11013)
);

ninexnine_unit ninexnine_unit_1650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12013)
);

ninexnine_unit ninexnine_unit_1651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13013)
);

ninexnine_unit ninexnine_unit_1652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14013)
);

ninexnine_unit ninexnine_unit_1653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15013)
);

ninexnine_unit ninexnine_unit_1654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16013)
);

ninexnine_unit ninexnine_unit_1655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17013)
);

ninexnine_unit ninexnine_unit_1656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18013)
);

ninexnine_unit ninexnine_unit_1657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19013)
);

ninexnine_unit ninexnine_unit_1658(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A013)
);

ninexnine_unit ninexnine_unit_1659(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B013)
);

ninexnine_unit ninexnine_unit_1660(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C013)
);

ninexnine_unit ninexnine_unit_1661(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D013)
);

ninexnine_unit ninexnine_unit_1662(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E013)
);

ninexnine_unit ninexnine_unit_1663(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F013)
);

assign C1013=c10013+c11013+c12013+c13013+c14013+c15013+c16013+c17013+c18013+c19013+c1A013+c1B013+c1C013+c1D013+c1E013+c1F013;
assign A1013=(C1013>=0)?1:0;

assign P2013=A1013;

ninexnine_unit ninexnine_unit_1664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10023)
);

ninexnine_unit ninexnine_unit_1665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11023)
);

ninexnine_unit ninexnine_unit_1666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12023)
);

ninexnine_unit ninexnine_unit_1667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13023)
);

ninexnine_unit ninexnine_unit_1668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14023)
);

ninexnine_unit ninexnine_unit_1669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15023)
);

ninexnine_unit ninexnine_unit_1670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16023)
);

ninexnine_unit ninexnine_unit_1671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17023)
);

ninexnine_unit ninexnine_unit_1672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18023)
);

ninexnine_unit ninexnine_unit_1673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19023)
);

ninexnine_unit ninexnine_unit_1674(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A023)
);

ninexnine_unit ninexnine_unit_1675(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B023)
);

ninexnine_unit ninexnine_unit_1676(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C023)
);

ninexnine_unit ninexnine_unit_1677(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D023)
);

ninexnine_unit ninexnine_unit_1678(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E023)
);

ninexnine_unit ninexnine_unit_1679(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F023)
);

assign C1023=c10023+c11023+c12023+c13023+c14023+c15023+c16023+c17023+c18023+c19023+c1A023+c1B023+c1C023+c1D023+c1E023+c1F023;
assign A1023=(C1023>=0)?1:0;

assign P2023=A1023;

ninexnine_unit ninexnine_unit_1680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10103)
);

ninexnine_unit ninexnine_unit_1681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11103)
);

ninexnine_unit ninexnine_unit_1682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12103)
);

ninexnine_unit ninexnine_unit_1683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13103)
);

ninexnine_unit ninexnine_unit_1684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14103)
);

ninexnine_unit ninexnine_unit_1685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15103)
);

ninexnine_unit ninexnine_unit_1686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16103)
);

ninexnine_unit ninexnine_unit_1687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17103)
);

ninexnine_unit ninexnine_unit_1688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18103)
);

ninexnine_unit ninexnine_unit_1689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19103)
);

ninexnine_unit ninexnine_unit_1690(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A103)
);

ninexnine_unit ninexnine_unit_1691(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B103)
);

ninexnine_unit ninexnine_unit_1692(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C103)
);

ninexnine_unit ninexnine_unit_1693(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D103)
);

ninexnine_unit ninexnine_unit_1694(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E103)
);

ninexnine_unit ninexnine_unit_1695(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F103)
);

assign C1103=c10103+c11103+c12103+c13103+c14103+c15103+c16103+c17103+c18103+c19103+c1A103+c1B103+c1C103+c1D103+c1E103+c1F103;
assign A1103=(C1103>=0)?1:0;

assign P2103=A1103;

ninexnine_unit ninexnine_unit_1696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10113)
);

ninexnine_unit ninexnine_unit_1697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11113)
);

ninexnine_unit ninexnine_unit_1698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12113)
);

ninexnine_unit ninexnine_unit_1699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13113)
);

ninexnine_unit ninexnine_unit_1700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14113)
);

ninexnine_unit ninexnine_unit_1701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15113)
);

ninexnine_unit ninexnine_unit_1702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16113)
);

ninexnine_unit ninexnine_unit_1703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17113)
);

ninexnine_unit ninexnine_unit_1704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18113)
);

ninexnine_unit ninexnine_unit_1705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19113)
);

ninexnine_unit ninexnine_unit_1706(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A113)
);

ninexnine_unit ninexnine_unit_1707(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B113)
);

ninexnine_unit ninexnine_unit_1708(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C113)
);

ninexnine_unit ninexnine_unit_1709(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D113)
);

ninexnine_unit ninexnine_unit_1710(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E113)
);

ninexnine_unit ninexnine_unit_1711(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F113)
);

assign C1113=c10113+c11113+c12113+c13113+c14113+c15113+c16113+c17113+c18113+c19113+c1A113+c1B113+c1C113+c1D113+c1E113+c1F113;
assign A1113=(C1113>=0)?1:0;

assign P2113=A1113;

ninexnine_unit ninexnine_unit_1712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10123)
);

ninexnine_unit ninexnine_unit_1713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11123)
);

ninexnine_unit ninexnine_unit_1714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12123)
);

ninexnine_unit ninexnine_unit_1715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13123)
);

ninexnine_unit ninexnine_unit_1716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14123)
);

ninexnine_unit ninexnine_unit_1717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15123)
);

ninexnine_unit ninexnine_unit_1718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16123)
);

ninexnine_unit ninexnine_unit_1719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17123)
);

ninexnine_unit ninexnine_unit_1720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18123)
);

ninexnine_unit ninexnine_unit_1721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19123)
);

ninexnine_unit ninexnine_unit_1722(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A123)
);

ninexnine_unit ninexnine_unit_1723(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B123)
);

ninexnine_unit ninexnine_unit_1724(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C123)
);

ninexnine_unit ninexnine_unit_1725(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D123)
);

ninexnine_unit ninexnine_unit_1726(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E123)
);

ninexnine_unit ninexnine_unit_1727(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F123)
);

assign C1123=c10123+c11123+c12123+c13123+c14123+c15123+c16123+c17123+c18123+c19123+c1A123+c1B123+c1C123+c1D123+c1E123+c1F123;
assign A1123=(C1123>=0)?1:0;

assign P2123=A1123;

ninexnine_unit ninexnine_unit_1728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10203)
);

ninexnine_unit ninexnine_unit_1729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11203)
);

ninexnine_unit ninexnine_unit_1730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12203)
);

ninexnine_unit ninexnine_unit_1731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13203)
);

ninexnine_unit ninexnine_unit_1732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14203)
);

ninexnine_unit ninexnine_unit_1733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15203)
);

ninexnine_unit ninexnine_unit_1734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16203)
);

ninexnine_unit ninexnine_unit_1735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17203)
);

ninexnine_unit ninexnine_unit_1736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18203)
);

ninexnine_unit ninexnine_unit_1737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19203)
);

ninexnine_unit ninexnine_unit_1738(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A203)
);

ninexnine_unit ninexnine_unit_1739(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B203)
);

ninexnine_unit ninexnine_unit_1740(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C203)
);

ninexnine_unit ninexnine_unit_1741(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D203)
);

ninexnine_unit ninexnine_unit_1742(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E203)
);

ninexnine_unit ninexnine_unit_1743(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F203)
);

assign C1203=c10203+c11203+c12203+c13203+c14203+c15203+c16203+c17203+c18203+c19203+c1A203+c1B203+c1C203+c1D203+c1E203+c1F203;
assign A1203=(C1203>=0)?1:0;

assign P2203=A1203;

ninexnine_unit ninexnine_unit_1744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10213)
);

ninexnine_unit ninexnine_unit_1745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11213)
);

ninexnine_unit ninexnine_unit_1746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12213)
);

ninexnine_unit ninexnine_unit_1747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13213)
);

ninexnine_unit ninexnine_unit_1748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14213)
);

ninexnine_unit ninexnine_unit_1749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15213)
);

ninexnine_unit ninexnine_unit_1750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16213)
);

ninexnine_unit ninexnine_unit_1751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17213)
);

ninexnine_unit ninexnine_unit_1752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18213)
);

ninexnine_unit ninexnine_unit_1753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19213)
);

ninexnine_unit ninexnine_unit_1754(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A213)
);

ninexnine_unit ninexnine_unit_1755(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B213)
);

ninexnine_unit ninexnine_unit_1756(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C213)
);

ninexnine_unit ninexnine_unit_1757(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D213)
);

ninexnine_unit ninexnine_unit_1758(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E213)
);

ninexnine_unit ninexnine_unit_1759(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F213)
);

assign C1213=c10213+c11213+c12213+c13213+c14213+c15213+c16213+c17213+c18213+c19213+c1A213+c1B213+c1C213+c1D213+c1E213+c1F213;
assign A1213=(C1213>=0)?1:0;

assign P2213=A1213;

ninexnine_unit ninexnine_unit_1760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10223)
);

ninexnine_unit ninexnine_unit_1761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11223)
);

ninexnine_unit ninexnine_unit_1762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12223)
);

ninexnine_unit ninexnine_unit_1763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W13003),
				.b1(W13013),
				.b2(W13023),
				.b3(W13103),
				.b4(W13113),
				.b5(W13123),
				.b6(W13203),
				.b7(W13213),
				.b8(W13223),
				.c(c13223)
);

ninexnine_unit ninexnine_unit_1764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W13004),
				.b1(W13014),
				.b2(W13024),
				.b3(W13104),
				.b4(W13114),
				.b5(W13124),
				.b6(W13204),
				.b7(W13214),
				.b8(W13224),
				.c(c14223)
);

ninexnine_unit ninexnine_unit_1765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W13005),
				.b1(W13015),
				.b2(W13025),
				.b3(W13105),
				.b4(W13115),
				.b5(W13125),
				.b6(W13205),
				.b7(W13215),
				.b8(W13225),
				.c(c15223)
);

ninexnine_unit ninexnine_unit_1766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W13006),
				.b1(W13016),
				.b2(W13026),
				.b3(W13106),
				.b4(W13116),
				.b5(W13126),
				.b6(W13206),
				.b7(W13216),
				.b8(W13226),
				.c(c16223)
);

ninexnine_unit ninexnine_unit_1767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W13007),
				.b1(W13017),
				.b2(W13027),
				.b3(W13107),
				.b4(W13117),
				.b5(W13127),
				.b6(W13207),
				.b7(W13217),
				.b8(W13227),
				.c(c17223)
);

ninexnine_unit ninexnine_unit_1768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W13008),
				.b1(W13018),
				.b2(W13028),
				.b3(W13108),
				.b4(W13118),
				.b5(W13128),
				.b6(W13208),
				.b7(W13218),
				.b8(W13228),
				.c(c18223)
);

ninexnine_unit ninexnine_unit_1769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W13009),
				.b1(W13019),
				.b2(W13029),
				.b3(W13109),
				.b4(W13119),
				.b5(W13129),
				.b6(W13209),
				.b7(W13219),
				.b8(W13229),
				.c(c19223)
);

ninexnine_unit ninexnine_unit_1770(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1300A),
				.b1(W1301A),
				.b2(W1302A),
				.b3(W1310A),
				.b4(W1311A),
				.b5(W1312A),
				.b6(W1320A),
				.b7(W1321A),
				.b8(W1322A),
				.c(c1A223)
);

ninexnine_unit ninexnine_unit_1771(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1300B),
				.b1(W1301B),
				.b2(W1302B),
				.b3(W1310B),
				.b4(W1311B),
				.b5(W1312B),
				.b6(W1320B),
				.b7(W1321B),
				.b8(W1322B),
				.c(c1B223)
);

ninexnine_unit ninexnine_unit_1772(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1300C),
				.b1(W1301C),
				.b2(W1302C),
				.b3(W1310C),
				.b4(W1311C),
				.b5(W1312C),
				.b6(W1320C),
				.b7(W1321C),
				.b8(W1322C),
				.c(c1C223)
);

ninexnine_unit ninexnine_unit_1773(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1300D),
				.b1(W1301D),
				.b2(W1302D),
				.b3(W1310D),
				.b4(W1311D),
				.b5(W1312D),
				.b6(W1320D),
				.b7(W1321D),
				.b8(W1322D),
				.c(c1D223)
);

ninexnine_unit ninexnine_unit_1774(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1300E),
				.b1(W1301E),
				.b2(W1302E),
				.b3(W1310E),
				.b4(W1311E),
				.b5(W1312E),
				.b6(W1320E),
				.b7(W1321E),
				.b8(W1322E),
				.c(c1E223)
);

ninexnine_unit ninexnine_unit_1775(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1300F),
				.b1(W1301F),
				.b2(W1302F),
				.b3(W1310F),
				.b4(W1311F),
				.b5(W1312F),
				.b6(W1320F),
				.b7(W1321F),
				.b8(W1322F),
				.c(c1F223)
);

assign C1223=c10223+c11223+c12223+c13223+c14223+c15223+c16223+c17223+c18223+c19223+c1A223+c1B223+c1C223+c1D223+c1E223+c1F223;
assign A1223=(C1223>=0)?1:0;

assign P2223=A1223;

ninexnine_unit ninexnine_unit_1776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10004)
);

ninexnine_unit ninexnine_unit_1777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11004)
);

ninexnine_unit ninexnine_unit_1778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12004)
);

ninexnine_unit ninexnine_unit_1779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13004)
);

ninexnine_unit ninexnine_unit_1780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14004)
);

ninexnine_unit ninexnine_unit_1781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15004)
);

ninexnine_unit ninexnine_unit_1782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16004)
);

ninexnine_unit ninexnine_unit_1783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17004)
);

ninexnine_unit ninexnine_unit_1784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18004)
);

ninexnine_unit ninexnine_unit_1785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19004)
);

ninexnine_unit ninexnine_unit_1786(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A004)
);

ninexnine_unit ninexnine_unit_1787(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B004)
);

ninexnine_unit ninexnine_unit_1788(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C004)
);

ninexnine_unit ninexnine_unit_1789(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D004)
);

ninexnine_unit ninexnine_unit_1790(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E004)
);

ninexnine_unit ninexnine_unit_1791(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F004)
);

assign C1004=c10004+c11004+c12004+c13004+c14004+c15004+c16004+c17004+c18004+c19004+c1A004+c1B004+c1C004+c1D004+c1E004+c1F004;
assign A1004=(C1004>=0)?1:0;

assign P2004=A1004;

ninexnine_unit ninexnine_unit_1792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10014)
);

ninexnine_unit ninexnine_unit_1793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11014)
);

ninexnine_unit ninexnine_unit_1794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12014)
);

ninexnine_unit ninexnine_unit_1795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13014)
);

ninexnine_unit ninexnine_unit_1796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14014)
);

ninexnine_unit ninexnine_unit_1797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15014)
);

ninexnine_unit ninexnine_unit_1798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16014)
);

ninexnine_unit ninexnine_unit_1799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17014)
);

ninexnine_unit ninexnine_unit_1800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18014)
);

ninexnine_unit ninexnine_unit_1801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19014)
);

ninexnine_unit ninexnine_unit_1802(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A014)
);

ninexnine_unit ninexnine_unit_1803(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B014)
);

ninexnine_unit ninexnine_unit_1804(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C014)
);

ninexnine_unit ninexnine_unit_1805(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D014)
);

ninexnine_unit ninexnine_unit_1806(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E014)
);

ninexnine_unit ninexnine_unit_1807(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F014)
);

assign C1014=c10014+c11014+c12014+c13014+c14014+c15014+c16014+c17014+c18014+c19014+c1A014+c1B014+c1C014+c1D014+c1E014+c1F014;
assign A1014=(C1014>=0)?1:0;

assign P2014=A1014;

ninexnine_unit ninexnine_unit_1808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10024)
);

ninexnine_unit ninexnine_unit_1809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11024)
);

ninexnine_unit ninexnine_unit_1810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12024)
);

ninexnine_unit ninexnine_unit_1811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13024)
);

ninexnine_unit ninexnine_unit_1812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14024)
);

ninexnine_unit ninexnine_unit_1813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15024)
);

ninexnine_unit ninexnine_unit_1814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16024)
);

ninexnine_unit ninexnine_unit_1815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17024)
);

ninexnine_unit ninexnine_unit_1816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18024)
);

ninexnine_unit ninexnine_unit_1817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19024)
);

ninexnine_unit ninexnine_unit_1818(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A024)
);

ninexnine_unit ninexnine_unit_1819(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B024)
);

ninexnine_unit ninexnine_unit_1820(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C024)
);

ninexnine_unit ninexnine_unit_1821(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D024)
);

ninexnine_unit ninexnine_unit_1822(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E024)
);

ninexnine_unit ninexnine_unit_1823(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F024)
);

assign C1024=c10024+c11024+c12024+c13024+c14024+c15024+c16024+c17024+c18024+c19024+c1A024+c1B024+c1C024+c1D024+c1E024+c1F024;
assign A1024=(C1024>=0)?1:0;

assign P2024=A1024;

ninexnine_unit ninexnine_unit_1824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10104)
);

ninexnine_unit ninexnine_unit_1825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11104)
);

ninexnine_unit ninexnine_unit_1826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12104)
);

ninexnine_unit ninexnine_unit_1827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13104)
);

ninexnine_unit ninexnine_unit_1828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14104)
);

ninexnine_unit ninexnine_unit_1829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15104)
);

ninexnine_unit ninexnine_unit_1830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16104)
);

ninexnine_unit ninexnine_unit_1831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17104)
);

ninexnine_unit ninexnine_unit_1832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18104)
);

ninexnine_unit ninexnine_unit_1833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19104)
);

ninexnine_unit ninexnine_unit_1834(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A104)
);

ninexnine_unit ninexnine_unit_1835(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B104)
);

ninexnine_unit ninexnine_unit_1836(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C104)
);

ninexnine_unit ninexnine_unit_1837(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D104)
);

ninexnine_unit ninexnine_unit_1838(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E104)
);

ninexnine_unit ninexnine_unit_1839(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F104)
);

assign C1104=c10104+c11104+c12104+c13104+c14104+c15104+c16104+c17104+c18104+c19104+c1A104+c1B104+c1C104+c1D104+c1E104+c1F104;
assign A1104=(C1104>=0)?1:0;

assign P2104=A1104;

ninexnine_unit ninexnine_unit_1840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10114)
);

ninexnine_unit ninexnine_unit_1841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11114)
);

ninexnine_unit ninexnine_unit_1842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12114)
);

ninexnine_unit ninexnine_unit_1843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13114)
);

ninexnine_unit ninexnine_unit_1844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14114)
);

ninexnine_unit ninexnine_unit_1845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15114)
);

ninexnine_unit ninexnine_unit_1846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16114)
);

ninexnine_unit ninexnine_unit_1847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17114)
);

ninexnine_unit ninexnine_unit_1848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18114)
);

ninexnine_unit ninexnine_unit_1849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19114)
);

ninexnine_unit ninexnine_unit_1850(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A114)
);

ninexnine_unit ninexnine_unit_1851(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B114)
);

ninexnine_unit ninexnine_unit_1852(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C114)
);

ninexnine_unit ninexnine_unit_1853(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D114)
);

ninexnine_unit ninexnine_unit_1854(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E114)
);

ninexnine_unit ninexnine_unit_1855(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F114)
);

assign C1114=c10114+c11114+c12114+c13114+c14114+c15114+c16114+c17114+c18114+c19114+c1A114+c1B114+c1C114+c1D114+c1E114+c1F114;
assign A1114=(C1114>=0)?1:0;

assign P2114=A1114;

ninexnine_unit ninexnine_unit_1856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10124)
);

ninexnine_unit ninexnine_unit_1857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11124)
);

ninexnine_unit ninexnine_unit_1858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12124)
);

ninexnine_unit ninexnine_unit_1859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13124)
);

ninexnine_unit ninexnine_unit_1860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14124)
);

ninexnine_unit ninexnine_unit_1861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15124)
);

ninexnine_unit ninexnine_unit_1862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16124)
);

ninexnine_unit ninexnine_unit_1863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17124)
);

ninexnine_unit ninexnine_unit_1864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18124)
);

ninexnine_unit ninexnine_unit_1865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19124)
);

ninexnine_unit ninexnine_unit_1866(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A124)
);

ninexnine_unit ninexnine_unit_1867(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B124)
);

ninexnine_unit ninexnine_unit_1868(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C124)
);

ninexnine_unit ninexnine_unit_1869(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D124)
);

ninexnine_unit ninexnine_unit_1870(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E124)
);

ninexnine_unit ninexnine_unit_1871(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F124)
);

assign C1124=c10124+c11124+c12124+c13124+c14124+c15124+c16124+c17124+c18124+c19124+c1A124+c1B124+c1C124+c1D124+c1E124+c1F124;
assign A1124=(C1124>=0)?1:0;

assign P2124=A1124;

ninexnine_unit ninexnine_unit_1872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10204)
);

ninexnine_unit ninexnine_unit_1873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11204)
);

ninexnine_unit ninexnine_unit_1874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12204)
);

ninexnine_unit ninexnine_unit_1875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13204)
);

ninexnine_unit ninexnine_unit_1876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14204)
);

ninexnine_unit ninexnine_unit_1877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15204)
);

ninexnine_unit ninexnine_unit_1878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16204)
);

ninexnine_unit ninexnine_unit_1879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17204)
);

ninexnine_unit ninexnine_unit_1880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18204)
);

ninexnine_unit ninexnine_unit_1881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19204)
);

ninexnine_unit ninexnine_unit_1882(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A204)
);

ninexnine_unit ninexnine_unit_1883(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B204)
);

ninexnine_unit ninexnine_unit_1884(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C204)
);

ninexnine_unit ninexnine_unit_1885(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D204)
);

ninexnine_unit ninexnine_unit_1886(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E204)
);

ninexnine_unit ninexnine_unit_1887(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F204)
);

assign C1204=c10204+c11204+c12204+c13204+c14204+c15204+c16204+c17204+c18204+c19204+c1A204+c1B204+c1C204+c1D204+c1E204+c1F204;
assign A1204=(C1204>=0)?1:0;

assign P2204=A1204;

ninexnine_unit ninexnine_unit_1888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10214)
);

ninexnine_unit ninexnine_unit_1889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11214)
);

ninexnine_unit ninexnine_unit_1890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12214)
);

ninexnine_unit ninexnine_unit_1891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13214)
);

ninexnine_unit ninexnine_unit_1892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14214)
);

ninexnine_unit ninexnine_unit_1893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15214)
);

ninexnine_unit ninexnine_unit_1894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16214)
);

ninexnine_unit ninexnine_unit_1895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17214)
);

ninexnine_unit ninexnine_unit_1896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18214)
);

ninexnine_unit ninexnine_unit_1897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19214)
);

ninexnine_unit ninexnine_unit_1898(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A214)
);

ninexnine_unit ninexnine_unit_1899(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B214)
);

ninexnine_unit ninexnine_unit_1900(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C214)
);

ninexnine_unit ninexnine_unit_1901(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D214)
);

ninexnine_unit ninexnine_unit_1902(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E214)
);

ninexnine_unit ninexnine_unit_1903(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F214)
);

assign C1214=c10214+c11214+c12214+c13214+c14214+c15214+c16214+c17214+c18214+c19214+c1A214+c1B214+c1C214+c1D214+c1E214+c1F214;
assign A1214=(C1214>=0)?1:0;

assign P2214=A1214;

ninexnine_unit ninexnine_unit_1904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10224)
);

ninexnine_unit ninexnine_unit_1905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11224)
);

ninexnine_unit ninexnine_unit_1906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12224)
);

ninexnine_unit ninexnine_unit_1907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W14003),
				.b1(W14013),
				.b2(W14023),
				.b3(W14103),
				.b4(W14113),
				.b5(W14123),
				.b6(W14203),
				.b7(W14213),
				.b8(W14223),
				.c(c13224)
);

ninexnine_unit ninexnine_unit_1908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W14004),
				.b1(W14014),
				.b2(W14024),
				.b3(W14104),
				.b4(W14114),
				.b5(W14124),
				.b6(W14204),
				.b7(W14214),
				.b8(W14224),
				.c(c14224)
);

ninexnine_unit ninexnine_unit_1909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W14005),
				.b1(W14015),
				.b2(W14025),
				.b3(W14105),
				.b4(W14115),
				.b5(W14125),
				.b6(W14205),
				.b7(W14215),
				.b8(W14225),
				.c(c15224)
);

ninexnine_unit ninexnine_unit_1910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W14006),
				.b1(W14016),
				.b2(W14026),
				.b3(W14106),
				.b4(W14116),
				.b5(W14126),
				.b6(W14206),
				.b7(W14216),
				.b8(W14226),
				.c(c16224)
);

ninexnine_unit ninexnine_unit_1911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W14007),
				.b1(W14017),
				.b2(W14027),
				.b3(W14107),
				.b4(W14117),
				.b5(W14127),
				.b6(W14207),
				.b7(W14217),
				.b8(W14227),
				.c(c17224)
);

ninexnine_unit ninexnine_unit_1912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W14008),
				.b1(W14018),
				.b2(W14028),
				.b3(W14108),
				.b4(W14118),
				.b5(W14128),
				.b6(W14208),
				.b7(W14218),
				.b8(W14228),
				.c(c18224)
);

ninexnine_unit ninexnine_unit_1913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W14009),
				.b1(W14019),
				.b2(W14029),
				.b3(W14109),
				.b4(W14119),
				.b5(W14129),
				.b6(W14209),
				.b7(W14219),
				.b8(W14229),
				.c(c19224)
);

ninexnine_unit ninexnine_unit_1914(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1400A),
				.b1(W1401A),
				.b2(W1402A),
				.b3(W1410A),
				.b4(W1411A),
				.b5(W1412A),
				.b6(W1420A),
				.b7(W1421A),
				.b8(W1422A),
				.c(c1A224)
);

ninexnine_unit ninexnine_unit_1915(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1400B),
				.b1(W1401B),
				.b2(W1402B),
				.b3(W1410B),
				.b4(W1411B),
				.b5(W1412B),
				.b6(W1420B),
				.b7(W1421B),
				.b8(W1422B),
				.c(c1B224)
);

ninexnine_unit ninexnine_unit_1916(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1400C),
				.b1(W1401C),
				.b2(W1402C),
				.b3(W1410C),
				.b4(W1411C),
				.b5(W1412C),
				.b6(W1420C),
				.b7(W1421C),
				.b8(W1422C),
				.c(c1C224)
);

ninexnine_unit ninexnine_unit_1917(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1400D),
				.b1(W1401D),
				.b2(W1402D),
				.b3(W1410D),
				.b4(W1411D),
				.b5(W1412D),
				.b6(W1420D),
				.b7(W1421D),
				.b8(W1422D),
				.c(c1D224)
);

ninexnine_unit ninexnine_unit_1918(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1400E),
				.b1(W1401E),
				.b2(W1402E),
				.b3(W1410E),
				.b4(W1411E),
				.b5(W1412E),
				.b6(W1420E),
				.b7(W1421E),
				.b8(W1422E),
				.c(c1E224)
);

ninexnine_unit ninexnine_unit_1919(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1400F),
				.b1(W1401F),
				.b2(W1402F),
				.b3(W1410F),
				.b4(W1411F),
				.b5(W1412F),
				.b6(W1420F),
				.b7(W1421F),
				.b8(W1422F),
				.c(c1F224)
);

assign C1224=c10224+c11224+c12224+c13224+c14224+c15224+c16224+c17224+c18224+c19224+c1A224+c1B224+c1C224+c1D224+c1E224+c1F224;
assign A1224=(C1224>=0)?1:0;

assign P2224=A1224;

ninexnine_unit ninexnine_unit_1920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10005)
);

ninexnine_unit ninexnine_unit_1921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11005)
);

ninexnine_unit ninexnine_unit_1922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12005)
);

ninexnine_unit ninexnine_unit_1923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13005)
);

ninexnine_unit ninexnine_unit_1924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14005)
);

ninexnine_unit ninexnine_unit_1925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15005)
);

ninexnine_unit ninexnine_unit_1926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16005)
);

ninexnine_unit ninexnine_unit_1927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17005)
);

ninexnine_unit ninexnine_unit_1928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18005)
);

ninexnine_unit ninexnine_unit_1929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19005)
);

ninexnine_unit ninexnine_unit_1930(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A005)
);

ninexnine_unit ninexnine_unit_1931(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B005)
);

ninexnine_unit ninexnine_unit_1932(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C005)
);

ninexnine_unit ninexnine_unit_1933(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D005)
);

ninexnine_unit ninexnine_unit_1934(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E005)
);

ninexnine_unit ninexnine_unit_1935(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F005)
);

assign C1005=c10005+c11005+c12005+c13005+c14005+c15005+c16005+c17005+c18005+c19005+c1A005+c1B005+c1C005+c1D005+c1E005+c1F005;
assign A1005=(C1005>=0)?1:0;

assign P2005=A1005;

ninexnine_unit ninexnine_unit_1936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10015)
);

ninexnine_unit ninexnine_unit_1937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11015)
);

ninexnine_unit ninexnine_unit_1938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12015)
);

ninexnine_unit ninexnine_unit_1939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13015)
);

ninexnine_unit ninexnine_unit_1940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14015)
);

ninexnine_unit ninexnine_unit_1941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15015)
);

ninexnine_unit ninexnine_unit_1942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16015)
);

ninexnine_unit ninexnine_unit_1943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17015)
);

ninexnine_unit ninexnine_unit_1944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18015)
);

ninexnine_unit ninexnine_unit_1945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19015)
);

ninexnine_unit ninexnine_unit_1946(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A015)
);

ninexnine_unit ninexnine_unit_1947(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B015)
);

ninexnine_unit ninexnine_unit_1948(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C015)
);

ninexnine_unit ninexnine_unit_1949(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D015)
);

ninexnine_unit ninexnine_unit_1950(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E015)
);

ninexnine_unit ninexnine_unit_1951(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F015)
);

assign C1015=c10015+c11015+c12015+c13015+c14015+c15015+c16015+c17015+c18015+c19015+c1A015+c1B015+c1C015+c1D015+c1E015+c1F015;
assign A1015=(C1015>=0)?1:0;

assign P2015=A1015;

ninexnine_unit ninexnine_unit_1952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10025)
);

ninexnine_unit ninexnine_unit_1953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11025)
);

ninexnine_unit ninexnine_unit_1954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12025)
);

ninexnine_unit ninexnine_unit_1955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13025)
);

ninexnine_unit ninexnine_unit_1956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14025)
);

ninexnine_unit ninexnine_unit_1957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15025)
);

ninexnine_unit ninexnine_unit_1958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16025)
);

ninexnine_unit ninexnine_unit_1959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17025)
);

ninexnine_unit ninexnine_unit_1960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18025)
);

ninexnine_unit ninexnine_unit_1961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19025)
);

ninexnine_unit ninexnine_unit_1962(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A025)
);

ninexnine_unit ninexnine_unit_1963(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B025)
);

ninexnine_unit ninexnine_unit_1964(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C025)
);

ninexnine_unit ninexnine_unit_1965(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D025)
);

ninexnine_unit ninexnine_unit_1966(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E025)
);

ninexnine_unit ninexnine_unit_1967(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F025)
);

assign C1025=c10025+c11025+c12025+c13025+c14025+c15025+c16025+c17025+c18025+c19025+c1A025+c1B025+c1C025+c1D025+c1E025+c1F025;
assign A1025=(C1025>=0)?1:0;

assign P2025=A1025;

ninexnine_unit ninexnine_unit_1968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10105)
);

ninexnine_unit ninexnine_unit_1969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11105)
);

ninexnine_unit ninexnine_unit_1970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12105)
);

ninexnine_unit ninexnine_unit_1971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13105)
);

ninexnine_unit ninexnine_unit_1972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14105)
);

ninexnine_unit ninexnine_unit_1973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15105)
);

ninexnine_unit ninexnine_unit_1974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16105)
);

ninexnine_unit ninexnine_unit_1975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17105)
);

ninexnine_unit ninexnine_unit_1976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18105)
);

ninexnine_unit ninexnine_unit_1977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19105)
);

ninexnine_unit ninexnine_unit_1978(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A105)
);

ninexnine_unit ninexnine_unit_1979(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B105)
);

ninexnine_unit ninexnine_unit_1980(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C105)
);

ninexnine_unit ninexnine_unit_1981(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D105)
);

ninexnine_unit ninexnine_unit_1982(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E105)
);

ninexnine_unit ninexnine_unit_1983(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F105)
);

assign C1105=c10105+c11105+c12105+c13105+c14105+c15105+c16105+c17105+c18105+c19105+c1A105+c1B105+c1C105+c1D105+c1E105+c1F105;
assign A1105=(C1105>=0)?1:0;

assign P2105=A1105;

ninexnine_unit ninexnine_unit_1984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10115)
);

ninexnine_unit ninexnine_unit_1985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11115)
);

ninexnine_unit ninexnine_unit_1986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12115)
);

ninexnine_unit ninexnine_unit_1987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13115)
);

ninexnine_unit ninexnine_unit_1988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14115)
);

ninexnine_unit ninexnine_unit_1989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15115)
);

ninexnine_unit ninexnine_unit_1990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16115)
);

ninexnine_unit ninexnine_unit_1991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17115)
);

ninexnine_unit ninexnine_unit_1992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18115)
);

ninexnine_unit ninexnine_unit_1993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19115)
);

ninexnine_unit ninexnine_unit_1994(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A115)
);

ninexnine_unit ninexnine_unit_1995(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B115)
);

ninexnine_unit ninexnine_unit_1996(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C115)
);

ninexnine_unit ninexnine_unit_1997(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D115)
);

ninexnine_unit ninexnine_unit_1998(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E115)
);

ninexnine_unit ninexnine_unit_1999(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F115)
);

assign C1115=c10115+c11115+c12115+c13115+c14115+c15115+c16115+c17115+c18115+c19115+c1A115+c1B115+c1C115+c1D115+c1E115+c1F115;
assign A1115=(C1115>=0)?1:0;

assign P2115=A1115;

ninexnine_unit ninexnine_unit_2000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10125)
);

ninexnine_unit ninexnine_unit_2001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11125)
);

ninexnine_unit ninexnine_unit_2002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12125)
);

ninexnine_unit ninexnine_unit_2003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13125)
);

ninexnine_unit ninexnine_unit_2004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14125)
);

ninexnine_unit ninexnine_unit_2005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15125)
);

ninexnine_unit ninexnine_unit_2006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16125)
);

ninexnine_unit ninexnine_unit_2007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17125)
);

ninexnine_unit ninexnine_unit_2008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18125)
);

ninexnine_unit ninexnine_unit_2009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19125)
);

ninexnine_unit ninexnine_unit_2010(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A125)
);

ninexnine_unit ninexnine_unit_2011(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B125)
);

ninexnine_unit ninexnine_unit_2012(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C125)
);

ninexnine_unit ninexnine_unit_2013(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D125)
);

ninexnine_unit ninexnine_unit_2014(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E125)
);

ninexnine_unit ninexnine_unit_2015(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F125)
);

assign C1125=c10125+c11125+c12125+c13125+c14125+c15125+c16125+c17125+c18125+c19125+c1A125+c1B125+c1C125+c1D125+c1E125+c1F125;
assign A1125=(C1125>=0)?1:0;

assign P2125=A1125;

ninexnine_unit ninexnine_unit_2016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10205)
);

ninexnine_unit ninexnine_unit_2017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11205)
);

ninexnine_unit ninexnine_unit_2018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12205)
);

ninexnine_unit ninexnine_unit_2019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13205)
);

ninexnine_unit ninexnine_unit_2020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14205)
);

ninexnine_unit ninexnine_unit_2021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15205)
);

ninexnine_unit ninexnine_unit_2022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16205)
);

ninexnine_unit ninexnine_unit_2023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17205)
);

ninexnine_unit ninexnine_unit_2024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18205)
);

ninexnine_unit ninexnine_unit_2025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19205)
);

ninexnine_unit ninexnine_unit_2026(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A205)
);

ninexnine_unit ninexnine_unit_2027(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B205)
);

ninexnine_unit ninexnine_unit_2028(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C205)
);

ninexnine_unit ninexnine_unit_2029(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D205)
);

ninexnine_unit ninexnine_unit_2030(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E205)
);

ninexnine_unit ninexnine_unit_2031(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F205)
);

assign C1205=c10205+c11205+c12205+c13205+c14205+c15205+c16205+c17205+c18205+c19205+c1A205+c1B205+c1C205+c1D205+c1E205+c1F205;
assign A1205=(C1205>=0)?1:0;

assign P2205=A1205;

ninexnine_unit ninexnine_unit_2032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10215)
);

ninexnine_unit ninexnine_unit_2033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11215)
);

ninexnine_unit ninexnine_unit_2034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12215)
);

ninexnine_unit ninexnine_unit_2035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13215)
);

ninexnine_unit ninexnine_unit_2036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14215)
);

ninexnine_unit ninexnine_unit_2037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15215)
);

ninexnine_unit ninexnine_unit_2038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16215)
);

ninexnine_unit ninexnine_unit_2039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17215)
);

ninexnine_unit ninexnine_unit_2040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18215)
);

ninexnine_unit ninexnine_unit_2041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19215)
);

ninexnine_unit ninexnine_unit_2042(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A215)
);

ninexnine_unit ninexnine_unit_2043(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B215)
);

ninexnine_unit ninexnine_unit_2044(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C215)
);

ninexnine_unit ninexnine_unit_2045(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D215)
);

ninexnine_unit ninexnine_unit_2046(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E215)
);

ninexnine_unit ninexnine_unit_2047(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F215)
);

assign C1215=c10215+c11215+c12215+c13215+c14215+c15215+c16215+c17215+c18215+c19215+c1A215+c1B215+c1C215+c1D215+c1E215+c1F215;
assign A1215=(C1215>=0)?1:0;

assign P2215=A1215;

ninexnine_unit ninexnine_unit_2048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10225)
);

ninexnine_unit ninexnine_unit_2049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11225)
);

ninexnine_unit ninexnine_unit_2050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12225)
);

ninexnine_unit ninexnine_unit_2051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W15003),
				.b1(W15013),
				.b2(W15023),
				.b3(W15103),
				.b4(W15113),
				.b5(W15123),
				.b6(W15203),
				.b7(W15213),
				.b8(W15223),
				.c(c13225)
);

ninexnine_unit ninexnine_unit_2052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W15004),
				.b1(W15014),
				.b2(W15024),
				.b3(W15104),
				.b4(W15114),
				.b5(W15124),
				.b6(W15204),
				.b7(W15214),
				.b8(W15224),
				.c(c14225)
);

ninexnine_unit ninexnine_unit_2053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W15005),
				.b1(W15015),
				.b2(W15025),
				.b3(W15105),
				.b4(W15115),
				.b5(W15125),
				.b6(W15205),
				.b7(W15215),
				.b8(W15225),
				.c(c15225)
);

ninexnine_unit ninexnine_unit_2054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W15006),
				.b1(W15016),
				.b2(W15026),
				.b3(W15106),
				.b4(W15116),
				.b5(W15126),
				.b6(W15206),
				.b7(W15216),
				.b8(W15226),
				.c(c16225)
);

ninexnine_unit ninexnine_unit_2055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W15007),
				.b1(W15017),
				.b2(W15027),
				.b3(W15107),
				.b4(W15117),
				.b5(W15127),
				.b6(W15207),
				.b7(W15217),
				.b8(W15227),
				.c(c17225)
);

ninexnine_unit ninexnine_unit_2056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W15008),
				.b1(W15018),
				.b2(W15028),
				.b3(W15108),
				.b4(W15118),
				.b5(W15128),
				.b6(W15208),
				.b7(W15218),
				.b8(W15228),
				.c(c18225)
);

ninexnine_unit ninexnine_unit_2057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W15009),
				.b1(W15019),
				.b2(W15029),
				.b3(W15109),
				.b4(W15119),
				.b5(W15129),
				.b6(W15209),
				.b7(W15219),
				.b8(W15229),
				.c(c19225)
);

ninexnine_unit ninexnine_unit_2058(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1500A),
				.b1(W1501A),
				.b2(W1502A),
				.b3(W1510A),
				.b4(W1511A),
				.b5(W1512A),
				.b6(W1520A),
				.b7(W1521A),
				.b8(W1522A),
				.c(c1A225)
);

ninexnine_unit ninexnine_unit_2059(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1500B),
				.b1(W1501B),
				.b2(W1502B),
				.b3(W1510B),
				.b4(W1511B),
				.b5(W1512B),
				.b6(W1520B),
				.b7(W1521B),
				.b8(W1522B),
				.c(c1B225)
);

ninexnine_unit ninexnine_unit_2060(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1500C),
				.b1(W1501C),
				.b2(W1502C),
				.b3(W1510C),
				.b4(W1511C),
				.b5(W1512C),
				.b6(W1520C),
				.b7(W1521C),
				.b8(W1522C),
				.c(c1C225)
);

ninexnine_unit ninexnine_unit_2061(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1500D),
				.b1(W1501D),
				.b2(W1502D),
				.b3(W1510D),
				.b4(W1511D),
				.b5(W1512D),
				.b6(W1520D),
				.b7(W1521D),
				.b8(W1522D),
				.c(c1D225)
);

ninexnine_unit ninexnine_unit_2062(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1500E),
				.b1(W1501E),
				.b2(W1502E),
				.b3(W1510E),
				.b4(W1511E),
				.b5(W1512E),
				.b6(W1520E),
				.b7(W1521E),
				.b8(W1522E),
				.c(c1E225)
);

ninexnine_unit ninexnine_unit_2063(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1500F),
				.b1(W1501F),
				.b2(W1502F),
				.b3(W1510F),
				.b4(W1511F),
				.b5(W1512F),
				.b6(W1520F),
				.b7(W1521F),
				.b8(W1522F),
				.c(c1F225)
);

assign C1225=c10225+c11225+c12225+c13225+c14225+c15225+c16225+c17225+c18225+c19225+c1A225+c1B225+c1C225+c1D225+c1E225+c1F225;
assign A1225=(C1225>=0)?1:0;

assign P2225=A1225;

ninexnine_unit ninexnine_unit_2064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10006)
);

ninexnine_unit ninexnine_unit_2065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11006)
);

ninexnine_unit ninexnine_unit_2066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12006)
);

ninexnine_unit ninexnine_unit_2067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13006)
);

ninexnine_unit ninexnine_unit_2068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14006)
);

ninexnine_unit ninexnine_unit_2069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15006)
);

ninexnine_unit ninexnine_unit_2070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16006)
);

ninexnine_unit ninexnine_unit_2071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17006)
);

ninexnine_unit ninexnine_unit_2072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18006)
);

ninexnine_unit ninexnine_unit_2073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19006)
);

ninexnine_unit ninexnine_unit_2074(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A006)
);

ninexnine_unit ninexnine_unit_2075(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B006)
);

ninexnine_unit ninexnine_unit_2076(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C006)
);

ninexnine_unit ninexnine_unit_2077(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D006)
);

ninexnine_unit ninexnine_unit_2078(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E006)
);

ninexnine_unit ninexnine_unit_2079(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F006)
);

assign C1006=c10006+c11006+c12006+c13006+c14006+c15006+c16006+c17006+c18006+c19006+c1A006+c1B006+c1C006+c1D006+c1E006+c1F006;
assign A1006=(C1006>=0)?1:0;

assign P2006=A1006;

ninexnine_unit ninexnine_unit_2080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10016)
);

ninexnine_unit ninexnine_unit_2081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11016)
);

ninexnine_unit ninexnine_unit_2082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12016)
);

ninexnine_unit ninexnine_unit_2083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13016)
);

ninexnine_unit ninexnine_unit_2084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14016)
);

ninexnine_unit ninexnine_unit_2085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15016)
);

ninexnine_unit ninexnine_unit_2086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16016)
);

ninexnine_unit ninexnine_unit_2087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17016)
);

ninexnine_unit ninexnine_unit_2088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18016)
);

ninexnine_unit ninexnine_unit_2089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19016)
);

ninexnine_unit ninexnine_unit_2090(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A016)
);

ninexnine_unit ninexnine_unit_2091(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B016)
);

ninexnine_unit ninexnine_unit_2092(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C016)
);

ninexnine_unit ninexnine_unit_2093(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D016)
);

ninexnine_unit ninexnine_unit_2094(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E016)
);

ninexnine_unit ninexnine_unit_2095(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F016)
);

assign C1016=c10016+c11016+c12016+c13016+c14016+c15016+c16016+c17016+c18016+c19016+c1A016+c1B016+c1C016+c1D016+c1E016+c1F016;
assign A1016=(C1016>=0)?1:0;

assign P2016=A1016;

ninexnine_unit ninexnine_unit_2096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10026)
);

ninexnine_unit ninexnine_unit_2097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11026)
);

ninexnine_unit ninexnine_unit_2098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12026)
);

ninexnine_unit ninexnine_unit_2099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13026)
);

ninexnine_unit ninexnine_unit_2100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14026)
);

ninexnine_unit ninexnine_unit_2101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15026)
);

ninexnine_unit ninexnine_unit_2102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16026)
);

ninexnine_unit ninexnine_unit_2103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17026)
);

ninexnine_unit ninexnine_unit_2104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18026)
);

ninexnine_unit ninexnine_unit_2105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19026)
);

ninexnine_unit ninexnine_unit_2106(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A026)
);

ninexnine_unit ninexnine_unit_2107(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B026)
);

ninexnine_unit ninexnine_unit_2108(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C026)
);

ninexnine_unit ninexnine_unit_2109(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D026)
);

ninexnine_unit ninexnine_unit_2110(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E026)
);

ninexnine_unit ninexnine_unit_2111(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F026)
);

assign C1026=c10026+c11026+c12026+c13026+c14026+c15026+c16026+c17026+c18026+c19026+c1A026+c1B026+c1C026+c1D026+c1E026+c1F026;
assign A1026=(C1026>=0)?1:0;

assign P2026=A1026;

ninexnine_unit ninexnine_unit_2112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10106)
);

ninexnine_unit ninexnine_unit_2113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11106)
);

ninexnine_unit ninexnine_unit_2114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12106)
);

ninexnine_unit ninexnine_unit_2115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13106)
);

ninexnine_unit ninexnine_unit_2116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14106)
);

ninexnine_unit ninexnine_unit_2117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15106)
);

ninexnine_unit ninexnine_unit_2118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16106)
);

ninexnine_unit ninexnine_unit_2119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17106)
);

ninexnine_unit ninexnine_unit_2120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18106)
);

ninexnine_unit ninexnine_unit_2121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19106)
);

ninexnine_unit ninexnine_unit_2122(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A106)
);

ninexnine_unit ninexnine_unit_2123(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B106)
);

ninexnine_unit ninexnine_unit_2124(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C106)
);

ninexnine_unit ninexnine_unit_2125(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D106)
);

ninexnine_unit ninexnine_unit_2126(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E106)
);

ninexnine_unit ninexnine_unit_2127(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F106)
);

assign C1106=c10106+c11106+c12106+c13106+c14106+c15106+c16106+c17106+c18106+c19106+c1A106+c1B106+c1C106+c1D106+c1E106+c1F106;
assign A1106=(C1106>=0)?1:0;

assign P2106=A1106;

ninexnine_unit ninexnine_unit_2128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10116)
);

ninexnine_unit ninexnine_unit_2129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11116)
);

ninexnine_unit ninexnine_unit_2130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12116)
);

ninexnine_unit ninexnine_unit_2131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13116)
);

ninexnine_unit ninexnine_unit_2132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14116)
);

ninexnine_unit ninexnine_unit_2133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15116)
);

ninexnine_unit ninexnine_unit_2134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16116)
);

ninexnine_unit ninexnine_unit_2135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17116)
);

ninexnine_unit ninexnine_unit_2136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18116)
);

ninexnine_unit ninexnine_unit_2137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19116)
);

ninexnine_unit ninexnine_unit_2138(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A116)
);

ninexnine_unit ninexnine_unit_2139(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B116)
);

ninexnine_unit ninexnine_unit_2140(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C116)
);

ninexnine_unit ninexnine_unit_2141(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D116)
);

ninexnine_unit ninexnine_unit_2142(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E116)
);

ninexnine_unit ninexnine_unit_2143(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F116)
);

assign C1116=c10116+c11116+c12116+c13116+c14116+c15116+c16116+c17116+c18116+c19116+c1A116+c1B116+c1C116+c1D116+c1E116+c1F116;
assign A1116=(C1116>=0)?1:0;

assign P2116=A1116;

ninexnine_unit ninexnine_unit_2144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10126)
);

ninexnine_unit ninexnine_unit_2145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11126)
);

ninexnine_unit ninexnine_unit_2146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12126)
);

ninexnine_unit ninexnine_unit_2147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13126)
);

ninexnine_unit ninexnine_unit_2148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14126)
);

ninexnine_unit ninexnine_unit_2149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15126)
);

ninexnine_unit ninexnine_unit_2150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16126)
);

ninexnine_unit ninexnine_unit_2151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17126)
);

ninexnine_unit ninexnine_unit_2152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18126)
);

ninexnine_unit ninexnine_unit_2153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19126)
);

ninexnine_unit ninexnine_unit_2154(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A126)
);

ninexnine_unit ninexnine_unit_2155(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B126)
);

ninexnine_unit ninexnine_unit_2156(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C126)
);

ninexnine_unit ninexnine_unit_2157(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D126)
);

ninexnine_unit ninexnine_unit_2158(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E126)
);

ninexnine_unit ninexnine_unit_2159(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F126)
);

assign C1126=c10126+c11126+c12126+c13126+c14126+c15126+c16126+c17126+c18126+c19126+c1A126+c1B126+c1C126+c1D126+c1E126+c1F126;
assign A1126=(C1126>=0)?1:0;

assign P2126=A1126;

ninexnine_unit ninexnine_unit_2160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10206)
);

ninexnine_unit ninexnine_unit_2161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11206)
);

ninexnine_unit ninexnine_unit_2162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12206)
);

ninexnine_unit ninexnine_unit_2163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13206)
);

ninexnine_unit ninexnine_unit_2164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14206)
);

ninexnine_unit ninexnine_unit_2165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15206)
);

ninexnine_unit ninexnine_unit_2166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16206)
);

ninexnine_unit ninexnine_unit_2167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17206)
);

ninexnine_unit ninexnine_unit_2168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18206)
);

ninexnine_unit ninexnine_unit_2169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19206)
);

ninexnine_unit ninexnine_unit_2170(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A206)
);

ninexnine_unit ninexnine_unit_2171(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B206)
);

ninexnine_unit ninexnine_unit_2172(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C206)
);

ninexnine_unit ninexnine_unit_2173(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D206)
);

ninexnine_unit ninexnine_unit_2174(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E206)
);

ninexnine_unit ninexnine_unit_2175(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F206)
);

assign C1206=c10206+c11206+c12206+c13206+c14206+c15206+c16206+c17206+c18206+c19206+c1A206+c1B206+c1C206+c1D206+c1E206+c1F206;
assign A1206=(C1206>=0)?1:0;

assign P2206=A1206;

ninexnine_unit ninexnine_unit_2176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10216)
);

ninexnine_unit ninexnine_unit_2177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11216)
);

ninexnine_unit ninexnine_unit_2178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12216)
);

ninexnine_unit ninexnine_unit_2179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13216)
);

ninexnine_unit ninexnine_unit_2180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14216)
);

ninexnine_unit ninexnine_unit_2181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15216)
);

ninexnine_unit ninexnine_unit_2182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16216)
);

ninexnine_unit ninexnine_unit_2183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17216)
);

ninexnine_unit ninexnine_unit_2184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18216)
);

ninexnine_unit ninexnine_unit_2185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19216)
);

ninexnine_unit ninexnine_unit_2186(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A216)
);

ninexnine_unit ninexnine_unit_2187(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B216)
);

ninexnine_unit ninexnine_unit_2188(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C216)
);

ninexnine_unit ninexnine_unit_2189(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D216)
);

ninexnine_unit ninexnine_unit_2190(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E216)
);

ninexnine_unit ninexnine_unit_2191(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F216)
);

assign C1216=c10216+c11216+c12216+c13216+c14216+c15216+c16216+c17216+c18216+c19216+c1A216+c1B216+c1C216+c1D216+c1E216+c1F216;
assign A1216=(C1216>=0)?1:0;

assign P2216=A1216;

ninexnine_unit ninexnine_unit_2192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10226)
);

ninexnine_unit ninexnine_unit_2193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11226)
);

ninexnine_unit ninexnine_unit_2194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12226)
);

ninexnine_unit ninexnine_unit_2195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W16003),
				.b1(W16013),
				.b2(W16023),
				.b3(W16103),
				.b4(W16113),
				.b5(W16123),
				.b6(W16203),
				.b7(W16213),
				.b8(W16223),
				.c(c13226)
);

ninexnine_unit ninexnine_unit_2196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W16004),
				.b1(W16014),
				.b2(W16024),
				.b3(W16104),
				.b4(W16114),
				.b5(W16124),
				.b6(W16204),
				.b7(W16214),
				.b8(W16224),
				.c(c14226)
);

ninexnine_unit ninexnine_unit_2197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W16005),
				.b1(W16015),
				.b2(W16025),
				.b3(W16105),
				.b4(W16115),
				.b5(W16125),
				.b6(W16205),
				.b7(W16215),
				.b8(W16225),
				.c(c15226)
);

ninexnine_unit ninexnine_unit_2198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W16006),
				.b1(W16016),
				.b2(W16026),
				.b3(W16106),
				.b4(W16116),
				.b5(W16126),
				.b6(W16206),
				.b7(W16216),
				.b8(W16226),
				.c(c16226)
);

ninexnine_unit ninexnine_unit_2199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W16007),
				.b1(W16017),
				.b2(W16027),
				.b3(W16107),
				.b4(W16117),
				.b5(W16127),
				.b6(W16207),
				.b7(W16217),
				.b8(W16227),
				.c(c17226)
);

ninexnine_unit ninexnine_unit_2200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W16008),
				.b1(W16018),
				.b2(W16028),
				.b3(W16108),
				.b4(W16118),
				.b5(W16128),
				.b6(W16208),
				.b7(W16218),
				.b8(W16228),
				.c(c18226)
);

ninexnine_unit ninexnine_unit_2201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W16009),
				.b1(W16019),
				.b2(W16029),
				.b3(W16109),
				.b4(W16119),
				.b5(W16129),
				.b6(W16209),
				.b7(W16219),
				.b8(W16229),
				.c(c19226)
);

ninexnine_unit ninexnine_unit_2202(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1600A),
				.b1(W1601A),
				.b2(W1602A),
				.b3(W1610A),
				.b4(W1611A),
				.b5(W1612A),
				.b6(W1620A),
				.b7(W1621A),
				.b8(W1622A),
				.c(c1A226)
);

ninexnine_unit ninexnine_unit_2203(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1600B),
				.b1(W1601B),
				.b2(W1602B),
				.b3(W1610B),
				.b4(W1611B),
				.b5(W1612B),
				.b6(W1620B),
				.b7(W1621B),
				.b8(W1622B),
				.c(c1B226)
);

ninexnine_unit ninexnine_unit_2204(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1600C),
				.b1(W1601C),
				.b2(W1602C),
				.b3(W1610C),
				.b4(W1611C),
				.b5(W1612C),
				.b6(W1620C),
				.b7(W1621C),
				.b8(W1622C),
				.c(c1C226)
);

ninexnine_unit ninexnine_unit_2205(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1600D),
				.b1(W1601D),
				.b2(W1602D),
				.b3(W1610D),
				.b4(W1611D),
				.b5(W1612D),
				.b6(W1620D),
				.b7(W1621D),
				.b8(W1622D),
				.c(c1D226)
);

ninexnine_unit ninexnine_unit_2206(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1600E),
				.b1(W1601E),
				.b2(W1602E),
				.b3(W1610E),
				.b4(W1611E),
				.b5(W1612E),
				.b6(W1620E),
				.b7(W1621E),
				.b8(W1622E),
				.c(c1E226)
);

ninexnine_unit ninexnine_unit_2207(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1600F),
				.b1(W1601F),
				.b2(W1602F),
				.b3(W1610F),
				.b4(W1611F),
				.b5(W1612F),
				.b6(W1620F),
				.b7(W1621F),
				.b8(W1622F),
				.c(c1F226)
);

assign C1226=c10226+c11226+c12226+c13226+c14226+c15226+c16226+c17226+c18226+c19226+c1A226+c1B226+c1C226+c1D226+c1E226+c1F226;
assign A1226=(C1226>=0)?1:0;

assign P2226=A1226;

ninexnine_unit ninexnine_unit_2208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10007)
);

ninexnine_unit ninexnine_unit_2209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11007)
);

ninexnine_unit ninexnine_unit_2210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12007)
);

ninexnine_unit ninexnine_unit_2211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13007)
);

ninexnine_unit ninexnine_unit_2212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14007)
);

ninexnine_unit ninexnine_unit_2213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15007)
);

ninexnine_unit ninexnine_unit_2214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16007)
);

ninexnine_unit ninexnine_unit_2215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17007)
);

ninexnine_unit ninexnine_unit_2216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18007)
);

ninexnine_unit ninexnine_unit_2217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19007)
);

ninexnine_unit ninexnine_unit_2218(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A007)
);

ninexnine_unit ninexnine_unit_2219(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B007)
);

ninexnine_unit ninexnine_unit_2220(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C007)
);

ninexnine_unit ninexnine_unit_2221(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D007)
);

ninexnine_unit ninexnine_unit_2222(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E007)
);

ninexnine_unit ninexnine_unit_2223(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F007)
);

assign C1007=c10007+c11007+c12007+c13007+c14007+c15007+c16007+c17007+c18007+c19007+c1A007+c1B007+c1C007+c1D007+c1E007+c1F007;
assign A1007=(C1007>=0)?1:0;

assign P2007=A1007;

ninexnine_unit ninexnine_unit_2224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10017)
);

ninexnine_unit ninexnine_unit_2225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11017)
);

ninexnine_unit ninexnine_unit_2226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12017)
);

ninexnine_unit ninexnine_unit_2227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13017)
);

ninexnine_unit ninexnine_unit_2228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14017)
);

ninexnine_unit ninexnine_unit_2229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15017)
);

ninexnine_unit ninexnine_unit_2230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16017)
);

ninexnine_unit ninexnine_unit_2231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17017)
);

ninexnine_unit ninexnine_unit_2232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18017)
);

ninexnine_unit ninexnine_unit_2233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19017)
);

ninexnine_unit ninexnine_unit_2234(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A017)
);

ninexnine_unit ninexnine_unit_2235(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B017)
);

ninexnine_unit ninexnine_unit_2236(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C017)
);

ninexnine_unit ninexnine_unit_2237(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D017)
);

ninexnine_unit ninexnine_unit_2238(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E017)
);

ninexnine_unit ninexnine_unit_2239(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F017)
);

assign C1017=c10017+c11017+c12017+c13017+c14017+c15017+c16017+c17017+c18017+c19017+c1A017+c1B017+c1C017+c1D017+c1E017+c1F017;
assign A1017=(C1017>=0)?1:0;

assign P2017=A1017;

ninexnine_unit ninexnine_unit_2240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10027)
);

ninexnine_unit ninexnine_unit_2241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11027)
);

ninexnine_unit ninexnine_unit_2242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12027)
);

ninexnine_unit ninexnine_unit_2243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13027)
);

ninexnine_unit ninexnine_unit_2244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14027)
);

ninexnine_unit ninexnine_unit_2245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15027)
);

ninexnine_unit ninexnine_unit_2246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16027)
);

ninexnine_unit ninexnine_unit_2247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17027)
);

ninexnine_unit ninexnine_unit_2248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18027)
);

ninexnine_unit ninexnine_unit_2249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19027)
);

ninexnine_unit ninexnine_unit_2250(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A027)
);

ninexnine_unit ninexnine_unit_2251(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B027)
);

ninexnine_unit ninexnine_unit_2252(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C027)
);

ninexnine_unit ninexnine_unit_2253(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D027)
);

ninexnine_unit ninexnine_unit_2254(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E027)
);

ninexnine_unit ninexnine_unit_2255(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F027)
);

assign C1027=c10027+c11027+c12027+c13027+c14027+c15027+c16027+c17027+c18027+c19027+c1A027+c1B027+c1C027+c1D027+c1E027+c1F027;
assign A1027=(C1027>=0)?1:0;

assign P2027=A1027;

ninexnine_unit ninexnine_unit_2256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10107)
);

ninexnine_unit ninexnine_unit_2257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11107)
);

ninexnine_unit ninexnine_unit_2258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12107)
);

ninexnine_unit ninexnine_unit_2259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13107)
);

ninexnine_unit ninexnine_unit_2260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14107)
);

ninexnine_unit ninexnine_unit_2261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15107)
);

ninexnine_unit ninexnine_unit_2262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16107)
);

ninexnine_unit ninexnine_unit_2263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17107)
);

ninexnine_unit ninexnine_unit_2264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18107)
);

ninexnine_unit ninexnine_unit_2265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19107)
);

ninexnine_unit ninexnine_unit_2266(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A107)
);

ninexnine_unit ninexnine_unit_2267(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B107)
);

ninexnine_unit ninexnine_unit_2268(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C107)
);

ninexnine_unit ninexnine_unit_2269(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D107)
);

ninexnine_unit ninexnine_unit_2270(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E107)
);

ninexnine_unit ninexnine_unit_2271(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F107)
);

assign C1107=c10107+c11107+c12107+c13107+c14107+c15107+c16107+c17107+c18107+c19107+c1A107+c1B107+c1C107+c1D107+c1E107+c1F107;
assign A1107=(C1107>=0)?1:0;

assign P2107=A1107;

ninexnine_unit ninexnine_unit_2272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10117)
);

ninexnine_unit ninexnine_unit_2273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11117)
);

ninexnine_unit ninexnine_unit_2274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12117)
);

ninexnine_unit ninexnine_unit_2275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13117)
);

ninexnine_unit ninexnine_unit_2276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14117)
);

ninexnine_unit ninexnine_unit_2277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15117)
);

ninexnine_unit ninexnine_unit_2278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16117)
);

ninexnine_unit ninexnine_unit_2279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17117)
);

ninexnine_unit ninexnine_unit_2280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18117)
);

ninexnine_unit ninexnine_unit_2281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19117)
);

ninexnine_unit ninexnine_unit_2282(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A117)
);

ninexnine_unit ninexnine_unit_2283(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B117)
);

ninexnine_unit ninexnine_unit_2284(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C117)
);

ninexnine_unit ninexnine_unit_2285(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D117)
);

ninexnine_unit ninexnine_unit_2286(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E117)
);

ninexnine_unit ninexnine_unit_2287(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F117)
);

assign C1117=c10117+c11117+c12117+c13117+c14117+c15117+c16117+c17117+c18117+c19117+c1A117+c1B117+c1C117+c1D117+c1E117+c1F117;
assign A1117=(C1117>=0)?1:0;

assign P2117=A1117;

ninexnine_unit ninexnine_unit_2288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10127)
);

ninexnine_unit ninexnine_unit_2289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11127)
);

ninexnine_unit ninexnine_unit_2290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12127)
);

ninexnine_unit ninexnine_unit_2291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13127)
);

ninexnine_unit ninexnine_unit_2292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14127)
);

ninexnine_unit ninexnine_unit_2293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15127)
);

ninexnine_unit ninexnine_unit_2294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16127)
);

ninexnine_unit ninexnine_unit_2295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17127)
);

ninexnine_unit ninexnine_unit_2296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18127)
);

ninexnine_unit ninexnine_unit_2297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19127)
);

ninexnine_unit ninexnine_unit_2298(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A127)
);

ninexnine_unit ninexnine_unit_2299(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B127)
);

ninexnine_unit ninexnine_unit_2300(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C127)
);

ninexnine_unit ninexnine_unit_2301(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D127)
);

ninexnine_unit ninexnine_unit_2302(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E127)
);

ninexnine_unit ninexnine_unit_2303(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F127)
);

assign C1127=c10127+c11127+c12127+c13127+c14127+c15127+c16127+c17127+c18127+c19127+c1A127+c1B127+c1C127+c1D127+c1E127+c1F127;
assign A1127=(C1127>=0)?1:0;

assign P2127=A1127;

ninexnine_unit ninexnine_unit_2304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10207)
);

ninexnine_unit ninexnine_unit_2305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11207)
);

ninexnine_unit ninexnine_unit_2306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12207)
);

ninexnine_unit ninexnine_unit_2307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13207)
);

ninexnine_unit ninexnine_unit_2308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14207)
);

ninexnine_unit ninexnine_unit_2309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15207)
);

ninexnine_unit ninexnine_unit_2310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16207)
);

ninexnine_unit ninexnine_unit_2311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17207)
);

ninexnine_unit ninexnine_unit_2312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18207)
);

ninexnine_unit ninexnine_unit_2313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19207)
);

ninexnine_unit ninexnine_unit_2314(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A207)
);

ninexnine_unit ninexnine_unit_2315(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B207)
);

ninexnine_unit ninexnine_unit_2316(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C207)
);

ninexnine_unit ninexnine_unit_2317(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D207)
);

ninexnine_unit ninexnine_unit_2318(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E207)
);

ninexnine_unit ninexnine_unit_2319(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F207)
);

assign C1207=c10207+c11207+c12207+c13207+c14207+c15207+c16207+c17207+c18207+c19207+c1A207+c1B207+c1C207+c1D207+c1E207+c1F207;
assign A1207=(C1207>=0)?1:0;

assign P2207=A1207;

ninexnine_unit ninexnine_unit_2320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10217)
);

ninexnine_unit ninexnine_unit_2321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11217)
);

ninexnine_unit ninexnine_unit_2322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12217)
);

ninexnine_unit ninexnine_unit_2323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13217)
);

ninexnine_unit ninexnine_unit_2324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14217)
);

ninexnine_unit ninexnine_unit_2325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15217)
);

ninexnine_unit ninexnine_unit_2326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16217)
);

ninexnine_unit ninexnine_unit_2327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17217)
);

ninexnine_unit ninexnine_unit_2328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18217)
);

ninexnine_unit ninexnine_unit_2329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19217)
);

ninexnine_unit ninexnine_unit_2330(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A217)
);

ninexnine_unit ninexnine_unit_2331(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B217)
);

ninexnine_unit ninexnine_unit_2332(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C217)
);

ninexnine_unit ninexnine_unit_2333(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D217)
);

ninexnine_unit ninexnine_unit_2334(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E217)
);

ninexnine_unit ninexnine_unit_2335(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F217)
);

assign C1217=c10217+c11217+c12217+c13217+c14217+c15217+c16217+c17217+c18217+c19217+c1A217+c1B217+c1C217+c1D217+c1E217+c1F217;
assign A1217=(C1217>=0)?1:0;

assign P2217=A1217;

ninexnine_unit ninexnine_unit_2336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10227)
);

ninexnine_unit ninexnine_unit_2337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11227)
);

ninexnine_unit ninexnine_unit_2338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12227)
);

ninexnine_unit ninexnine_unit_2339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W17003),
				.b1(W17013),
				.b2(W17023),
				.b3(W17103),
				.b4(W17113),
				.b5(W17123),
				.b6(W17203),
				.b7(W17213),
				.b8(W17223),
				.c(c13227)
);

ninexnine_unit ninexnine_unit_2340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W17004),
				.b1(W17014),
				.b2(W17024),
				.b3(W17104),
				.b4(W17114),
				.b5(W17124),
				.b6(W17204),
				.b7(W17214),
				.b8(W17224),
				.c(c14227)
);

ninexnine_unit ninexnine_unit_2341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W17005),
				.b1(W17015),
				.b2(W17025),
				.b3(W17105),
				.b4(W17115),
				.b5(W17125),
				.b6(W17205),
				.b7(W17215),
				.b8(W17225),
				.c(c15227)
);

ninexnine_unit ninexnine_unit_2342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W17006),
				.b1(W17016),
				.b2(W17026),
				.b3(W17106),
				.b4(W17116),
				.b5(W17126),
				.b6(W17206),
				.b7(W17216),
				.b8(W17226),
				.c(c16227)
);

ninexnine_unit ninexnine_unit_2343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W17007),
				.b1(W17017),
				.b2(W17027),
				.b3(W17107),
				.b4(W17117),
				.b5(W17127),
				.b6(W17207),
				.b7(W17217),
				.b8(W17227),
				.c(c17227)
);

ninexnine_unit ninexnine_unit_2344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W17008),
				.b1(W17018),
				.b2(W17028),
				.b3(W17108),
				.b4(W17118),
				.b5(W17128),
				.b6(W17208),
				.b7(W17218),
				.b8(W17228),
				.c(c18227)
);

ninexnine_unit ninexnine_unit_2345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W17009),
				.b1(W17019),
				.b2(W17029),
				.b3(W17109),
				.b4(W17119),
				.b5(W17129),
				.b6(W17209),
				.b7(W17219),
				.b8(W17229),
				.c(c19227)
);

ninexnine_unit ninexnine_unit_2346(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1700A),
				.b1(W1701A),
				.b2(W1702A),
				.b3(W1710A),
				.b4(W1711A),
				.b5(W1712A),
				.b6(W1720A),
				.b7(W1721A),
				.b8(W1722A),
				.c(c1A227)
);

ninexnine_unit ninexnine_unit_2347(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1700B),
				.b1(W1701B),
				.b2(W1702B),
				.b3(W1710B),
				.b4(W1711B),
				.b5(W1712B),
				.b6(W1720B),
				.b7(W1721B),
				.b8(W1722B),
				.c(c1B227)
);

ninexnine_unit ninexnine_unit_2348(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1700C),
				.b1(W1701C),
				.b2(W1702C),
				.b3(W1710C),
				.b4(W1711C),
				.b5(W1712C),
				.b6(W1720C),
				.b7(W1721C),
				.b8(W1722C),
				.c(c1C227)
);

ninexnine_unit ninexnine_unit_2349(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1700D),
				.b1(W1701D),
				.b2(W1702D),
				.b3(W1710D),
				.b4(W1711D),
				.b5(W1712D),
				.b6(W1720D),
				.b7(W1721D),
				.b8(W1722D),
				.c(c1D227)
);

ninexnine_unit ninexnine_unit_2350(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1700E),
				.b1(W1701E),
				.b2(W1702E),
				.b3(W1710E),
				.b4(W1711E),
				.b5(W1712E),
				.b6(W1720E),
				.b7(W1721E),
				.b8(W1722E),
				.c(c1E227)
);

ninexnine_unit ninexnine_unit_2351(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1700F),
				.b1(W1701F),
				.b2(W1702F),
				.b3(W1710F),
				.b4(W1711F),
				.b5(W1712F),
				.b6(W1720F),
				.b7(W1721F),
				.b8(W1722F),
				.c(c1F227)
);

assign C1227=c10227+c11227+c12227+c13227+c14227+c15227+c16227+c17227+c18227+c19227+c1A227+c1B227+c1C227+c1D227+c1E227+c1F227;
assign A1227=(C1227>=0)?1:0;

assign P2227=A1227;

ninexnine_unit ninexnine_unit_2352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10008)
);

ninexnine_unit ninexnine_unit_2353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11008)
);

ninexnine_unit ninexnine_unit_2354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12008)
);

ninexnine_unit ninexnine_unit_2355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13008)
);

ninexnine_unit ninexnine_unit_2356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14008)
);

ninexnine_unit ninexnine_unit_2357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15008)
);

ninexnine_unit ninexnine_unit_2358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16008)
);

ninexnine_unit ninexnine_unit_2359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17008)
);

ninexnine_unit ninexnine_unit_2360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18008)
);

ninexnine_unit ninexnine_unit_2361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19008)
);

ninexnine_unit ninexnine_unit_2362(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A008)
);

ninexnine_unit ninexnine_unit_2363(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B008)
);

ninexnine_unit ninexnine_unit_2364(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C008)
);

ninexnine_unit ninexnine_unit_2365(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D008)
);

ninexnine_unit ninexnine_unit_2366(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E008)
);

ninexnine_unit ninexnine_unit_2367(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F008)
);

assign C1008=c10008+c11008+c12008+c13008+c14008+c15008+c16008+c17008+c18008+c19008+c1A008+c1B008+c1C008+c1D008+c1E008+c1F008;
assign A1008=(C1008>=0)?1:0;

assign P2008=A1008;

ninexnine_unit ninexnine_unit_2368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10018)
);

ninexnine_unit ninexnine_unit_2369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11018)
);

ninexnine_unit ninexnine_unit_2370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12018)
);

ninexnine_unit ninexnine_unit_2371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13018)
);

ninexnine_unit ninexnine_unit_2372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14018)
);

ninexnine_unit ninexnine_unit_2373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15018)
);

ninexnine_unit ninexnine_unit_2374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16018)
);

ninexnine_unit ninexnine_unit_2375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17018)
);

ninexnine_unit ninexnine_unit_2376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18018)
);

ninexnine_unit ninexnine_unit_2377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19018)
);

ninexnine_unit ninexnine_unit_2378(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A018)
);

ninexnine_unit ninexnine_unit_2379(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B018)
);

ninexnine_unit ninexnine_unit_2380(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C018)
);

ninexnine_unit ninexnine_unit_2381(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D018)
);

ninexnine_unit ninexnine_unit_2382(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E018)
);

ninexnine_unit ninexnine_unit_2383(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F018)
);

assign C1018=c10018+c11018+c12018+c13018+c14018+c15018+c16018+c17018+c18018+c19018+c1A018+c1B018+c1C018+c1D018+c1E018+c1F018;
assign A1018=(C1018>=0)?1:0;

assign P2018=A1018;

ninexnine_unit ninexnine_unit_2384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10028)
);

ninexnine_unit ninexnine_unit_2385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11028)
);

ninexnine_unit ninexnine_unit_2386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12028)
);

ninexnine_unit ninexnine_unit_2387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13028)
);

ninexnine_unit ninexnine_unit_2388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14028)
);

ninexnine_unit ninexnine_unit_2389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15028)
);

ninexnine_unit ninexnine_unit_2390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16028)
);

ninexnine_unit ninexnine_unit_2391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17028)
);

ninexnine_unit ninexnine_unit_2392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18028)
);

ninexnine_unit ninexnine_unit_2393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19028)
);

ninexnine_unit ninexnine_unit_2394(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A028)
);

ninexnine_unit ninexnine_unit_2395(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B028)
);

ninexnine_unit ninexnine_unit_2396(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C028)
);

ninexnine_unit ninexnine_unit_2397(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D028)
);

ninexnine_unit ninexnine_unit_2398(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E028)
);

ninexnine_unit ninexnine_unit_2399(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F028)
);

assign C1028=c10028+c11028+c12028+c13028+c14028+c15028+c16028+c17028+c18028+c19028+c1A028+c1B028+c1C028+c1D028+c1E028+c1F028;
assign A1028=(C1028>=0)?1:0;

assign P2028=A1028;

ninexnine_unit ninexnine_unit_2400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10108)
);

ninexnine_unit ninexnine_unit_2401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11108)
);

ninexnine_unit ninexnine_unit_2402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12108)
);

ninexnine_unit ninexnine_unit_2403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13108)
);

ninexnine_unit ninexnine_unit_2404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14108)
);

ninexnine_unit ninexnine_unit_2405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15108)
);

ninexnine_unit ninexnine_unit_2406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16108)
);

ninexnine_unit ninexnine_unit_2407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17108)
);

ninexnine_unit ninexnine_unit_2408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18108)
);

ninexnine_unit ninexnine_unit_2409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19108)
);

ninexnine_unit ninexnine_unit_2410(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A108)
);

ninexnine_unit ninexnine_unit_2411(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B108)
);

ninexnine_unit ninexnine_unit_2412(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C108)
);

ninexnine_unit ninexnine_unit_2413(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D108)
);

ninexnine_unit ninexnine_unit_2414(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E108)
);

ninexnine_unit ninexnine_unit_2415(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F108)
);

assign C1108=c10108+c11108+c12108+c13108+c14108+c15108+c16108+c17108+c18108+c19108+c1A108+c1B108+c1C108+c1D108+c1E108+c1F108;
assign A1108=(C1108>=0)?1:0;

assign P2108=A1108;

ninexnine_unit ninexnine_unit_2416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10118)
);

ninexnine_unit ninexnine_unit_2417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11118)
);

ninexnine_unit ninexnine_unit_2418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12118)
);

ninexnine_unit ninexnine_unit_2419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13118)
);

ninexnine_unit ninexnine_unit_2420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14118)
);

ninexnine_unit ninexnine_unit_2421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15118)
);

ninexnine_unit ninexnine_unit_2422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16118)
);

ninexnine_unit ninexnine_unit_2423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17118)
);

ninexnine_unit ninexnine_unit_2424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18118)
);

ninexnine_unit ninexnine_unit_2425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19118)
);

ninexnine_unit ninexnine_unit_2426(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A118)
);

ninexnine_unit ninexnine_unit_2427(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B118)
);

ninexnine_unit ninexnine_unit_2428(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C118)
);

ninexnine_unit ninexnine_unit_2429(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D118)
);

ninexnine_unit ninexnine_unit_2430(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E118)
);

ninexnine_unit ninexnine_unit_2431(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F118)
);

assign C1118=c10118+c11118+c12118+c13118+c14118+c15118+c16118+c17118+c18118+c19118+c1A118+c1B118+c1C118+c1D118+c1E118+c1F118;
assign A1118=(C1118>=0)?1:0;

assign P2118=A1118;

ninexnine_unit ninexnine_unit_2432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10128)
);

ninexnine_unit ninexnine_unit_2433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11128)
);

ninexnine_unit ninexnine_unit_2434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12128)
);

ninexnine_unit ninexnine_unit_2435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13128)
);

ninexnine_unit ninexnine_unit_2436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14128)
);

ninexnine_unit ninexnine_unit_2437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15128)
);

ninexnine_unit ninexnine_unit_2438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16128)
);

ninexnine_unit ninexnine_unit_2439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17128)
);

ninexnine_unit ninexnine_unit_2440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18128)
);

ninexnine_unit ninexnine_unit_2441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19128)
);

ninexnine_unit ninexnine_unit_2442(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A128)
);

ninexnine_unit ninexnine_unit_2443(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B128)
);

ninexnine_unit ninexnine_unit_2444(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C128)
);

ninexnine_unit ninexnine_unit_2445(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D128)
);

ninexnine_unit ninexnine_unit_2446(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E128)
);

ninexnine_unit ninexnine_unit_2447(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F128)
);

assign C1128=c10128+c11128+c12128+c13128+c14128+c15128+c16128+c17128+c18128+c19128+c1A128+c1B128+c1C128+c1D128+c1E128+c1F128;
assign A1128=(C1128>=0)?1:0;

assign P2128=A1128;

ninexnine_unit ninexnine_unit_2448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10208)
);

ninexnine_unit ninexnine_unit_2449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11208)
);

ninexnine_unit ninexnine_unit_2450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12208)
);

ninexnine_unit ninexnine_unit_2451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13208)
);

ninexnine_unit ninexnine_unit_2452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14208)
);

ninexnine_unit ninexnine_unit_2453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15208)
);

ninexnine_unit ninexnine_unit_2454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16208)
);

ninexnine_unit ninexnine_unit_2455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17208)
);

ninexnine_unit ninexnine_unit_2456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18208)
);

ninexnine_unit ninexnine_unit_2457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19208)
);

ninexnine_unit ninexnine_unit_2458(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A208)
);

ninexnine_unit ninexnine_unit_2459(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B208)
);

ninexnine_unit ninexnine_unit_2460(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C208)
);

ninexnine_unit ninexnine_unit_2461(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D208)
);

ninexnine_unit ninexnine_unit_2462(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E208)
);

ninexnine_unit ninexnine_unit_2463(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F208)
);

assign C1208=c10208+c11208+c12208+c13208+c14208+c15208+c16208+c17208+c18208+c19208+c1A208+c1B208+c1C208+c1D208+c1E208+c1F208;
assign A1208=(C1208>=0)?1:0;

assign P2208=A1208;

ninexnine_unit ninexnine_unit_2464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10218)
);

ninexnine_unit ninexnine_unit_2465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11218)
);

ninexnine_unit ninexnine_unit_2466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12218)
);

ninexnine_unit ninexnine_unit_2467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13218)
);

ninexnine_unit ninexnine_unit_2468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14218)
);

ninexnine_unit ninexnine_unit_2469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15218)
);

ninexnine_unit ninexnine_unit_2470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16218)
);

ninexnine_unit ninexnine_unit_2471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17218)
);

ninexnine_unit ninexnine_unit_2472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18218)
);

ninexnine_unit ninexnine_unit_2473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19218)
);

ninexnine_unit ninexnine_unit_2474(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A218)
);

ninexnine_unit ninexnine_unit_2475(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B218)
);

ninexnine_unit ninexnine_unit_2476(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C218)
);

ninexnine_unit ninexnine_unit_2477(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D218)
);

ninexnine_unit ninexnine_unit_2478(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E218)
);

ninexnine_unit ninexnine_unit_2479(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F218)
);

assign C1218=c10218+c11218+c12218+c13218+c14218+c15218+c16218+c17218+c18218+c19218+c1A218+c1B218+c1C218+c1D218+c1E218+c1F218;
assign A1218=(C1218>=0)?1:0;

assign P2218=A1218;

ninexnine_unit ninexnine_unit_2480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10228)
);

ninexnine_unit ninexnine_unit_2481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11228)
);

ninexnine_unit ninexnine_unit_2482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12228)
);

ninexnine_unit ninexnine_unit_2483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W18003),
				.b1(W18013),
				.b2(W18023),
				.b3(W18103),
				.b4(W18113),
				.b5(W18123),
				.b6(W18203),
				.b7(W18213),
				.b8(W18223),
				.c(c13228)
);

ninexnine_unit ninexnine_unit_2484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W18004),
				.b1(W18014),
				.b2(W18024),
				.b3(W18104),
				.b4(W18114),
				.b5(W18124),
				.b6(W18204),
				.b7(W18214),
				.b8(W18224),
				.c(c14228)
);

ninexnine_unit ninexnine_unit_2485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W18005),
				.b1(W18015),
				.b2(W18025),
				.b3(W18105),
				.b4(W18115),
				.b5(W18125),
				.b6(W18205),
				.b7(W18215),
				.b8(W18225),
				.c(c15228)
);

ninexnine_unit ninexnine_unit_2486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W18006),
				.b1(W18016),
				.b2(W18026),
				.b3(W18106),
				.b4(W18116),
				.b5(W18126),
				.b6(W18206),
				.b7(W18216),
				.b8(W18226),
				.c(c16228)
);

ninexnine_unit ninexnine_unit_2487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W18007),
				.b1(W18017),
				.b2(W18027),
				.b3(W18107),
				.b4(W18117),
				.b5(W18127),
				.b6(W18207),
				.b7(W18217),
				.b8(W18227),
				.c(c17228)
);

ninexnine_unit ninexnine_unit_2488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W18008),
				.b1(W18018),
				.b2(W18028),
				.b3(W18108),
				.b4(W18118),
				.b5(W18128),
				.b6(W18208),
				.b7(W18218),
				.b8(W18228),
				.c(c18228)
);

ninexnine_unit ninexnine_unit_2489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W18009),
				.b1(W18019),
				.b2(W18029),
				.b3(W18109),
				.b4(W18119),
				.b5(W18129),
				.b6(W18209),
				.b7(W18219),
				.b8(W18229),
				.c(c19228)
);

ninexnine_unit ninexnine_unit_2490(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1800A),
				.b1(W1801A),
				.b2(W1802A),
				.b3(W1810A),
				.b4(W1811A),
				.b5(W1812A),
				.b6(W1820A),
				.b7(W1821A),
				.b8(W1822A),
				.c(c1A228)
);

ninexnine_unit ninexnine_unit_2491(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1800B),
				.b1(W1801B),
				.b2(W1802B),
				.b3(W1810B),
				.b4(W1811B),
				.b5(W1812B),
				.b6(W1820B),
				.b7(W1821B),
				.b8(W1822B),
				.c(c1B228)
);

ninexnine_unit ninexnine_unit_2492(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1800C),
				.b1(W1801C),
				.b2(W1802C),
				.b3(W1810C),
				.b4(W1811C),
				.b5(W1812C),
				.b6(W1820C),
				.b7(W1821C),
				.b8(W1822C),
				.c(c1C228)
);

ninexnine_unit ninexnine_unit_2493(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1800D),
				.b1(W1801D),
				.b2(W1802D),
				.b3(W1810D),
				.b4(W1811D),
				.b5(W1812D),
				.b6(W1820D),
				.b7(W1821D),
				.b8(W1822D),
				.c(c1D228)
);

ninexnine_unit ninexnine_unit_2494(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1800E),
				.b1(W1801E),
				.b2(W1802E),
				.b3(W1810E),
				.b4(W1811E),
				.b5(W1812E),
				.b6(W1820E),
				.b7(W1821E),
				.b8(W1822E),
				.c(c1E228)
);

ninexnine_unit ninexnine_unit_2495(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1800F),
				.b1(W1801F),
				.b2(W1802F),
				.b3(W1810F),
				.b4(W1811F),
				.b5(W1812F),
				.b6(W1820F),
				.b7(W1821F),
				.b8(W1822F),
				.c(c1F228)
);

assign C1228=c10228+c11228+c12228+c13228+c14228+c15228+c16228+c17228+c18228+c19228+c1A228+c1B228+c1C228+c1D228+c1E228+c1F228;
assign A1228=(C1228>=0)?1:0;

assign P2228=A1228;

ninexnine_unit ninexnine_unit_2496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10009)
);

ninexnine_unit ninexnine_unit_2497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11009)
);

ninexnine_unit ninexnine_unit_2498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12009)
);

ninexnine_unit ninexnine_unit_2499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13009)
);

ninexnine_unit ninexnine_unit_2500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14009)
);

ninexnine_unit ninexnine_unit_2501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15009)
);

ninexnine_unit ninexnine_unit_2502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16009)
);

ninexnine_unit ninexnine_unit_2503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17009)
);

ninexnine_unit ninexnine_unit_2504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18009)
);

ninexnine_unit ninexnine_unit_2505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19009)
);

ninexnine_unit ninexnine_unit_2506(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A009)
);

ninexnine_unit ninexnine_unit_2507(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B009)
);

ninexnine_unit ninexnine_unit_2508(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C009)
);

ninexnine_unit ninexnine_unit_2509(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D009)
);

ninexnine_unit ninexnine_unit_2510(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E009)
);

ninexnine_unit ninexnine_unit_2511(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F009)
);

assign C1009=c10009+c11009+c12009+c13009+c14009+c15009+c16009+c17009+c18009+c19009+c1A009+c1B009+c1C009+c1D009+c1E009+c1F009;
assign A1009=(C1009>=0)?1:0;

assign P2009=A1009;

ninexnine_unit ninexnine_unit_2512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10019)
);

ninexnine_unit ninexnine_unit_2513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11019)
);

ninexnine_unit ninexnine_unit_2514(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12019)
);

ninexnine_unit ninexnine_unit_2515(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13019)
);

ninexnine_unit ninexnine_unit_2516(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14019)
);

ninexnine_unit ninexnine_unit_2517(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15019)
);

ninexnine_unit ninexnine_unit_2518(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16019)
);

ninexnine_unit ninexnine_unit_2519(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17019)
);

ninexnine_unit ninexnine_unit_2520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18019)
);

ninexnine_unit ninexnine_unit_2521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19019)
);

ninexnine_unit ninexnine_unit_2522(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A019)
);

ninexnine_unit ninexnine_unit_2523(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B019)
);

ninexnine_unit ninexnine_unit_2524(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C019)
);

ninexnine_unit ninexnine_unit_2525(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D019)
);

ninexnine_unit ninexnine_unit_2526(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E019)
);

ninexnine_unit ninexnine_unit_2527(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F019)
);

assign C1019=c10019+c11019+c12019+c13019+c14019+c15019+c16019+c17019+c18019+c19019+c1A019+c1B019+c1C019+c1D019+c1E019+c1F019;
assign A1019=(C1019>=0)?1:0;

assign P2019=A1019;

ninexnine_unit ninexnine_unit_2528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10029)
);

ninexnine_unit ninexnine_unit_2529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11029)
);

ninexnine_unit ninexnine_unit_2530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12029)
);

ninexnine_unit ninexnine_unit_2531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13029)
);

ninexnine_unit ninexnine_unit_2532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14029)
);

ninexnine_unit ninexnine_unit_2533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15029)
);

ninexnine_unit ninexnine_unit_2534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16029)
);

ninexnine_unit ninexnine_unit_2535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17029)
);

ninexnine_unit ninexnine_unit_2536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18029)
);

ninexnine_unit ninexnine_unit_2537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19029)
);

ninexnine_unit ninexnine_unit_2538(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A029)
);

ninexnine_unit ninexnine_unit_2539(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B029)
);

ninexnine_unit ninexnine_unit_2540(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C029)
);

ninexnine_unit ninexnine_unit_2541(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D029)
);

ninexnine_unit ninexnine_unit_2542(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E029)
);

ninexnine_unit ninexnine_unit_2543(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F029)
);

assign C1029=c10029+c11029+c12029+c13029+c14029+c15029+c16029+c17029+c18029+c19029+c1A029+c1B029+c1C029+c1D029+c1E029+c1F029;
assign A1029=(C1029>=0)?1:0;

assign P2029=A1029;

ninexnine_unit ninexnine_unit_2544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10109)
);

ninexnine_unit ninexnine_unit_2545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11109)
);

ninexnine_unit ninexnine_unit_2546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12109)
);

ninexnine_unit ninexnine_unit_2547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13109)
);

ninexnine_unit ninexnine_unit_2548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14109)
);

ninexnine_unit ninexnine_unit_2549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15109)
);

ninexnine_unit ninexnine_unit_2550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16109)
);

ninexnine_unit ninexnine_unit_2551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17109)
);

ninexnine_unit ninexnine_unit_2552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18109)
);

ninexnine_unit ninexnine_unit_2553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19109)
);

ninexnine_unit ninexnine_unit_2554(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A109)
);

ninexnine_unit ninexnine_unit_2555(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B109)
);

ninexnine_unit ninexnine_unit_2556(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C109)
);

ninexnine_unit ninexnine_unit_2557(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D109)
);

ninexnine_unit ninexnine_unit_2558(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E109)
);

ninexnine_unit ninexnine_unit_2559(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F109)
);

assign C1109=c10109+c11109+c12109+c13109+c14109+c15109+c16109+c17109+c18109+c19109+c1A109+c1B109+c1C109+c1D109+c1E109+c1F109;
assign A1109=(C1109>=0)?1:0;

assign P2109=A1109;

ninexnine_unit ninexnine_unit_2560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10119)
);

ninexnine_unit ninexnine_unit_2561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11119)
);

ninexnine_unit ninexnine_unit_2562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12119)
);

ninexnine_unit ninexnine_unit_2563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13119)
);

ninexnine_unit ninexnine_unit_2564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14119)
);

ninexnine_unit ninexnine_unit_2565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15119)
);

ninexnine_unit ninexnine_unit_2566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16119)
);

ninexnine_unit ninexnine_unit_2567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17119)
);

ninexnine_unit ninexnine_unit_2568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18119)
);

ninexnine_unit ninexnine_unit_2569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19119)
);

ninexnine_unit ninexnine_unit_2570(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A119)
);

ninexnine_unit ninexnine_unit_2571(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B119)
);

ninexnine_unit ninexnine_unit_2572(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C119)
);

ninexnine_unit ninexnine_unit_2573(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D119)
);

ninexnine_unit ninexnine_unit_2574(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E119)
);

ninexnine_unit ninexnine_unit_2575(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F119)
);

assign C1119=c10119+c11119+c12119+c13119+c14119+c15119+c16119+c17119+c18119+c19119+c1A119+c1B119+c1C119+c1D119+c1E119+c1F119;
assign A1119=(C1119>=0)?1:0;

assign P2119=A1119;

ninexnine_unit ninexnine_unit_2576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10129)
);

ninexnine_unit ninexnine_unit_2577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11129)
);

ninexnine_unit ninexnine_unit_2578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12129)
);

ninexnine_unit ninexnine_unit_2579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13129)
);

ninexnine_unit ninexnine_unit_2580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14129)
);

ninexnine_unit ninexnine_unit_2581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15129)
);

ninexnine_unit ninexnine_unit_2582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16129)
);

ninexnine_unit ninexnine_unit_2583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17129)
);

ninexnine_unit ninexnine_unit_2584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18129)
);

ninexnine_unit ninexnine_unit_2585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19129)
);

ninexnine_unit ninexnine_unit_2586(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A129)
);

ninexnine_unit ninexnine_unit_2587(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B129)
);

ninexnine_unit ninexnine_unit_2588(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C129)
);

ninexnine_unit ninexnine_unit_2589(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D129)
);

ninexnine_unit ninexnine_unit_2590(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E129)
);

ninexnine_unit ninexnine_unit_2591(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F129)
);

assign C1129=c10129+c11129+c12129+c13129+c14129+c15129+c16129+c17129+c18129+c19129+c1A129+c1B129+c1C129+c1D129+c1E129+c1F129;
assign A1129=(C1129>=0)?1:0;

assign P2129=A1129;

ninexnine_unit ninexnine_unit_2592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10209)
);

ninexnine_unit ninexnine_unit_2593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11209)
);

ninexnine_unit ninexnine_unit_2594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12209)
);

ninexnine_unit ninexnine_unit_2595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13209)
);

ninexnine_unit ninexnine_unit_2596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14209)
);

ninexnine_unit ninexnine_unit_2597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15209)
);

ninexnine_unit ninexnine_unit_2598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16209)
);

ninexnine_unit ninexnine_unit_2599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17209)
);

ninexnine_unit ninexnine_unit_2600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18209)
);

ninexnine_unit ninexnine_unit_2601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19209)
);

ninexnine_unit ninexnine_unit_2602(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A209)
);

ninexnine_unit ninexnine_unit_2603(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B209)
);

ninexnine_unit ninexnine_unit_2604(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C209)
);

ninexnine_unit ninexnine_unit_2605(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D209)
);

ninexnine_unit ninexnine_unit_2606(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E209)
);

ninexnine_unit ninexnine_unit_2607(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F209)
);

assign C1209=c10209+c11209+c12209+c13209+c14209+c15209+c16209+c17209+c18209+c19209+c1A209+c1B209+c1C209+c1D209+c1E209+c1F209;
assign A1209=(C1209>=0)?1:0;

assign P2209=A1209;

ninexnine_unit ninexnine_unit_2608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10219)
);

ninexnine_unit ninexnine_unit_2609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11219)
);

ninexnine_unit ninexnine_unit_2610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12219)
);

ninexnine_unit ninexnine_unit_2611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13219)
);

ninexnine_unit ninexnine_unit_2612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14219)
);

ninexnine_unit ninexnine_unit_2613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15219)
);

ninexnine_unit ninexnine_unit_2614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16219)
);

ninexnine_unit ninexnine_unit_2615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17219)
);

ninexnine_unit ninexnine_unit_2616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18219)
);

ninexnine_unit ninexnine_unit_2617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19219)
);

ninexnine_unit ninexnine_unit_2618(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A219)
);

ninexnine_unit ninexnine_unit_2619(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B219)
);

ninexnine_unit ninexnine_unit_2620(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C219)
);

ninexnine_unit ninexnine_unit_2621(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D219)
);

ninexnine_unit ninexnine_unit_2622(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E219)
);

ninexnine_unit ninexnine_unit_2623(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F219)
);

assign C1219=c10219+c11219+c12219+c13219+c14219+c15219+c16219+c17219+c18219+c19219+c1A219+c1B219+c1C219+c1D219+c1E219+c1F219;
assign A1219=(C1219>=0)?1:0;

assign P2219=A1219;

ninexnine_unit ninexnine_unit_2624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10229)
);

ninexnine_unit ninexnine_unit_2625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11229)
);

ninexnine_unit ninexnine_unit_2626(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12229)
);

ninexnine_unit ninexnine_unit_2627(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W19003),
				.b1(W19013),
				.b2(W19023),
				.b3(W19103),
				.b4(W19113),
				.b5(W19123),
				.b6(W19203),
				.b7(W19213),
				.b8(W19223),
				.c(c13229)
);

ninexnine_unit ninexnine_unit_2628(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W19004),
				.b1(W19014),
				.b2(W19024),
				.b3(W19104),
				.b4(W19114),
				.b5(W19124),
				.b6(W19204),
				.b7(W19214),
				.b8(W19224),
				.c(c14229)
);

ninexnine_unit ninexnine_unit_2629(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W19005),
				.b1(W19015),
				.b2(W19025),
				.b3(W19105),
				.b4(W19115),
				.b5(W19125),
				.b6(W19205),
				.b7(W19215),
				.b8(W19225),
				.c(c15229)
);

ninexnine_unit ninexnine_unit_2630(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W19006),
				.b1(W19016),
				.b2(W19026),
				.b3(W19106),
				.b4(W19116),
				.b5(W19126),
				.b6(W19206),
				.b7(W19216),
				.b8(W19226),
				.c(c16229)
);

ninexnine_unit ninexnine_unit_2631(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W19007),
				.b1(W19017),
				.b2(W19027),
				.b3(W19107),
				.b4(W19117),
				.b5(W19127),
				.b6(W19207),
				.b7(W19217),
				.b8(W19227),
				.c(c17229)
);

ninexnine_unit ninexnine_unit_2632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W19008),
				.b1(W19018),
				.b2(W19028),
				.b3(W19108),
				.b4(W19118),
				.b5(W19128),
				.b6(W19208),
				.b7(W19218),
				.b8(W19228),
				.c(c18229)
);

ninexnine_unit ninexnine_unit_2633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W19009),
				.b1(W19019),
				.b2(W19029),
				.b3(W19109),
				.b4(W19119),
				.b5(W19129),
				.b6(W19209),
				.b7(W19219),
				.b8(W19229),
				.c(c19229)
);

ninexnine_unit ninexnine_unit_2634(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1900A),
				.b1(W1901A),
				.b2(W1902A),
				.b3(W1910A),
				.b4(W1911A),
				.b5(W1912A),
				.b6(W1920A),
				.b7(W1921A),
				.b8(W1922A),
				.c(c1A229)
);

ninexnine_unit ninexnine_unit_2635(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1900B),
				.b1(W1901B),
				.b2(W1902B),
				.b3(W1910B),
				.b4(W1911B),
				.b5(W1912B),
				.b6(W1920B),
				.b7(W1921B),
				.b8(W1922B),
				.c(c1B229)
);

ninexnine_unit ninexnine_unit_2636(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1900C),
				.b1(W1901C),
				.b2(W1902C),
				.b3(W1910C),
				.b4(W1911C),
				.b5(W1912C),
				.b6(W1920C),
				.b7(W1921C),
				.b8(W1922C),
				.c(c1C229)
);

ninexnine_unit ninexnine_unit_2637(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1900D),
				.b1(W1901D),
				.b2(W1902D),
				.b3(W1910D),
				.b4(W1911D),
				.b5(W1912D),
				.b6(W1920D),
				.b7(W1921D),
				.b8(W1922D),
				.c(c1D229)
);

ninexnine_unit ninexnine_unit_2638(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1900E),
				.b1(W1901E),
				.b2(W1902E),
				.b3(W1910E),
				.b4(W1911E),
				.b5(W1912E),
				.b6(W1920E),
				.b7(W1921E),
				.b8(W1922E),
				.c(c1E229)
);

ninexnine_unit ninexnine_unit_2639(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1900F),
				.b1(W1901F),
				.b2(W1902F),
				.b3(W1910F),
				.b4(W1911F),
				.b5(W1912F),
				.b6(W1920F),
				.b7(W1921F),
				.b8(W1922F),
				.c(c1F229)
);

assign C1229=c10229+c11229+c12229+c13229+c14229+c15229+c16229+c17229+c18229+c19229+c1A229+c1B229+c1C229+c1D229+c1E229+c1F229;
assign A1229=(C1229>=0)?1:0;

assign P2229=A1229;

ninexnine_unit ninexnine_unit_2640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1000A)
);

ninexnine_unit ninexnine_unit_2641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1100A)
);

ninexnine_unit ninexnine_unit_2642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1200A)
);

ninexnine_unit ninexnine_unit_2643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1300A)
);

ninexnine_unit ninexnine_unit_2644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1400A)
);

ninexnine_unit ninexnine_unit_2645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1500A)
);

ninexnine_unit ninexnine_unit_2646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1600A)
);

ninexnine_unit ninexnine_unit_2647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1700A)
);

ninexnine_unit ninexnine_unit_2648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1800A)
);

ninexnine_unit ninexnine_unit_2649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1900A)
);

ninexnine_unit ninexnine_unit_2650(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A00A)
);

ninexnine_unit ninexnine_unit_2651(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B00A)
);

ninexnine_unit ninexnine_unit_2652(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C00A)
);

ninexnine_unit ninexnine_unit_2653(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D00A)
);

ninexnine_unit ninexnine_unit_2654(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E00A)
);

ninexnine_unit ninexnine_unit_2655(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F00A)
);

assign C100A=c1000A+c1100A+c1200A+c1300A+c1400A+c1500A+c1600A+c1700A+c1800A+c1900A+c1A00A+c1B00A+c1C00A+c1D00A+c1E00A+c1F00A;
assign A100A=(C100A>=0)?1:0;

assign P200A=A100A;

ninexnine_unit ninexnine_unit_2656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1001A)
);

ninexnine_unit ninexnine_unit_2657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1101A)
);

ninexnine_unit ninexnine_unit_2658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1201A)
);

ninexnine_unit ninexnine_unit_2659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1301A)
);

ninexnine_unit ninexnine_unit_2660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1401A)
);

ninexnine_unit ninexnine_unit_2661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1501A)
);

ninexnine_unit ninexnine_unit_2662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1601A)
);

ninexnine_unit ninexnine_unit_2663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1701A)
);

ninexnine_unit ninexnine_unit_2664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1801A)
);

ninexnine_unit ninexnine_unit_2665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1901A)
);

ninexnine_unit ninexnine_unit_2666(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A01A)
);

ninexnine_unit ninexnine_unit_2667(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B01A)
);

ninexnine_unit ninexnine_unit_2668(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C01A)
);

ninexnine_unit ninexnine_unit_2669(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D01A)
);

ninexnine_unit ninexnine_unit_2670(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E01A)
);

ninexnine_unit ninexnine_unit_2671(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F01A)
);

assign C101A=c1001A+c1101A+c1201A+c1301A+c1401A+c1501A+c1601A+c1701A+c1801A+c1901A+c1A01A+c1B01A+c1C01A+c1D01A+c1E01A+c1F01A;
assign A101A=(C101A>=0)?1:0;

assign P201A=A101A;

ninexnine_unit ninexnine_unit_2672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1002A)
);

ninexnine_unit ninexnine_unit_2673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1102A)
);

ninexnine_unit ninexnine_unit_2674(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1202A)
);

ninexnine_unit ninexnine_unit_2675(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1302A)
);

ninexnine_unit ninexnine_unit_2676(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1402A)
);

ninexnine_unit ninexnine_unit_2677(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1502A)
);

ninexnine_unit ninexnine_unit_2678(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1602A)
);

ninexnine_unit ninexnine_unit_2679(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1702A)
);

ninexnine_unit ninexnine_unit_2680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1802A)
);

ninexnine_unit ninexnine_unit_2681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1902A)
);

ninexnine_unit ninexnine_unit_2682(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A02A)
);

ninexnine_unit ninexnine_unit_2683(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B02A)
);

ninexnine_unit ninexnine_unit_2684(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C02A)
);

ninexnine_unit ninexnine_unit_2685(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D02A)
);

ninexnine_unit ninexnine_unit_2686(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E02A)
);

ninexnine_unit ninexnine_unit_2687(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F02A)
);

assign C102A=c1002A+c1102A+c1202A+c1302A+c1402A+c1502A+c1602A+c1702A+c1802A+c1902A+c1A02A+c1B02A+c1C02A+c1D02A+c1E02A+c1F02A;
assign A102A=(C102A>=0)?1:0;

assign P202A=A102A;

ninexnine_unit ninexnine_unit_2688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1010A)
);

ninexnine_unit ninexnine_unit_2689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1110A)
);

ninexnine_unit ninexnine_unit_2690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1210A)
);

ninexnine_unit ninexnine_unit_2691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1310A)
);

ninexnine_unit ninexnine_unit_2692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1410A)
);

ninexnine_unit ninexnine_unit_2693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1510A)
);

ninexnine_unit ninexnine_unit_2694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1610A)
);

ninexnine_unit ninexnine_unit_2695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1710A)
);

ninexnine_unit ninexnine_unit_2696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1810A)
);

ninexnine_unit ninexnine_unit_2697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1910A)
);

ninexnine_unit ninexnine_unit_2698(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A10A)
);

ninexnine_unit ninexnine_unit_2699(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B10A)
);

ninexnine_unit ninexnine_unit_2700(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C10A)
);

ninexnine_unit ninexnine_unit_2701(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D10A)
);

ninexnine_unit ninexnine_unit_2702(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E10A)
);

ninexnine_unit ninexnine_unit_2703(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F10A)
);

assign C110A=c1010A+c1110A+c1210A+c1310A+c1410A+c1510A+c1610A+c1710A+c1810A+c1910A+c1A10A+c1B10A+c1C10A+c1D10A+c1E10A+c1F10A;
assign A110A=(C110A>=0)?1:0;

assign P210A=A110A;

ninexnine_unit ninexnine_unit_2704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1011A)
);

ninexnine_unit ninexnine_unit_2705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1111A)
);

ninexnine_unit ninexnine_unit_2706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1211A)
);

ninexnine_unit ninexnine_unit_2707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1311A)
);

ninexnine_unit ninexnine_unit_2708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1411A)
);

ninexnine_unit ninexnine_unit_2709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1511A)
);

ninexnine_unit ninexnine_unit_2710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1611A)
);

ninexnine_unit ninexnine_unit_2711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1711A)
);

ninexnine_unit ninexnine_unit_2712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1811A)
);

ninexnine_unit ninexnine_unit_2713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1911A)
);

ninexnine_unit ninexnine_unit_2714(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A11A)
);

ninexnine_unit ninexnine_unit_2715(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B11A)
);

ninexnine_unit ninexnine_unit_2716(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C11A)
);

ninexnine_unit ninexnine_unit_2717(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D11A)
);

ninexnine_unit ninexnine_unit_2718(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E11A)
);

ninexnine_unit ninexnine_unit_2719(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F11A)
);

assign C111A=c1011A+c1111A+c1211A+c1311A+c1411A+c1511A+c1611A+c1711A+c1811A+c1911A+c1A11A+c1B11A+c1C11A+c1D11A+c1E11A+c1F11A;
assign A111A=(C111A>=0)?1:0;

assign P211A=A111A;

ninexnine_unit ninexnine_unit_2720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1012A)
);

ninexnine_unit ninexnine_unit_2721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1112A)
);

ninexnine_unit ninexnine_unit_2722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1212A)
);

ninexnine_unit ninexnine_unit_2723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1312A)
);

ninexnine_unit ninexnine_unit_2724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1412A)
);

ninexnine_unit ninexnine_unit_2725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1512A)
);

ninexnine_unit ninexnine_unit_2726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1612A)
);

ninexnine_unit ninexnine_unit_2727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1712A)
);

ninexnine_unit ninexnine_unit_2728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1812A)
);

ninexnine_unit ninexnine_unit_2729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1912A)
);

ninexnine_unit ninexnine_unit_2730(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A12A)
);

ninexnine_unit ninexnine_unit_2731(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B12A)
);

ninexnine_unit ninexnine_unit_2732(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C12A)
);

ninexnine_unit ninexnine_unit_2733(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D12A)
);

ninexnine_unit ninexnine_unit_2734(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E12A)
);

ninexnine_unit ninexnine_unit_2735(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F12A)
);

assign C112A=c1012A+c1112A+c1212A+c1312A+c1412A+c1512A+c1612A+c1712A+c1812A+c1912A+c1A12A+c1B12A+c1C12A+c1D12A+c1E12A+c1F12A;
assign A112A=(C112A>=0)?1:0;

assign P212A=A112A;

ninexnine_unit ninexnine_unit_2736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1020A)
);

ninexnine_unit ninexnine_unit_2737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1120A)
);

ninexnine_unit ninexnine_unit_2738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1220A)
);

ninexnine_unit ninexnine_unit_2739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1320A)
);

ninexnine_unit ninexnine_unit_2740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1420A)
);

ninexnine_unit ninexnine_unit_2741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1520A)
);

ninexnine_unit ninexnine_unit_2742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1620A)
);

ninexnine_unit ninexnine_unit_2743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1720A)
);

ninexnine_unit ninexnine_unit_2744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1820A)
);

ninexnine_unit ninexnine_unit_2745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1920A)
);

ninexnine_unit ninexnine_unit_2746(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A20A)
);

ninexnine_unit ninexnine_unit_2747(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B20A)
);

ninexnine_unit ninexnine_unit_2748(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C20A)
);

ninexnine_unit ninexnine_unit_2749(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D20A)
);

ninexnine_unit ninexnine_unit_2750(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E20A)
);

ninexnine_unit ninexnine_unit_2751(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F20A)
);

assign C120A=c1020A+c1120A+c1220A+c1320A+c1420A+c1520A+c1620A+c1720A+c1820A+c1920A+c1A20A+c1B20A+c1C20A+c1D20A+c1E20A+c1F20A;
assign A120A=(C120A>=0)?1:0;

assign P220A=A120A;

ninexnine_unit ninexnine_unit_2752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1021A)
);

ninexnine_unit ninexnine_unit_2753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1121A)
);

ninexnine_unit ninexnine_unit_2754(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1221A)
);

ninexnine_unit ninexnine_unit_2755(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1321A)
);

ninexnine_unit ninexnine_unit_2756(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1421A)
);

ninexnine_unit ninexnine_unit_2757(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1521A)
);

ninexnine_unit ninexnine_unit_2758(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1621A)
);

ninexnine_unit ninexnine_unit_2759(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1721A)
);

ninexnine_unit ninexnine_unit_2760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1821A)
);

ninexnine_unit ninexnine_unit_2761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1921A)
);

ninexnine_unit ninexnine_unit_2762(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A21A)
);

ninexnine_unit ninexnine_unit_2763(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B21A)
);

ninexnine_unit ninexnine_unit_2764(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C21A)
);

ninexnine_unit ninexnine_unit_2765(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D21A)
);

ninexnine_unit ninexnine_unit_2766(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E21A)
);

ninexnine_unit ninexnine_unit_2767(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F21A)
);

assign C121A=c1021A+c1121A+c1221A+c1321A+c1421A+c1521A+c1621A+c1721A+c1821A+c1921A+c1A21A+c1B21A+c1C21A+c1D21A+c1E21A+c1F21A;
assign A121A=(C121A>=0)?1:0;

assign P221A=A121A;

ninexnine_unit ninexnine_unit_2768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1022A)
);

ninexnine_unit ninexnine_unit_2769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1122A)
);

ninexnine_unit ninexnine_unit_2770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1222A)
);

ninexnine_unit ninexnine_unit_2771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1A003),
				.b1(W1A013),
				.b2(W1A023),
				.b3(W1A103),
				.b4(W1A113),
				.b5(W1A123),
				.b6(W1A203),
				.b7(W1A213),
				.b8(W1A223),
				.c(c1322A)
);

ninexnine_unit ninexnine_unit_2772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1A004),
				.b1(W1A014),
				.b2(W1A024),
				.b3(W1A104),
				.b4(W1A114),
				.b5(W1A124),
				.b6(W1A204),
				.b7(W1A214),
				.b8(W1A224),
				.c(c1422A)
);

ninexnine_unit ninexnine_unit_2773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1A005),
				.b1(W1A015),
				.b2(W1A025),
				.b3(W1A105),
				.b4(W1A115),
				.b5(W1A125),
				.b6(W1A205),
				.b7(W1A215),
				.b8(W1A225),
				.c(c1522A)
);

ninexnine_unit ninexnine_unit_2774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1A006),
				.b1(W1A016),
				.b2(W1A026),
				.b3(W1A106),
				.b4(W1A116),
				.b5(W1A126),
				.b6(W1A206),
				.b7(W1A216),
				.b8(W1A226),
				.c(c1622A)
);

ninexnine_unit ninexnine_unit_2775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1A007),
				.b1(W1A017),
				.b2(W1A027),
				.b3(W1A107),
				.b4(W1A117),
				.b5(W1A127),
				.b6(W1A207),
				.b7(W1A217),
				.b8(W1A227),
				.c(c1722A)
);

ninexnine_unit ninexnine_unit_2776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1A008),
				.b1(W1A018),
				.b2(W1A028),
				.b3(W1A108),
				.b4(W1A118),
				.b5(W1A128),
				.b6(W1A208),
				.b7(W1A218),
				.b8(W1A228),
				.c(c1822A)
);

ninexnine_unit ninexnine_unit_2777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1A009),
				.b1(W1A019),
				.b2(W1A029),
				.b3(W1A109),
				.b4(W1A119),
				.b5(W1A129),
				.b6(W1A209),
				.b7(W1A219),
				.b8(W1A229),
				.c(c1922A)
);

ninexnine_unit ninexnine_unit_2778(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1A00A),
				.b1(W1A01A),
				.b2(W1A02A),
				.b3(W1A10A),
				.b4(W1A11A),
				.b5(W1A12A),
				.b6(W1A20A),
				.b7(W1A21A),
				.b8(W1A22A),
				.c(c1A22A)
);

ninexnine_unit ninexnine_unit_2779(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1A00B),
				.b1(W1A01B),
				.b2(W1A02B),
				.b3(W1A10B),
				.b4(W1A11B),
				.b5(W1A12B),
				.b6(W1A20B),
				.b7(W1A21B),
				.b8(W1A22B),
				.c(c1B22A)
);

ninexnine_unit ninexnine_unit_2780(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1A00C),
				.b1(W1A01C),
				.b2(W1A02C),
				.b3(W1A10C),
				.b4(W1A11C),
				.b5(W1A12C),
				.b6(W1A20C),
				.b7(W1A21C),
				.b8(W1A22C),
				.c(c1C22A)
);

ninexnine_unit ninexnine_unit_2781(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1A00D),
				.b1(W1A01D),
				.b2(W1A02D),
				.b3(W1A10D),
				.b4(W1A11D),
				.b5(W1A12D),
				.b6(W1A20D),
				.b7(W1A21D),
				.b8(W1A22D),
				.c(c1D22A)
);

ninexnine_unit ninexnine_unit_2782(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1A00E),
				.b1(W1A01E),
				.b2(W1A02E),
				.b3(W1A10E),
				.b4(W1A11E),
				.b5(W1A12E),
				.b6(W1A20E),
				.b7(W1A21E),
				.b8(W1A22E),
				.c(c1E22A)
);

ninexnine_unit ninexnine_unit_2783(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1A00F),
				.b1(W1A01F),
				.b2(W1A02F),
				.b3(W1A10F),
				.b4(W1A11F),
				.b5(W1A12F),
				.b6(W1A20F),
				.b7(W1A21F),
				.b8(W1A22F),
				.c(c1F22A)
);

assign C122A=c1022A+c1122A+c1222A+c1322A+c1422A+c1522A+c1622A+c1722A+c1822A+c1922A+c1A22A+c1B22A+c1C22A+c1D22A+c1E22A+c1F22A;
assign A122A=(C122A>=0)?1:0;

assign P222A=A122A;

ninexnine_unit ninexnine_unit_2784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1000B)
);

ninexnine_unit ninexnine_unit_2785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1100B)
);

ninexnine_unit ninexnine_unit_2786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1200B)
);

ninexnine_unit ninexnine_unit_2787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1300B)
);

ninexnine_unit ninexnine_unit_2788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1400B)
);

ninexnine_unit ninexnine_unit_2789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1500B)
);

ninexnine_unit ninexnine_unit_2790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1600B)
);

ninexnine_unit ninexnine_unit_2791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1700B)
);

ninexnine_unit ninexnine_unit_2792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1800B)
);

ninexnine_unit ninexnine_unit_2793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1900B)
);

ninexnine_unit ninexnine_unit_2794(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A00B)
);

ninexnine_unit ninexnine_unit_2795(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B00B)
);

ninexnine_unit ninexnine_unit_2796(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C00B)
);

ninexnine_unit ninexnine_unit_2797(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D00B)
);

ninexnine_unit ninexnine_unit_2798(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E00B)
);

ninexnine_unit ninexnine_unit_2799(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F00B)
);

assign C100B=c1000B+c1100B+c1200B+c1300B+c1400B+c1500B+c1600B+c1700B+c1800B+c1900B+c1A00B+c1B00B+c1C00B+c1D00B+c1E00B+c1F00B;
assign A100B=(C100B>=0)?1:0;

assign P200B=A100B;

ninexnine_unit ninexnine_unit_2800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1001B)
);

ninexnine_unit ninexnine_unit_2801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1101B)
);

ninexnine_unit ninexnine_unit_2802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1201B)
);

ninexnine_unit ninexnine_unit_2803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1301B)
);

ninexnine_unit ninexnine_unit_2804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1401B)
);

ninexnine_unit ninexnine_unit_2805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1501B)
);

ninexnine_unit ninexnine_unit_2806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1601B)
);

ninexnine_unit ninexnine_unit_2807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1701B)
);

ninexnine_unit ninexnine_unit_2808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1801B)
);

ninexnine_unit ninexnine_unit_2809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1901B)
);

ninexnine_unit ninexnine_unit_2810(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A01B)
);

ninexnine_unit ninexnine_unit_2811(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B01B)
);

ninexnine_unit ninexnine_unit_2812(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C01B)
);

ninexnine_unit ninexnine_unit_2813(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D01B)
);

ninexnine_unit ninexnine_unit_2814(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E01B)
);

ninexnine_unit ninexnine_unit_2815(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F01B)
);

assign C101B=c1001B+c1101B+c1201B+c1301B+c1401B+c1501B+c1601B+c1701B+c1801B+c1901B+c1A01B+c1B01B+c1C01B+c1D01B+c1E01B+c1F01B;
assign A101B=(C101B>=0)?1:0;

assign P201B=A101B;

ninexnine_unit ninexnine_unit_2816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1002B)
);

ninexnine_unit ninexnine_unit_2817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1102B)
);

ninexnine_unit ninexnine_unit_2818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1202B)
);

ninexnine_unit ninexnine_unit_2819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1302B)
);

ninexnine_unit ninexnine_unit_2820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1402B)
);

ninexnine_unit ninexnine_unit_2821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1502B)
);

ninexnine_unit ninexnine_unit_2822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1602B)
);

ninexnine_unit ninexnine_unit_2823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1702B)
);

ninexnine_unit ninexnine_unit_2824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1802B)
);

ninexnine_unit ninexnine_unit_2825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1902B)
);

ninexnine_unit ninexnine_unit_2826(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A02B)
);

ninexnine_unit ninexnine_unit_2827(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B02B)
);

ninexnine_unit ninexnine_unit_2828(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C02B)
);

ninexnine_unit ninexnine_unit_2829(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D02B)
);

ninexnine_unit ninexnine_unit_2830(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E02B)
);

ninexnine_unit ninexnine_unit_2831(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F02B)
);

assign C102B=c1002B+c1102B+c1202B+c1302B+c1402B+c1502B+c1602B+c1702B+c1802B+c1902B+c1A02B+c1B02B+c1C02B+c1D02B+c1E02B+c1F02B;
assign A102B=(C102B>=0)?1:0;

assign P202B=A102B;

ninexnine_unit ninexnine_unit_2832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1010B)
);

ninexnine_unit ninexnine_unit_2833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1110B)
);

ninexnine_unit ninexnine_unit_2834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1210B)
);

ninexnine_unit ninexnine_unit_2835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1310B)
);

ninexnine_unit ninexnine_unit_2836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1410B)
);

ninexnine_unit ninexnine_unit_2837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1510B)
);

ninexnine_unit ninexnine_unit_2838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1610B)
);

ninexnine_unit ninexnine_unit_2839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1710B)
);

ninexnine_unit ninexnine_unit_2840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1810B)
);

ninexnine_unit ninexnine_unit_2841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1910B)
);

ninexnine_unit ninexnine_unit_2842(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A10B)
);

ninexnine_unit ninexnine_unit_2843(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B10B)
);

ninexnine_unit ninexnine_unit_2844(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C10B)
);

ninexnine_unit ninexnine_unit_2845(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D10B)
);

ninexnine_unit ninexnine_unit_2846(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E10B)
);

ninexnine_unit ninexnine_unit_2847(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F10B)
);

assign C110B=c1010B+c1110B+c1210B+c1310B+c1410B+c1510B+c1610B+c1710B+c1810B+c1910B+c1A10B+c1B10B+c1C10B+c1D10B+c1E10B+c1F10B;
assign A110B=(C110B>=0)?1:0;

assign P210B=A110B;

ninexnine_unit ninexnine_unit_2848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1011B)
);

ninexnine_unit ninexnine_unit_2849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1111B)
);

ninexnine_unit ninexnine_unit_2850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1211B)
);

ninexnine_unit ninexnine_unit_2851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1311B)
);

ninexnine_unit ninexnine_unit_2852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1411B)
);

ninexnine_unit ninexnine_unit_2853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1511B)
);

ninexnine_unit ninexnine_unit_2854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1611B)
);

ninexnine_unit ninexnine_unit_2855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1711B)
);

ninexnine_unit ninexnine_unit_2856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1811B)
);

ninexnine_unit ninexnine_unit_2857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1911B)
);

ninexnine_unit ninexnine_unit_2858(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A11B)
);

ninexnine_unit ninexnine_unit_2859(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B11B)
);

ninexnine_unit ninexnine_unit_2860(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C11B)
);

ninexnine_unit ninexnine_unit_2861(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D11B)
);

ninexnine_unit ninexnine_unit_2862(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E11B)
);

ninexnine_unit ninexnine_unit_2863(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F11B)
);

assign C111B=c1011B+c1111B+c1211B+c1311B+c1411B+c1511B+c1611B+c1711B+c1811B+c1911B+c1A11B+c1B11B+c1C11B+c1D11B+c1E11B+c1F11B;
assign A111B=(C111B>=0)?1:0;

assign P211B=A111B;

ninexnine_unit ninexnine_unit_2864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1012B)
);

ninexnine_unit ninexnine_unit_2865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1112B)
);

ninexnine_unit ninexnine_unit_2866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1212B)
);

ninexnine_unit ninexnine_unit_2867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1312B)
);

ninexnine_unit ninexnine_unit_2868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1412B)
);

ninexnine_unit ninexnine_unit_2869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1512B)
);

ninexnine_unit ninexnine_unit_2870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1612B)
);

ninexnine_unit ninexnine_unit_2871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1712B)
);

ninexnine_unit ninexnine_unit_2872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1812B)
);

ninexnine_unit ninexnine_unit_2873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1912B)
);

ninexnine_unit ninexnine_unit_2874(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A12B)
);

ninexnine_unit ninexnine_unit_2875(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B12B)
);

ninexnine_unit ninexnine_unit_2876(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C12B)
);

ninexnine_unit ninexnine_unit_2877(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D12B)
);

ninexnine_unit ninexnine_unit_2878(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E12B)
);

ninexnine_unit ninexnine_unit_2879(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F12B)
);

assign C112B=c1012B+c1112B+c1212B+c1312B+c1412B+c1512B+c1612B+c1712B+c1812B+c1912B+c1A12B+c1B12B+c1C12B+c1D12B+c1E12B+c1F12B;
assign A112B=(C112B>=0)?1:0;

assign P212B=A112B;

ninexnine_unit ninexnine_unit_2880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1020B)
);

ninexnine_unit ninexnine_unit_2881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1120B)
);

ninexnine_unit ninexnine_unit_2882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1220B)
);

ninexnine_unit ninexnine_unit_2883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1320B)
);

ninexnine_unit ninexnine_unit_2884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1420B)
);

ninexnine_unit ninexnine_unit_2885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1520B)
);

ninexnine_unit ninexnine_unit_2886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1620B)
);

ninexnine_unit ninexnine_unit_2887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1720B)
);

ninexnine_unit ninexnine_unit_2888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1820B)
);

ninexnine_unit ninexnine_unit_2889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1920B)
);

ninexnine_unit ninexnine_unit_2890(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A20B)
);

ninexnine_unit ninexnine_unit_2891(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B20B)
);

ninexnine_unit ninexnine_unit_2892(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C20B)
);

ninexnine_unit ninexnine_unit_2893(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D20B)
);

ninexnine_unit ninexnine_unit_2894(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E20B)
);

ninexnine_unit ninexnine_unit_2895(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F20B)
);

assign C120B=c1020B+c1120B+c1220B+c1320B+c1420B+c1520B+c1620B+c1720B+c1820B+c1920B+c1A20B+c1B20B+c1C20B+c1D20B+c1E20B+c1F20B;
assign A120B=(C120B>=0)?1:0;

assign P220B=A120B;

ninexnine_unit ninexnine_unit_2896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1021B)
);

ninexnine_unit ninexnine_unit_2897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1121B)
);

ninexnine_unit ninexnine_unit_2898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1221B)
);

ninexnine_unit ninexnine_unit_2899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1321B)
);

ninexnine_unit ninexnine_unit_2900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1421B)
);

ninexnine_unit ninexnine_unit_2901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1521B)
);

ninexnine_unit ninexnine_unit_2902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1621B)
);

ninexnine_unit ninexnine_unit_2903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1721B)
);

ninexnine_unit ninexnine_unit_2904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1821B)
);

ninexnine_unit ninexnine_unit_2905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1921B)
);

ninexnine_unit ninexnine_unit_2906(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A21B)
);

ninexnine_unit ninexnine_unit_2907(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B21B)
);

ninexnine_unit ninexnine_unit_2908(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C21B)
);

ninexnine_unit ninexnine_unit_2909(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D21B)
);

ninexnine_unit ninexnine_unit_2910(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E21B)
);

ninexnine_unit ninexnine_unit_2911(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F21B)
);

assign C121B=c1021B+c1121B+c1221B+c1321B+c1421B+c1521B+c1621B+c1721B+c1821B+c1921B+c1A21B+c1B21B+c1C21B+c1D21B+c1E21B+c1F21B;
assign A121B=(C121B>=0)?1:0;

assign P221B=A121B;

ninexnine_unit ninexnine_unit_2912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1022B)
);

ninexnine_unit ninexnine_unit_2913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1122B)
);

ninexnine_unit ninexnine_unit_2914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1222B)
);

ninexnine_unit ninexnine_unit_2915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1B003),
				.b1(W1B013),
				.b2(W1B023),
				.b3(W1B103),
				.b4(W1B113),
				.b5(W1B123),
				.b6(W1B203),
				.b7(W1B213),
				.b8(W1B223),
				.c(c1322B)
);

ninexnine_unit ninexnine_unit_2916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1B004),
				.b1(W1B014),
				.b2(W1B024),
				.b3(W1B104),
				.b4(W1B114),
				.b5(W1B124),
				.b6(W1B204),
				.b7(W1B214),
				.b8(W1B224),
				.c(c1422B)
);

ninexnine_unit ninexnine_unit_2917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1B005),
				.b1(W1B015),
				.b2(W1B025),
				.b3(W1B105),
				.b4(W1B115),
				.b5(W1B125),
				.b6(W1B205),
				.b7(W1B215),
				.b8(W1B225),
				.c(c1522B)
);

ninexnine_unit ninexnine_unit_2918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1B006),
				.b1(W1B016),
				.b2(W1B026),
				.b3(W1B106),
				.b4(W1B116),
				.b5(W1B126),
				.b6(W1B206),
				.b7(W1B216),
				.b8(W1B226),
				.c(c1622B)
);

ninexnine_unit ninexnine_unit_2919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1B007),
				.b1(W1B017),
				.b2(W1B027),
				.b3(W1B107),
				.b4(W1B117),
				.b5(W1B127),
				.b6(W1B207),
				.b7(W1B217),
				.b8(W1B227),
				.c(c1722B)
);

ninexnine_unit ninexnine_unit_2920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1B008),
				.b1(W1B018),
				.b2(W1B028),
				.b3(W1B108),
				.b4(W1B118),
				.b5(W1B128),
				.b6(W1B208),
				.b7(W1B218),
				.b8(W1B228),
				.c(c1822B)
);

ninexnine_unit ninexnine_unit_2921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1B009),
				.b1(W1B019),
				.b2(W1B029),
				.b3(W1B109),
				.b4(W1B119),
				.b5(W1B129),
				.b6(W1B209),
				.b7(W1B219),
				.b8(W1B229),
				.c(c1922B)
);

ninexnine_unit ninexnine_unit_2922(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1B00A),
				.b1(W1B01A),
				.b2(W1B02A),
				.b3(W1B10A),
				.b4(W1B11A),
				.b5(W1B12A),
				.b6(W1B20A),
				.b7(W1B21A),
				.b8(W1B22A),
				.c(c1A22B)
);

ninexnine_unit ninexnine_unit_2923(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1B00B),
				.b1(W1B01B),
				.b2(W1B02B),
				.b3(W1B10B),
				.b4(W1B11B),
				.b5(W1B12B),
				.b6(W1B20B),
				.b7(W1B21B),
				.b8(W1B22B),
				.c(c1B22B)
);

ninexnine_unit ninexnine_unit_2924(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1B00C),
				.b1(W1B01C),
				.b2(W1B02C),
				.b3(W1B10C),
				.b4(W1B11C),
				.b5(W1B12C),
				.b6(W1B20C),
				.b7(W1B21C),
				.b8(W1B22C),
				.c(c1C22B)
);

ninexnine_unit ninexnine_unit_2925(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1B00D),
				.b1(W1B01D),
				.b2(W1B02D),
				.b3(W1B10D),
				.b4(W1B11D),
				.b5(W1B12D),
				.b6(W1B20D),
				.b7(W1B21D),
				.b8(W1B22D),
				.c(c1D22B)
);

ninexnine_unit ninexnine_unit_2926(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1B00E),
				.b1(W1B01E),
				.b2(W1B02E),
				.b3(W1B10E),
				.b4(W1B11E),
				.b5(W1B12E),
				.b6(W1B20E),
				.b7(W1B21E),
				.b8(W1B22E),
				.c(c1E22B)
);

ninexnine_unit ninexnine_unit_2927(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1B00F),
				.b1(W1B01F),
				.b2(W1B02F),
				.b3(W1B10F),
				.b4(W1B11F),
				.b5(W1B12F),
				.b6(W1B20F),
				.b7(W1B21F),
				.b8(W1B22F),
				.c(c1F22B)
);

assign C122B=c1022B+c1122B+c1222B+c1322B+c1422B+c1522B+c1622B+c1722B+c1822B+c1922B+c1A22B+c1B22B+c1C22B+c1D22B+c1E22B+c1F22B;
assign A122B=(C122B>=0)?1:0;

assign P222B=A122B;

ninexnine_unit ninexnine_unit_2928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1000C)
);

ninexnine_unit ninexnine_unit_2929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1100C)
);

ninexnine_unit ninexnine_unit_2930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1200C)
);

ninexnine_unit ninexnine_unit_2931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1300C)
);

ninexnine_unit ninexnine_unit_2932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1400C)
);

ninexnine_unit ninexnine_unit_2933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1500C)
);

ninexnine_unit ninexnine_unit_2934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1600C)
);

ninexnine_unit ninexnine_unit_2935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1700C)
);

ninexnine_unit ninexnine_unit_2936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1800C)
);

ninexnine_unit ninexnine_unit_2937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1900C)
);

ninexnine_unit ninexnine_unit_2938(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A00C)
);

ninexnine_unit ninexnine_unit_2939(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B00C)
);

ninexnine_unit ninexnine_unit_2940(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C00C)
);

ninexnine_unit ninexnine_unit_2941(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D00C)
);

ninexnine_unit ninexnine_unit_2942(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E00C)
);

ninexnine_unit ninexnine_unit_2943(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F00C)
);

assign C100C=c1000C+c1100C+c1200C+c1300C+c1400C+c1500C+c1600C+c1700C+c1800C+c1900C+c1A00C+c1B00C+c1C00C+c1D00C+c1E00C+c1F00C;
assign A100C=(C100C>=0)?1:0;

assign P200C=A100C;

ninexnine_unit ninexnine_unit_2944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1001C)
);

ninexnine_unit ninexnine_unit_2945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1101C)
);

ninexnine_unit ninexnine_unit_2946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1201C)
);

ninexnine_unit ninexnine_unit_2947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1301C)
);

ninexnine_unit ninexnine_unit_2948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1401C)
);

ninexnine_unit ninexnine_unit_2949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1501C)
);

ninexnine_unit ninexnine_unit_2950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1601C)
);

ninexnine_unit ninexnine_unit_2951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1701C)
);

ninexnine_unit ninexnine_unit_2952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1801C)
);

ninexnine_unit ninexnine_unit_2953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1901C)
);

ninexnine_unit ninexnine_unit_2954(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A01C)
);

ninexnine_unit ninexnine_unit_2955(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B01C)
);

ninexnine_unit ninexnine_unit_2956(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C01C)
);

ninexnine_unit ninexnine_unit_2957(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D01C)
);

ninexnine_unit ninexnine_unit_2958(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E01C)
);

ninexnine_unit ninexnine_unit_2959(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F01C)
);

assign C101C=c1001C+c1101C+c1201C+c1301C+c1401C+c1501C+c1601C+c1701C+c1801C+c1901C+c1A01C+c1B01C+c1C01C+c1D01C+c1E01C+c1F01C;
assign A101C=(C101C>=0)?1:0;

assign P201C=A101C;

ninexnine_unit ninexnine_unit_2960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1002C)
);

ninexnine_unit ninexnine_unit_2961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1102C)
);

ninexnine_unit ninexnine_unit_2962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1202C)
);

ninexnine_unit ninexnine_unit_2963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1302C)
);

ninexnine_unit ninexnine_unit_2964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1402C)
);

ninexnine_unit ninexnine_unit_2965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1502C)
);

ninexnine_unit ninexnine_unit_2966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1602C)
);

ninexnine_unit ninexnine_unit_2967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1702C)
);

ninexnine_unit ninexnine_unit_2968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1802C)
);

ninexnine_unit ninexnine_unit_2969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1902C)
);

ninexnine_unit ninexnine_unit_2970(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A02C)
);

ninexnine_unit ninexnine_unit_2971(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B02C)
);

ninexnine_unit ninexnine_unit_2972(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C02C)
);

ninexnine_unit ninexnine_unit_2973(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D02C)
);

ninexnine_unit ninexnine_unit_2974(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E02C)
);

ninexnine_unit ninexnine_unit_2975(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F02C)
);

assign C102C=c1002C+c1102C+c1202C+c1302C+c1402C+c1502C+c1602C+c1702C+c1802C+c1902C+c1A02C+c1B02C+c1C02C+c1D02C+c1E02C+c1F02C;
assign A102C=(C102C>=0)?1:0;

assign P202C=A102C;

ninexnine_unit ninexnine_unit_2976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1010C)
);

ninexnine_unit ninexnine_unit_2977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1110C)
);

ninexnine_unit ninexnine_unit_2978(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1210C)
);

ninexnine_unit ninexnine_unit_2979(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1310C)
);

ninexnine_unit ninexnine_unit_2980(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1410C)
);

ninexnine_unit ninexnine_unit_2981(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1510C)
);

ninexnine_unit ninexnine_unit_2982(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1610C)
);

ninexnine_unit ninexnine_unit_2983(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1710C)
);

ninexnine_unit ninexnine_unit_2984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1810C)
);

ninexnine_unit ninexnine_unit_2985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1910C)
);

ninexnine_unit ninexnine_unit_2986(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A10C)
);

ninexnine_unit ninexnine_unit_2987(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B10C)
);

ninexnine_unit ninexnine_unit_2988(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C10C)
);

ninexnine_unit ninexnine_unit_2989(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D10C)
);

ninexnine_unit ninexnine_unit_2990(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E10C)
);

ninexnine_unit ninexnine_unit_2991(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F10C)
);

assign C110C=c1010C+c1110C+c1210C+c1310C+c1410C+c1510C+c1610C+c1710C+c1810C+c1910C+c1A10C+c1B10C+c1C10C+c1D10C+c1E10C+c1F10C;
assign A110C=(C110C>=0)?1:0;

assign P210C=A110C;

ninexnine_unit ninexnine_unit_2992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1011C)
);

ninexnine_unit ninexnine_unit_2993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1111C)
);

ninexnine_unit ninexnine_unit_2994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1211C)
);

ninexnine_unit ninexnine_unit_2995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1311C)
);

ninexnine_unit ninexnine_unit_2996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1411C)
);

ninexnine_unit ninexnine_unit_2997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1511C)
);

ninexnine_unit ninexnine_unit_2998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1611C)
);

ninexnine_unit ninexnine_unit_2999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1711C)
);

ninexnine_unit ninexnine_unit_3000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1811C)
);

ninexnine_unit ninexnine_unit_3001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1911C)
);

ninexnine_unit ninexnine_unit_3002(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A11C)
);

ninexnine_unit ninexnine_unit_3003(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B11C)
);

ninexnine_unit ninexnine_unit_3004(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C11C)
);

ninexnine_unit ninexnine_unit_3005(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D11C)
);

ninexnine_unit ninexnine_unit_3006(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E11C)
);

ninexnine_unit ninexnine_unit_3007(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F11C)
);

assign C111C=c1011C+c1111C+c1211C+c1311C+c1411C+c1511C+c1611C+c1711C+c1811C+c1911C+c1A11C+c1B11C+c1C11C+c1D11C+c1E11C+c1F11C;
assign A111C=(C111C>=0)?1:0;

assign P211C=A111C;

ninexnine_unit ninexnine_unit_3008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1012C)
);

ninexnine_unit ninexnine_unit_3009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1112C)
);

ninexnine_unit ninexnine_unit_3010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1212C)
);

ninexnine_unit ninexnine_unit_3011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1312C)
);

ninexnine_unit ninexnine_unit_3012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1412C)
);

ninexnine_unit ninexnine_unit_3013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1512C)
);

ninexnine_unit ninexnine_unit_3014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1612C)
);

ninexnine_unit ninexnine_unit_3015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1712C)
);

ninexnine_unit ninexnine_unit_3016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1812C)
);

ninexnine_unit ninexnine_unit_3017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1912C)
);

ninexnine_unit ninexnine_unit_3018(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A12C)
);

ninexnine_unit ninexnine_unit_3019(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B12C)
);

ninexnine_unit ninexnine_unit_3020(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C12C)
);

ninexnine_unit ninexnine_unit_3021(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D12C)
);

ninexnine_unit ninexnine_unit_3022(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E12C)
);

ninexnine_unit ninexnine_unit_3023(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F12C)
);

assign C112C=c1012C+c1112C+c1212C+c1312C+c1412C+c1512C+c1612C+c1712C+c1812C+c1912C+c1A12C+c1B12C+c1C12C+c1D12C+c1E12C+c1F12C;
assign A112C=(C112C>=0)?1:0;

assign P212C=A112C;

ninexnine_unit ninexnine_unit_3024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1020C)
);

ninexnine_unit ninexnine_unit_3025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1120C)
);

ninexnine_unit ninexnine_unit_3026(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1220C)
);

ninexnine_unit ninexnine_unit_3027(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1320C)
);

ninexnine_unit ninexnine_unit_3028(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1420C)
);

ninexnine_unit ninexnine_unit_3029(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1520C)
);

ninexnine_unit ninexnine_unit_3030(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1620C)
);

ninexnine_unit ninexnine_unit_3031(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1720C)
);

ninexnine_unit ninexnine_unit_3032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1820C)
);

ninexnine_unit ninexnine_unit_3033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1920C)
);

ninexnine_unit ninexnine_unit_3034(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A20C)
);

ninexnine_unit ninexnine_unit_3035(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B20C)
);

ninexnine_unit ninexnine_unit_3036(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C20C)
);

ninexnine_unit ninexnine_unit_3037(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D20C)
);

ninexnine_unit ninexnine_unit_3038(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E20C)
);

ninexnine_unit ninexnine_unit_3039(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F20C)
);

assign C120C=c1020C+c1120C+c1220C+c1320C+c1420C+c1520C+c1620C+c1720C+c1820C+c1920C+c1A20C+c1B20C+c1C20C+c1D20C+c1E20C+c1F20C;
assign A120C=(C120C>=0)?1:0;

assign P220C=A120C;

ninexnine_unit ninexnine_unit_3040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1021C)
);

ninexnine_unit ninexnine_unit_3041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1121C)
);

ninexnine_unit ninexnine_unit_3042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1221C)
);

ninexnine_unit ninexnine_unit_3043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1321C)
);

ninexnine_unit ninexnine_unit_3044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1421C)
);

ninexnine_unit ninexnine_unit_3045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1521C)
);

ninexnine_unit ninexnine_unit_3046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1621C)
);

ninexnine_unit ninexnine_unit_3047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1721C)
);

ninexnine_unit ninexnine_unit_3048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1821C)
);

ninexnine_unit ninexnine_unit_3049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1921C)
);

ninexnine_unit ninexnine_unit_3050(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A21C)
);

ninexnine_unit ninexnine_unit_3051(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B21C)
);

ninexnine_unit ninexnine_unit_3052(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C21C)
);

ninexnine_unit ninexnine_unit_3053(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D21C)
);

ninexnine_unit ninexnine_unit_3054(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E21C)
);

ninexnine_unit ninexnine_unit_3055(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F21C)
);

assign C121C=c1021C+c1121C+c1221C+c1321C+c1421C+c1521C+c1621C+c1721C+c1821C+c1921C+c1A21C+c1B21C+c1C21C+c1D21C+c1E21C+c1F21C;
assign A121C=(C121C>=0)?1:0;

assign P221C=A121C;

ninexnine_unit ninexnine_unit_3056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1022C)
);

ninexnine_unit ninexnine_unit_3057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1122C)
);

ninexnine_unit ninexnine_unit_3058(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1222C)
);

ninexnine_unit ninexnine_unit_3059(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1C003),
				.b1(W1C013),
				.b2(W1C023),
				.b3(W1C103),
				.b4(W1C113),
				.b5(W1C123),
				.b6(W1C203),
				.b7(W1C213),
				.b8(W1C223),
				.c(c1322C)
);

ninexnine_unit ninexnine_unit_3060(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1C004),
				.b1(W1C014),
				.b2(W1C024),
				.b3(W1C104),
				.b4(W1C114),
				.b5(W1C124),
				.b6(W1C204),
				.b7(W1C214),
				.b8(W1C224),
				.c(c1422C)
);

ninexnine_unit ninexnine_unit_3061(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1C005),
				.b1(W1C015),
				.b2(W1C025),
				.b3(W1C105),
				.b4(W1C115),
				.b5(W1C125),
				.b6(W1C205),
				.b7(W1C215),
				.b8(W1C225),
				.c(c1522C)
);

ninexnine_unit ninexnine_unit_3062(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1C006),
				.b1(W1C016),
				.b2(W1C026),
				.b3(W1C106),
				.b4(W1C116),
				.b5(W1C126),
				.b6(W1C206),
				.b7(W1C216),
				.b8(W1C226),
				.c(c1622C)
);

ninexnine_unit ninexnine_unit_3063(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1C007),
				.b1(W1C017),
				.b2(W1C027),
				.b3(W1C107),
				.b4(W1C117),
				.b5(W1C127),
				.b6(W1C207),
				.b7(W1C217),
				.b8(W1C227),
				.c(c1722C)
);

ninexnine_unit ninexnine_unit_3064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1C008),
				.b1(W1C018),
				.b2(W1C028),
				.b3(W1C108),
				.b4(W1C118),
				.b5(W1C128),
				.b6(W1C208),
				.b7(W1C218),
				.b8(W1C228),
				.c(c1822C)
);

ninexnine_unit ninexnine_unit_3065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1C009),
				.b1(W1C019),
				.b2(W1C029),
				.b3(W1C109),
				.b4(W1C119),
				.b5(W1C129),
				.b6(W1C209),
				.b7(W1C219),
				.b8(W1C229),
				.c(c1922C)
);

ninexnine_unit ninexnine_unit_3066(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1C00A),
				.b1(W1C01A),
				.b2(W1C02A),
				.b3(W1C10A),
				.b4(W1C11A),
				.b5(W1C12A),
				.b6(W1C20A),
				.b7(W1C21A),
				.b8(W1C22A),
				.c(c1A22C)
);

ninexnine_unit ninexnine_unit_3067(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1C00B),
				.b1(W1C01B),
				.b2(W1C02B),
				.b3(W1C10B),
				.b4(W1C11B),
				.b5(W1C12B),
				.b6(W1C20B),
				.b7(W1C21B),
				.b8(W1C22B),
				.c(c1B22C)
);

ninexnine_unit ninexnine_unit_3068(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1C00C),
				.b1(W1C01C),
				.b2(W1C02C),
				.b3(W1C10C),
				.b4(W1C11C),
				.b5(W1C12C),
				.b6(W1C20C),
				.b7(W1C21C),
				.b8(W1C22C),
				.c(c1C22C)
);

ninexnine_unit ninexnine_unit_3069(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1C00D),
				.b1(W1C01D),
				.b2(W1C02D),
				.b3(W1C10D),
				.b4(W1C11D),
				.b5(W1C12D),
				.b6(W1C20D),
				.b7(W1C21D),
				.b8(W1C22D),
				.c(c1D22C)
);

ninexnine_unit ninexnine_unit_3070(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1C00E),
				.b1(W1C01E),
				.b2(W1C02E),
				.b3(W1C10E),
				.b4(W1C11E),
				.b5(W1C12E),
				.b6(W1C20E),
				.b7(W1C21E),
				.b8(W1C22E),
				.c(c1E22C)
);

ninexnine_unit ninexnine_unit_3071(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1C00F),
				.b1(W1C01F),
				.b2(W1C02F),
				.b3(W1C10F),
				.b4(W1C11F),
				.b5(W1C12F),
				.b6(W1C20F),
				.b7(W1C21F),
				.b8(W1C22F),
				.c(c1F22C)
);

assign C122C=c1022C+c1122C+c1222C+c1322C+c1422C+c1522C+c1622C+c1722C+c1822C+c1922C+c1A22C+c1B22C+c1C22C+c1D22C+c1E22C+c1F22C;
assign A122C=(C122C>=0)?1:0;

assign P222C=A122C;

ninexnine_unit ninexnine_unit_3072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1000D)
);

ninexnine_unit ninexnine_unit_3073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1100D)
);

ninexnine_unit ninexnine_unit_3074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1200D)
);

ninexnine_unit ninexnine_unit_3075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1300D)
);

ninexnine_unit ninexnine_unit_3076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1400D)
);

ninexnine_unit ninexnine_unit_3077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1500D)
);

ninexnine_unit ninexnine_unit_3078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1600D)
);

ninexnine_unit ninexnine_unit_3079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1700D)
);

ninexnine_unit ninexnine_unit_3080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1800D)
);

ninexnine_unit ninexnine_unit_3081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1900D)
);

ninexnine_unit ninexnine_unit_3082(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A00D)
);

ninexnine_unit ninexnine_unit_3083(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B00D)
);

ninexnine_unit ninexnine_unit_3084(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C00D)
);

ninexnine_unit ninexnine_unit_3085(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D00D)
);

ninexnine_unit ninexnine_unit_3086(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E00D)
);

ninexnine_unit ninexnine_unit_3087(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F00D)
);

assign C100D=c1000D+c1100D+c1200D+c1300D+c1400D+c1500D+c1600D+c1700D+c1800D+c1900D+c1A00D+c1B00D+c1C00D+c1D00D+c1E00D+c1F00D;
assign A100D=(C100D>=0)?1:0;

assign P200D=A100D;

ninexnine_unit ninexnine_unit_3088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1001D)
);

ninexnine_unit ninexnine_unit_3089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1101D)
);

ninexnine_unit ninexnine_unit_3090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1201D)
);

ninexnine_unit ninexnine_unit_3091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1301D)
);

ninexnine_unit ninexnine_unit_3092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1401D)
);

ninexnine_unit ninexnine_unit_3093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1501D)
);

ninexnine_unit ninexnine_unit_3094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1601D)
);

ninexnine_unit ninexnine_unit_3095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1701D)
);

ninexnine_unit ninexnine_unit_3096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1801D)
);

ninexnine_unit ninexnine_unit_3097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1901D)
);

ninexnine_unit ninexnine_unit_3098(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A01D)
);

ninexnine_unit ninexnine_unit_3099(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B01D)
);

ninexnine_unit ninexnine_unit_3100(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C01D)
);

ninexnine_unit ninexnine_unit_3101(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D01D)
);

ninexnine_unit ninexnine_unit_3102(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E01D)
);

ninexnine_unit ninexnine_unit_3103(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F01D)
);

assign C101D=c1001D+c1101D+c1201D+c1301D+c1401D+c1501D+c1601D+c1701D+c1801D+c1901D+c1A01D+c1B01D+c1C01D+c1D01D+c1E01D+c1F01D;
assign A101D=(C101D>=0)?1:0;

assign P201D=A101D;

ninexnine_unit ninexnine_unit_3104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1002D)
);

ninexnine_unit ninexnine_unit_3105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1102D)
);

ninexnine_unit ninexnine_unit_3106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1202D)
);

ninexnine_unit ninexnine_unit_3107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1302D)
);

ninexnine_unit ninexnine_unit_3108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1402D)
);

ninexnine_unit ninexnine_unit_3109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1502D)
);

ninexnine_unit ninexnine_unit_3110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1602D)
);

ninexnine_unit ninexnine_unit_3111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1702D)
);

ninexnine_unit ninexnine_unit_3112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1802D)
);

ninexnine_unit ninexnine_unit_3113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1902D)
);

ninexnine_unit ninexnine_unit_3114(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A02D)
);

ninexnine_unit ninexnine_unit_3115(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B02D)
);

ninexnine_unit ninexnine_unit_3116(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C02D)
);

ninexnine_unit ninexnine_unit_3117(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D02D)
);

ninexnine_unit ninexnine_unit_3118(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E02D)
);

ninexnine_unit ninexnine_unit_3119(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F02D)
);

assign C102D=c1002D+c1102D+c1202D+c1302D+c1402D+c1502D+c1602D+c1702D+c1802D+c1902D+c1A02D+c1B02D+c1C02D+c1D02D+c1E02D+c1F02D;
assign A102D=(C102D>=0)?1:0;

assign P202D=A102D;

ninexnine_unit ninexnine_unit_3120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1010D)
);

ninexnine_unit ninexnine_unit_3121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1110D)
);

ninexnine_unit ninexnine_unit_3122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1210D)
);

ninexnine_unit ninexnine_unit_3123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1310D)
);

ninexnine_unit ninexnine_unit_3124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1410D)
);

ninexnine_unit ninexnine_unit_3125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1510D)
);

ninexnine_unit ninexnine_unit_3126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1610D)
);

ninexnine_unit ninexnine_unit_3127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1710D)
);

ninexnine_unit ninexnine_unit_3128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1810D)
);

ninexnine_unit ninexnine_unit_3129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1910D)
);

ninexnine_unit ninexnine_unit_3130(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A10D)
);

ninexnine_unit ninexnine_unit_3131(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B10D)
);

ninexnine_unit ninexnine_unit_3132(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C10D)
);

ninexnine_unit ninexnine_unit_3133(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D10D)
);

ninexnine_unit ninexnine_unit_3134(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E10D)
);

ninexnine_unit ninexnine_unit_3135(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F10D)
);

assign C110D=c1010D+c1110D+c1210D+c1310D+c1410D+c1510D+c1610D+c1710D+c1810D+c1910D+c1A10D+c1B10D+c1C10D+c1D10D+c1E10D+c1F10D;
assign A110D=(C110D>=0)?1:0;

assign P210D=A110D;

ninexnine_unit ninexnine_unit_3136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1011D)
);

ninexnine_unit ninexnine_unit_3137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1111D)
);

ninexnine_unit ninexnine_unit_3138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1211D)
);

ninexnine_unit ninexnine_unit_3139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1311D)
);

ninexnine_unit ninexnine_unit_3140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1411D)
);

ninexnine_unit ninexnine_unit_3141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1511D)
);

ninexnine_unit ninexnine_unit_3142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1611D)
);

ninexnine_unit ninexnine_unit_3143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1711D)
);

ninexnine_unit ninexnine_unit_3144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1811D)
);

ninexnine_unit ninexnine_unit_3145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1911D)
);

ninexnine_unit ninexnine_unit_3146(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A11D)
);

ninexnine_unit ninexnine_unit_3147(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B11D)
);

ninexnine_unit ninexnine_unit_3148(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C11D)
);

ninexnine_unit ninexnine_unit_3149(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D11D)
);

ninexnine_unit ninexnine_unit_3150(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E11D)
);

ninexnine_unit ninexnine_unit_3151(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F11D)
);

assign C111D=c1011D+c1111D+c1211D+c1311D+c1411D+c1511D+c1611D+c1711D+c1811D+c1911D+c1A11D+c1B11D+c1C11D+c1D11D+c1E11D+c1F11D;
assign A111D=(C111D>=0)?1:0;

assign P211D=A111D;

ninexnine_unit ninexnine_unit_3152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1012D)
);

ninexnine_unit ninexnine_unit_3153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1112D)
);

ninexnine_unit ninexnine_unit_3154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1212D)
);

ninexnine_unit ninexnine_unit_3155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1312D)
);

ninexnine_unit ninexnine_unit_3156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1412D)
);

ninexnine_unit ninexnine_unit_3157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1512D)
);

ninexnine_unit ninexnine_unit_3158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1612D)
);

ninexnine_unit ninexnine_unit_3159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1712D)
);

ninexnine_unit ninexnine_unit_3160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1812D)
);

ninexnine_unit ninexnine_unit_3161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1912D)
);

ninexnine_unit ninexnine_unit_3162(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A12D)
);

ninexnine_unit ninexnine_unit_3163(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B12D)
);

ninexnine_unit ninexnine_unit_3164(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C12D)
);

ninexnine_unit ninexnine_unit_3165(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D12D)
);

ninexnine_unit ninexnine_unit_3166(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E12D)
);

ninexnine_unit ninexnine_unit_3167(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F12D)
);

assign C112D=c1012D+c1112D+c1212D+c1312D+c1412D+c1512D+c1612D+c1712D+c1812D+c1912D+c1A12D+c1B12D+c1C12D+c1D12D+c1E12D+c1F12D;
assign A112D=(C112D>=0)?1:0;

assign P212D=A112D;

ninexnine_unit ninexnine_unit_3168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1020D)
);

ninexnine_unit ninexnine_unit_3169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1120D)
);

ninexnine_unit ninexnine_unit_3170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1220D)
);

ninexnine_unit ninexnine_unit_3171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1320D)
);

ninexnine_unit ninexnine_unit_3172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1420D)
);

ninexnine_unit ninexnine_unit_3173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1520D)
);

ninexnine_unit ninexnine_unit_3174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1620D)
);

ninexnine_unit ninexnine_unit_3175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1720D)
);

ninexnine_unit ninexnine_unit_3176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1820D)
);

ninexnine_unit ninexnine_unit_3177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1920D)
);

ninexnine_unit ninexnine_unit_3178(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A20D)
);

ninexnine_unit ninexnine_unit_3179(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B20D)
);

ninexnine_unit ninexnine_unit_3180(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C20D)
);

ninexnine_unit ninexnine_unit_3181(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D20D)
);

ninexnine_unit ninexnine_unit_3182(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E20D)
);

ninexnine_unit ninexnine_unit_3183(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F20D)
);

assign C120D=c1020D+c1120D+c1220D+c1320D+c1420D+c1520D+c1620D+c1720D+c1820D+c1920D+c1A20D+c1B20D+c1C20D+c1D20D+c1E20D+c1F20D;
assign A120D=(C120D>=0)?1:0;

assign P220D=A120D;

ninexnine_unit ninexnine_unit_3184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1021D)
);

ninexnine_unit ninexnine_unit_3185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1121D)
);

ninexnine_unit ninexnine_unit_3186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1221D)
);

ninexnine_unit ninexnine_unit_3187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1321D)
);

ninexnine_unit ninexnine_unit_3188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1421D)
);

ninexnine_unit ninexnine_unit_3189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1521D)
);

ninexnine_unit ninexnine_unit_3190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1621D)
);

ninexnine_unit ninexnine_unit_3191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1721D)
);

ninexnine_unit ninexnine_unit_3192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1821D)
);

ninexnine_unit ninexnine_unit_3193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1921D)
);

ninexnine_unit ninexnine_unit_3194(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A21D)
);

ninexnine_unit ninexnine_unit_3195(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B21D)
);

ninexnine_unit ninexnine_unit_3196(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C21D)
);

ninexnine_unit ninexnine_unit_3197(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D21D)
);

ninexnine_unit ninexnine_unit_3198(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E21D)
);

ninexnine_unit ninexnine_unit_3199(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F21D)
);

assign C121D=c1021D+c1121D+c1221D+c1321D+c1421D+c1521D+c1621D+c1721D+c1821D+c1921D+c1A21D+c1B21D+c1C21D+c1D21D+c1E21D+c1F21D;
assign A121D=(C121D>=0)?1:0;

assign P221D=A121D;

ninexnine_unit ninexnine_unit_3200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1022D)
);

ninexnine_unit ninexnine_unit_3201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1122D)
);

ninexnine_unit ninexnine_unit_3202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1222D)
);

ninexnine_unit ninexnine_unit_3203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1D003),
				.b1(W1D013),
				.b2(W1D023),
				.b3(W1D103),
				.b4(W1D113),
				.b5(W1D123),
				.b6(W1D203),
				.b7(W1D213),
				.b8(W1D223),
				.c(c1322D)
);

ninexnine_unit ninexnine_unit_3204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1D004),
				.b1(W1D014),
				.b2(W1D024),
				.b3(W1D104),
				.b4(W1D114),
				.b5(W1D124),
				.b6(W1D204),
				.b7(W1D214),
				.b8(W1D224),
				.c(c1422D)
);

ninexnine_unit ninexnine_unit_3205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1D005),
				.b1(W1D015),
				.b2(W1D025),
				.b3(W1D105),
				.b4(W1D115),
				.b5(W1D125),
				.b6(W1D205),
				.b7(W1D215),
				.b8(W1D225),
				.c(c1522D)
);

ninexnine_unit ninexnine_unit_3206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1D006),
				.b1(W1D016),
				.b2(W1D026),
				.b3(W1D106),
				.b4(W1D116),
				.b5(W1D126),
				.b6(W1D206),
				.b7(W1D216),
				.b8(W1D226),
				.c(c1622D)
);

ninexnine_unit ninexnine_unit_3207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1D007),
				.b1(W1D017),
				.b2(W1D027),
				.b3(W1D107),
				.b4(W1D117),
				.b5(W1D127),
				.b6(W1D207),
				.b7(W1D217),
				.b8(W1D227),
				.c(c1722D)
);

ninexnine_unit ninexnine_unit_3208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1D008),
				.b1(W1D018),
				.b2(W1D028),
				.b3(W1D108),
				.b4(W1D118),
				.b5(W1D128),
				.b6(W1D208),
				.b7(W1D218),
				.b8(W1D228),
				.c(c1822D)
);

ninexnine_unit ninexnine_unit_3209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1D009),
				.b1(W1D019),
				.b2(W1D029),
				.b3(W1D109),
				.b4(W1D119),
				.b5(W1D129),
				.b6(W1D209),
				.b7(W1D219),
				.b8(W1D229),
				.c(c1922D)
);

ninexnine_unit ninexnine_unit_3210(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1D00A),
				.b1(W1D01A),
				.b2(W1D02A),
				.b3(W1D10A),
				.b4(W1D11A),
				.b5(W1D12A),
				.b6(W1D20A),
				.b7(W1D21A),
				.b8(W1D22A),
				.c(c1A22D)
);

ninexnine_unit ninexnine_unit_3211(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1D00B),
				.b1(W1D01B),
				.b2(W1D02B),
				.b3(W1D10B),
				.b4(W1D11B),
				.b5(W1D12B),
				.b6(W1D20B),
				.b7(W1D21B),
				.b8(W1D22B),
				.c(c1B22D)
);

ninexnine_unit ninexnine_unit_3212(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1D00C),
				.b1(W1D01C),
				.b2(W1D02C),
				.b3(W1D10C),
				.b4(W1D11C),
				.b5(W1D12C),
				.b6(W1D20C),
				.b7(W1D21C),
				.b8(W1D22C),
				.c(c1C22D)
);

ninexnine_unit ninexnine_unit_3213(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1D00D),
				.b1(W1D01D),
				.b2(W1D02D),
				.b3(W1D10D),
				.b4(W1D11D),
				.b5(W1D12D),
				.b6(W1D20D),
				.b7(W1D21D),
				.b8(W1D22D),
				.c(c1D22D)
);

ninexnine_unit ninexnine_unit_3214(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1D00E),
				.b1(W1D01E),
				.b2(W1D02E),
				.b3(W1D10E),
				.b4(W1D11E),
				.b5(W1D12E),
				.b6(W1D20E),
				.b7(W1D21E),
				.b8(W1D22E),
				.c(c1E22D)
);

ninexnine_unit ninexnine_unit_3215(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1D00F),
				.b1(W1D01F),
				.b2(W1D02F),
				.b3(W1D10F),
				.b4(W1D11F),
				.b5(W1D12F),
				.b6(W1D20F),
				.b7(W1D21F),
				.b8(W1D22F),
				.c(c1F22D)
);

assign C122D=c1022D+c1122D+c1222D+c1322D+c1422D+c1522D+c1622D+c1722D+c1822D+c1922D+c1A22D+c1B22D+c1C22D+c1D22D+c1E22D+c1F22D;
assign A122D=(C122D>=0)?1:0;

assign P222D=A122D;

ninexnine_unit ninexnine_unit_3216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1000E)
);

ninexnine_unit ninexnine_unit_3217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1100E)
);

ninexnine_unit ninexnine_unit_3218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1200E)
);

ninexnine_unit ninexnine_unit_3219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1300E)
);

ninexnine_unit ninexnine_unit_3220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1400E)
);

ninexnine_unit ninexnine_unit_3221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1500E)
);

ninexnine_unit ninexnine_unit_3222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1600E)
);

ninexnine_unit ninexnine_unit_3223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1700E)
);

ninexnine_unit ninexnine_unit_3224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1800E)
);

ninexnine_unit ninexnine_unit_3225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1900E)
);

ninexnine_unit ninexnine_unit_3226(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A00E)
);

ninexnine_unit ninexnine_unit_3227(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B00E)
);

ninexnine_unit ninexnine_unit_3228(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C00E)
);

ninexnine_unit ninexnine_unit_3229(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D00E)
);

ninexnine_unit ninexnine_unit_3230(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E00E)
);

ninexnine_unit ninexnine_unit_3231(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F00E)
);

assign C100E=c1000E+c1100E+c1200E+c1300E+c1400E+c1500E+c1600E+c1700E+c1800E+c1900E+c1A00E+c1B00E+c1C00E+c1D00E+c1E00E+c1F00E;
assign A100E=(C100E>=0)?1:0;

assign P200E=A100E;

ninexnine_unit ninexnine_unit_3232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1001E)
);

ninexnine_unit ninexnine_unit_3233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1101E)
);

ninexnine_unit ninexnine_unit_3234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1201E)
);

ninexnine_unit ninexnine_unit_3235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1301E)
);

ninexnine_unit ninexnine_unit_3236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1401E)
);

ninexnine_unit ninexnine_unit_3237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1501E)
);

ninexnine_unit ninexnine_unit_3238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1601E)
);

ninexnine_unit ninexnine_unit_3239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1701E)
);

ninexnine_unit ninexnine_unit_3240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1801E)
);

ninexnine_unit ninexnine_unit_3241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1901E)
);

ninexnine_unit ninexnine_unit_3242(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A01E)
);

ninexnine_unit ninexnine_unit_3243(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B01E)
);

ninexnine_unit ninexnine_unit_3244(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C01E)
);

ninexnine_unit ninexnine_unit_3245(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D01E)
);

ninexnine_unit ninexnine_unit_3246(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E01E)
);

ninexnine_unit ninexnine_unit_3247(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F01E)
);

assign C101E=c1001E+c1101E+c1201E+c1301E+c1401E+c1501E+c1601E+c1701E+c1801E+c1901E+c1A01E+c1B01E+c1C01E+c1D01E+c1E01E+c1F01E;
assign A101E=(C101E>=0)?1:0;

assign P201E=A101E;

ninexnine_unit ninexnine_unit_3248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1002E)
);

ninexnine_unit ninexnine_unit_3249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1102E)
);

ninexnine_unit ninexnine_unit_3250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1202E)
);

ninexnine_unit ninexnine_unit_3251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1302E)
);

ninexnine_unit ninexnine_unit_3252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1402E)
);

ninexnine_unit ninexnine_unit_3253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1502E)
);

ninexnine_unit ninexnine_unit_3254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1602E)
);

ninexnine_unit ninexnine_unit_3255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1702E)
);

ninexnine_unit ninexnine_unit_3256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1802E)
);

ninexnine_unit ninexnine_unit_3257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1902E)
);

ninexnine_unit ninexnine_unit_3258(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A02E)
);

ninexnine_unit ninexnine_unit_3259(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B02E)
);

ninexnine_unit ninexnine_unit_3260(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C02E)
);

ninexnine_unit ninexnine_unit_3261(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D02E)
);

ninexnine_unit ninexnine_unit_3262(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E02E)
);

ninexnine_unit ninexnine_unit_3263(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F02E)
);

assign C102E=c1002E+c1102E+c1202E+c1302E+c1402E+c1502E+c1602E+c1702E+c1802E+c1902E+c1A02E+c1B02E+c1C02E+c1D02E+c1E02E+c1F02E;
assign A102E=(C102E>=0)?1:0;

assign P202E=A102E;

ninexnine_unit ninexnine_unit_3264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1010E)
);

ninexnine_unit ninexnine_unit_3265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1110E)
);

ninexnine_unit ninexnine_unit_3266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1210E)
);

ninexnine_unit ninexnine_unit_3267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1310E)
);

ninexnine_unit ninexnine_unit_3268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1410E)
);

ninexnine_unit ninexnine_unit_3269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1510E)
);

ninexnine_unit ninexnine_unit_3270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1610E)
);

ninexnine_unit ninexnine_unit_3271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1710E)
);

ninexnine_unit ninexnine_unit_3272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1810E)
);

ninexnine_unit ninexnine_unit_3273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1910E)
);

ninexnine_unit ninexnine_unit_3274(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A10E)
);

ninexnine_unit ninexnine_unit_3275(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B10E)
);

ninexnine_unit ninexnine_unit_3276(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C10E)
);

ninexnine_unit ninexnine_unit_3277(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D10E)
);

ninexnine_unit ninexnine_unit_3278(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E10E)
);

ninexnine_unit ninexnine_unit_3279(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F10E)
);

assign C110E=c1010E+c1110E+c1210E+c1310E+c1410E+c1510E+c1610E+c1710E+c1810E+c1910E+c1A10E+c1B10E+c1C10E+c1D10E+c1E10E+c1F10E;
assign A110E=(C110E>=0)?1:0;

assign P210E=A110E;

ninexnine_unit ninexnine_unit_3280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1011E)
);

ninexnine_unit ninexnine_unit_3281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1111E)
);

ninexnine_unit ninexnine_unit_3282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1211E)
);

ninexnine_unit ninexnine_unit_3283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1311E)
);

ninexnine_unit ninexnine_unit_3284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1411E)
);

ninexnine_unit ninexnine_unit_3285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1511E)
);

ninexnine_unit ninexnine_unit_3286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1611E)
);

ninexnine_unit ninexnine_unit_3287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1711E)
);

ninexnine_unit ninexnine_unit_3288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1811E)
);

ninexnine_unit ninexnine_unit_3289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1911E)
);

ninexnine_unit ninexnine_unit_3290(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A11E)
);

ninexnine_unit ninexnine_unit_3291(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B11E)
);

ninexnine_unit ninexnine_unit_3292(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C11E)
);

ninexnine_unit ninexnine_unit_3293(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D11E)
);

ninexnine_unit ninexnine_unit_3294(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E11E)
);

ninexnine_unit ninexnine_unit_3295(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F11E)
);

assign C111E=c1011E+c1111E+c1211E+c1311E+c1411E+c1511E+c1611E+c1711E+c1811E+c1911E+c1A11E+c1B11E+c1C11E+c1D11E+c1E11E+c1F11E;
assign A111E=(C111E>=0)?1:0;

assign P211E=A111E;

ninexnine_unit ninexnine_unit_3296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1012E)
);

ninexnine_unit ninexnine_unit_3297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1112E)
);

ninexnine_unit ninexnine_unit_3298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1212E)
);

ninexnine_unit ninexnine_unit_3299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1312E)
);

ninexnine_unit ninexnine_unit_3300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1412E)
);

ninexnine_unit ninexnine_unit_3301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1512E)
);

ninexnine_unit ninexnine_unit_3302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1612E)
);

ninexnine_unit ninexnine_unit_3303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1712E)
);

ninexnine_unit ninexnine_unit_3304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1812E)
);

ninexnine_unit ninexnine_unit_3305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1912E)
);

ninexnine_unit ninexnine_unit_3306(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A12E)
);

ninexnine_unit ninexnine_unit_3307(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B12E)
);

ninexnine_unit ninexnine_unit_3308(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C12E)
);

ninexnine_unit ninexnine_unit_3309(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D12E)
);

ninexnine_unit ninexnine_unit_3310(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E12E)
);

ninexnine_unit ninexnine_unit_3311(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F12E)
);

assign C112E=c1012E+c1112E+c1212E+c1312E+c1412E+c1512E+c1612E+c1712E+c1812E+c1912E+c1A12E+c1B12E+c1C12E+c1D12E+c1E12E+c1F12E;
assign A112E=(C112E>=0)?1:0;

assign P212E=A112E;

ninexnine_unit ninexnine_unit_3312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1020E)
);

ninexnine_unit ninexnine_unit_3313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1120E)
);

ninexnine_unit ninexnine_unit_3314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1220E)
);

ninexnine_unit ninexnine_unit_3315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1320E)
);

ninexnine_unit ninexnine_unit_3316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1420E)
);

ninexnine_unit ninexnine_unit_3317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1520E)
);

ninexnine_unit ninexnine_unit_3318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1620E)
);

ninexnine_unit ninexnine_unit_3319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1720E)
);

ninexnine_unit ninexnine_unit_3320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1820E)
);

ninexnine_unit ninexnine_unit_3321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1920E)
);

ninexnine_unit ninexnine_unit_3322(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A20E)
);

ninexnine_unit ninexnine_unit_3323(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B20E)
);

ninexnine_unit ninexnine_unit_3324(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C20E)
);

ninexnine_unit ninexnine_unit_3325(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D20E)
);

ninexnine_unit ninexnine_unit_3326(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E20E)
);

ninexnine_unit ninexnine_unit_3327(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F20E)
);

assign C120E=c1020E+c1120E+c1220E+c1320E+c1420E+c1520E+c1620E+c1720E+c1820E+c1920E+c1A20E+c1B20E+c1C20E+c1D20E+c1E20E+c1F20E;
assign A120E=(C120E>=0)?1:0;

assign P220E=A120E;

ninexnine_unit ninexnine_unit_3328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1021E)
);

ninexnine_unit ninexnine_unit_3329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1121E)
);

ninexnine_unit ninexnine_unit_3330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1221E)
);

ninexnine_unit ninexnine_unit_3331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1321E)
);

ninexnine_unit ninexnine_unit_3332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1421E)
);

ninexnine_unit ninexnine_unit_3333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1521E)
);

ninexnine_unit ninexnine_unit_3334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1621E)
);

ninexnine_unit ninexnine_unit_3335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1721E)
);

ninexnine_unit ninexnine_unit_3336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1821E)
);

ninexnine_unit ninexnine_unit_3337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1921E)
);

ninexnine_unit ninexnine_unit_3338(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A21E)
);

ninexnine_unit ninexnine_unit_3339(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B21E)
);

ninexnine_unit ninexnine_unit_3340(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C21E)
);

ninexnine_unit ninexnine_unit_3341(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D21E)
);

ninexnine_unit ninexnine_unit_3342(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E21E)
);

ninexnine_unit ninexnine_unit_3343(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F21E)
);

assign C121E=c1021E+c1121E+c1221E+c1321E+c1421E+c1521E+c1621E+c1721E+c1821E+c1921E+c1A21E+c1B21E+c1C21E+c1D21E+c1E21E+c1F21E;
assign A121E=(C121E>=0)?1:0;

assign P221E=A121E;

ninexnine_unit ninexnine_unit_3344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1022E)
);

ninexnine_unit ninexnine_unit_3345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1122E)
);

ninexnine_unit ninexnine_unit_3346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1222E)
);

ninexnine_unit ninexnine_unit_3347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1E003),
				.b1(W1E013),
				.b2(W1E023),
				.b3(W1E103),
				.b4(W1E113),
				.b5(W1E123),
				.b6(W1E203),
				.b7(W1E213),
				.b8(W1E223),
				.c(c1322E)
);

ninexnine_unit ninexnine_unit_3348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1E004),
				.b1(W1E014),
				.b2(W1E024),
				.b3(W1E104),
				.b4(W1E114),
				.b5(W1E124),
				.b6(W1E204),
				.b7(W1E214),
				.b8(W1E224),
				.c(c1422E)
);

ninexnine_unit ninexnine_unit_3349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1E005),
				.b1(W1E015),
				.b2(W1E025),
				.b3(W1E105),
				.b4(W1E115),
				.b5(W1E125),
				.b6(W1E205),
				.b7(W1E215),
				.b8(W1E225),
				.c(c1522E)
);

ninexnine_unit ninexnine_unit_3350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1E006),
				.b1(W1E016),
				.b2(W1E026),
				.b3(W1E106),
				.b4(W1E116),
				.b5(W1E126),
				.b6(W1E206),
				.b7(W1E216),
				.b8(W1E226),
				.c(c1622E)
);

ninexnine_unit ninexnine_unit_3351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1E007),
				.b1(W1E017),
				.b2(W1E027),
				.b3(W1E107),
				.b4(W1E117),
				.b5(W1E127),
				.b6(W1E207),
				.b7(W1E217),
				.b8(W1E227),
				.c(c1722E)
);

ninexnine_unit ninexnine_unit_3352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1E008),
				.b1(W1E018),
				.b2(W1E028),
				.b3(W1E108),
				.b4(W1E118),
				.b5(W1E128),
				.b6(W1E208),
				.b7(W1E218),
				.b8(W1E228),
				.c(c1822E)
);

ninexnine_unit ninexnine_unit_3353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1E009),
				.b1(W1E019),
				.b2(W1E029),
				.b3(W1E109),
				.b4(W1E119),
				.b5(W1E129),
				.b6(W1E209),
				.b7(W1E219),
				.b8(W1E229),
				.c(c1922E)
);

ninexnine_unit ninexnine_unit_3354(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1E00A),
				.b1(W1E01A),
				.b2(W1E02A),
				.b3(W1E10A),
				.b4(W1E11A),
				.b5(W1E12A),
				.b6(W1E20A),
				.b7(W1E21A),
				.b8(W1E22A),
				.c(c1A22E)
);

ninexnine_unit ninexnine_unit_3355(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1E00B),
				.b1(W1E01B),
				.b2(W1E02B),
				.b3(W1E10B),
				.b4(W1E11B),
				.b5(W1E12B),
				.b6(W1E20B),
				.b7(W1E21B),
				.b8(W1E22B),
				.c(c1B22E)
);

ninexnine_unit ninexnine_unit_3356(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1E00C),
				.b1(W1E01C),
				.b2(W1E02C),
				.b3(W1E10C),
				.b4(W1E11C),
				.b5(W1E12C),
				.b6(W1E20C),
				.b7(W1E21C),
				.b8(W1E22C),
				.c(c1C22E)
);

ninexnine_unit ninexnine_unit_3357(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1E00D),
				.b1(W1E01D),
				.b2(W1E02D),
				.b3(W1E10D),
				.b4(W1E11D),
				.b5(W1E12D),
				.b6(W1E20D),
				.b7(W1E21D),
				.b8(W1E22D),
				.c(c1D22E)
);

ninexnine_unit ninexnine_unit_3358(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1E00E),
				.b1(W1E01E),
				.b2(W1E02E),
				.b3(W1E10E),
				.b4(W1E11E),
				.b5(W1E12E),
				.b6(W1E20E),
				.b7(W1E21E),
				.b8(W1E22E),
				.c(c1E22E)
);

ninexnine_unit ninexnine_unit_3359(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1E00F),
				.b1(W1E01F),
				.b2(W1E02F),
				.b3(W1E10F),
				.b4(W1E11F),
				.b5(W1E12F),
				.b6(W1E20F),
				.b7(W1E21F),
				.b8(W1E22F),
				.c(c1F22E)
);

assign C122E=c1022E+c1122E+c1222E+c1322E+c1422E+c1522E+c1622E+c1722E+c1822E+c1922E+c1A22E+c1B22E+c1C22E+c1D22E+c1E22E+c1F22E;
assign A122E=(C122E>=0)?1:0;

assign P222E=A122E;

ninexnine_unit ninexnine_unit_3360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1000F)
);

ninexnine_unit ninexnine_unit_3361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1100F)
);

ninexnine_unit ninexnine_unit_3362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1200F)
);

ninexnine_unit ninexnine_unit_3363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1300F)
);

ninexnine_unit ninexnine_unit_3364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1400F)
);

ninexnine_unit ninexnine_unit_3365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1500F)
);

ninexnine_unit ninexnine_unit_3366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1600F)
);

ninexnine_unit ninexnine_unit_3367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1700F)
);

ninexnine_unit ninexnine_unit_3368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1800F)
);

ninexnine_unit ninexnine_unit_3369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1900F)
);

ninexnine_unit ninexnine_unit_3370(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A00F)
);

ninexnine_unit ninexnine_unit_3371(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B00F)
);

ninexnine_unit ninexnine_unit_3372(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C00F)
);

ninexnine_unit ninexnine_unit_3373(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D00F)
);

ninexnine_unit ninexnine_unit_3374(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E00F)
);

ninexnine_unit ninexnine_unit_3375(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F00F)
);

assign C100F=c1000F+c1100F+c1200F+c1300F+c1400F+c1500F+c1600F+c1700F+c1800F+c1900F+c1A00F+c1B00F+c1C00F+c1D00F+c1E00F+c1F00F;
assign A100F=(C100F>=0)?1:0;

assign P200F=A100F;

ninexnine_unit ninexnine_unit_3376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1001F)
);

ninexnine_unit ninexnine_unit_3377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1101F)
);

ninexnine_unit ninexnine_unit_3378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1201F)
);

ninexnine_unit ninexnine_unit_3379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1301F)
);

ninexnine_unit ninexnine_unit_3380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1401F)
);

ninexnine_unit ninexnine_unit_3381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1501F)
);

ninexnine_unit ninexnine_unit_3382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1601F)
);

ninexnine_unit ninexnine_unit_3383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1701F)
);

ninexnine_unit ninexnine_unit_3384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1801F)
);

ninexnine_unit ninexnine_unit_3385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1901F)
);

ninexnine_unit ninexnine_unit_3386(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A01F)
);

ninexnine_unit ninexnine_unit_3387(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B01F)
);

ninexnine_unit ninexnine_unit_3388(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C01F)
);

ninexnine_unit ninexnine_unit_3389(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D01F)
);

ninexnine_unit ninexnine_unit_3390(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E01F)
);

ninexnine_unit ninexnine_unit_3391(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F01F)
);

assign C101F=c1001F+c1101F+c1201F+c1301F+c1401F+c1501F+c1601F+c1701F+c1801F+c1901F+c1A01F+c1B01F+c1C01F+c1D01F+c1E01F+c1F01F;
assign A101F=(C101F>=0)?1:0;

assign P201F=A101F;

ninexnine_unit ninexnine_unit_3392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1002F)
);

ninexnine_unit ninexnine_unit_3393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1102F)
);

ninexnine_unit ninexnine_unit_3394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1202F)
);

ninexnine_unit ninexnine_unit_3395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1302F)
);

ninexnine_unit ninexnine_unit_3396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1402F)
);

ninexnine_unit ninexnine_unit_3397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1502F)
);

ninexnine_unit ninexnine_unit_3398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1602F)
);

ninexnine_unit ninexnine_unit_3399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1702F)
);

ninexnine_unit ninexnine_unit_3400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1802F)
);

ninexnine_unit ninexnine_unit_3401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1902F)
);

ninexnine_unit ninexnine_unit_3402(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A02F)
);

ninexnine_unit ninexnine_unit_3403(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B02F)
);

ninexnine_unit ninexnine_unit_3404(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C02F)
);

ninexnine_unit ninexnine_unit_3405(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D02F)
);

ninexnine_unit ninexnine_unit_3406(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E02F)
);

ninexnine_unit ninexnine_unit_3407(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F02F)
);

assign C102F=c1002F+c1102F+c1202F+c1302F+c1402F+c1502F+c1602F+c1702F+c1802F+c1902F+c1A02F+c1B02F+c1C02F+c1D02F+c1E02F+c1F02F;
assign A102F=(C102F>=0)?1:0;

assign P202F=A102F;

ninexnine_unit ninexnine_unit_3408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1010F)
);

ninexnine_unit ninexnine_unit_3409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1110F)
);

ninexnine_unit ninexnine_unit_3410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1210F)
);

ninexnine_unit ninexnine_unit_3411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1310F)
);

ninexnine_unit ninexnine_unit_3412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1410F)
);

ninexnine_unit ninexnine_unit_3413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1510F)
);

ninexnine_unit ninexnine_unit_3414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1610F)
);

ninexnine_unit ninexnine_unit_3415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1710F)
);

ninexnine_unit ninexnine_unit_3416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1810F)
);

ninexnine_unit ninexnine_unit_3417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1910F)
);

ninexnine_unit ninexnine_unit_3418(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A10F)
);

ninexnine_unit ninexnine_unit_3419(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B10F)
);

ninexnine_unit ninexnine_unit_3420(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C10F)
);

ninexnine_unit ninexnine_unit_3421(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D10F)
);

ninexnine_unit ninexnine_unit_3422(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E10F)
);

ninexnine_unit ninexnine_unit_3423(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F10F)
);

assign C110F=c1010F+c1110F+c1210F+c1310F+c1410F+c1510F+c1610F+c1710F+c1810F+c1910F+c1A10F+c1B10F+c1C10F+c1D10F+c1E10F+c1F10F;
assign A110F=(C110F>=0)?1:0;

assign P210F=A110F;

ninexnine_unit ninexnine_unit_3424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1011F)
);

ninexnine_unit ninexnine_unit_3425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1111F)
);

ninexnine_unit ninexnine_unit_3426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1211F)
);

ninexnine_unit ninexnine_unit_3427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1311F)
);

ninexnine_unit ninexnine_unit_3428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1411F)
);

ninexnine_unit ninexnine_unit_3429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1511F)
);

ninexnine_unit ninexnine_unit_3430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1611F)
);

ninexnine_unit ninexnine_unit_3431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1711F)
);

ninexnine_unit ninexnine_unit_3432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1811F)
);

ninexnine_unit ninexnine_unit_3433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1911F)
);

ninexnine_unit ninexnine_unit_3434(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A11F)
);

ninexnine_unit ninexnine_unit_3435(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B11F)
);

ninexnine_unit ninexnine_unit_3436(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C11F)
);

ninexnine_unit ninexnine_unit_3437(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D11F)
);

ninexnine_unit ninexnine_unit_3438(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E11F)
);

ninexnine_unit ninexnine_unit_3439(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F11F)
);

assign C111F=c1011F+c1111F+c1211F+c1311F+c1411F+c1511F+c1611F+c1711F+c1811F+c1911F+c1A11F+c1B11F+c1C11F+c1D11F+c1E11F+c1F11F;
assign A111F=(C111F>=0)?1:0;

assign P211F=A111F;

ninexnine_unit ninexnine_unit_3440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1012F)
);

ninexnine_unit ninexnine_unit_3441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1112F)
);

ninexnine_unit ninexnine_unit_3442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1212F)
);

ninexnine_unit ninexnine_unit_3443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1312F)
);

ninexnine_unit ninexnine_unit_3444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1412F)
);

ninexnine_unit ninexnine_unit_3445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1512F)
);

ninexnine_unit ninexnine_unit_3446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1612F)
);

ninexnine_unit ninexnine_unit_3447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1712F)
);

ninexnine_unit ninexnine_unit_3448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1812F)
);

ninexnine_unit ninexnine_unit_3449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1912F)
);

ninexnine_unit ninexnine_unit_3450(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A12F)
);

ninexnine_unit ninexnine_unit_3451(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B12F)
);

ninexnine_unit ninexnine_unit_3452(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C12F)
);

ninexnine_unit ninexnine_unit_3453(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D12F)
);

ninexnine_unit ninexnine_unit_3454(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E12F)
);

ninexnine_unit ninexnine_unit_3455(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F12F)
);

assign C112F=c1012F+c1112F+c1212F+c1312F+c1412F+c1512F+c1612F+c1712F+c1812F+c1912F+c1A12F+c1B12F+c1C12F+c1D12F+c1E12F+c1F12F;
assign A112F=(C112F>=0)?1:0;

assign P212F=A112F;

ninexnine_unit ninexnine_unit_3456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1020F)
);

ninexnine_unit ninexnine_unit_3457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1120F)
);

ninexnine_unit ninexnine_unit_3458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1220F)
);

ninexnine_unit ninexnine_unit_3459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1320F)
);

ninexnine_unit ninexnine_unit_3460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1420F)
);

ninexnine_unit ninexnine_unit_3461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1520F)
);

ninexnine_unit ninexnine_unit_3462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1620F)
);

ninexnine_unit ninexnine_unit_3463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1720F)
);

ninexnine_unit ninexnine_unit_3464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1820F)
);

ninexnine_unit ninexnine_unit_3465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1920F)
);

ninexnine_unit ninexnine_unit_3466(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A20F)
);

ninexnine_unit ninexnine_unit_3467(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B20F)
);

ninexnine_unit ninexnine_unit_3468(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C20F)
);

ninexnine_unit ninexnine_unit_3469(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D20F)
);

ninexnine_unit ninexnine_unit_3470(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E20F)
);

ninexnine_unit ninexnine_unit_3471(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F20F)
);

assign C120F=c1020F+c1120F+c1220F+c1320F+c1420F+c1520F+c1620F+c1720F+c1820F+c1920F+c1A20F+c1B20F+c1C20F+c1D20F+c1E20F+c1F20F;
assign A120F=(C120F>=0)?1:0;

assign P220F=A120F;

ninexnine_unit ninexnine_unit_3472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1021F)
);

ninexnine_unit ninexnine_unit_3473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1121F)
);

ninexnine_unit ninexnine_unit_3474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1221F)
);

ninexnine_unit ninexnine_unit_3475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1321F)
);

ninexnine_unit ninexnine_unit_3476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1421F)
);

ninexnine_unit ninexnine_unit_3477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1521F)
);

ninexnine_unit ninexnine_unit_3478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1621F)
);

ninexnine_unit ninexnine_unit_3479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1721F)
);

ninexnine_unit ninexnine_unit_3480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1821F)
);

ninexnine_unit ninexnine_unit_3481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1921F)
);

ninexnine_unit ninexnine_unit_3482(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A21F)
);

ninexnine_unit ninexnine_unit_3483(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B21F)
);

ninexnine_unit ninexnine_unit_3484(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C21F)
);

ninexnine_unit ninexnine_unit_3485(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D21F)
);

ninexnine_unit ninexnine_unit_3486(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E21F)
);

ninexnine_unit ninexnine_unit_3487(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F21F)
);

assign C121F=c1021F+c1121F+c1221F+c1321F+c1421F+c1521F+c1621F+c1721F+c1821F+c1921F+c1A21F+c1B21F+c1C21F+c1D21F+c1E21F+c1F21F;
assign A121F=(C121F>=0)?1:0;

assign P221F=A121F;

ninexnine_unit ninexnine_unit_3488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1022F)
);

ninexnine_unit ninexnine_unit_3489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1122F)
);

ninexnine_unit ninexnine_unit_3490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1222F)
);

ninexnine_unit ninexnine_unit_3491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1F003),
				.b1(W1F013),
				.b2(W1F023),
				.b3(W1F103),
				.b4(W1F113),
				.b5(W1F123),
				.b6(W1F203),
				.b7(W1F213),
				.b8(W1F223),
				.c(c1322F)
);

ninexnine_unit ninexnine_unit_3492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1F004),
				.b1(W1F014),
				.b2(W1F024),
				.b3(W1F104),
				.b4(W1F114),
				.b5(W1F124),
				.b6(W1F204),
				.b7(W1F214),
				.b8(W1F224),
				.c(c1422F)
);

ninexnine_unit ninexnine_unit_3493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1F005),
				.b1(W1F015),
				.b2(W1F025),
				.b3(W1F105),
				.b4(W1F115),
				.b5(W1F125),
				.b6(W1F205),
				.b7(W1F215),
				.b8(W1F225),
				.c(c1522F)
);

ninexnine_unit ninexnine_unit_3494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1F006),
				.b1(W1F016),
				.b2(W1F026),
				.b3(W1F106),
				.b4(W1F116),
				.b5(W1F126),
				.b6(W1F206),
				.b7(W1F216),
				.b8(W1F226),
				.c(c1622F)
);

ninexnine_unit ninexnine_unit_3495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1F007),
				.b1(W1F017),
				.b2(W1F027),
				.b3(W1F107),
				.b4(W1F117),
				.b5(W1F127),
				.b6(W1F207),
				.b7(W1F217),
				.b8(W1F227),
				.c(c1722F)
);

ninexnine_unit ninexnine_unit_3496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1F008),
				.b1(W1F018),
				.b2(W1F028),
				.b3(W1F108),
				.b4(W1F118),
				.b5(W1F128),
				.b6(W1F208),
				.b7(W1F218),
				.b8(W1F228),
				.c(c1822F)
);

ninexnine_unit ninexnine_unit_3497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1F009),
				.b1(W1F019),
				.b2(W1F029),
				.b3(W1F109),
				.b4(W1F119),
				.b5(W1F129),
				.b6(W1F209),
				.b7(W1F219),
				.b8(W1F229),
				.c(c1922F)
);

ninexnine_unit ninexnine_unit_3498(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1F00A),
				.b1(W1F01A),
				.b2(W1F02A),
				.b3(W1F10A),
				.b4(W1F11A),
				.b5(W1F12A),
				.b6(W1F20A),
				.b7(W1F21A),
				.b8(W1F22A),
				.c(c1A22F)
);

ninexnine_unit ninexnine_unit_3499(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1F00B),
				.b1(W1F01B),
				.b2(W1F02B),
				.b3(W1F10B),
				.b4(W1F11B),
				.b5(W1F12B),
				.b6(W1F20B),
				.b7(W1F21B),
				.b8(W1F22B),
				.c(c1B22F)
);

ninexnine_unit ninexnine_unit_3500(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1F00C),
				.b1(W1F01C),
				.b2(W1F02C),
				.b3(W1F10C),
				.b4(W1F11C),
				.b5(W1F12C),
				.b6(W1F20C),
				.b7(W1F21C),
				.b8(W1F22C),
				.c(c1C22F)
);

ninexnine_unit ninexnine_unit_3501(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1F00D),
				.b1(W1F01D),
				.b2(W1F02D),
				.b3(W1F10D),
				.b4(W1F11D),
				.b5(W1F12D),
				.b6(W1F20D),
				.b7(W1F21D),
				.b8(W1F22D),
				.c(c1D22F)
);

ninexnine_unit ninexnine_unit_3502(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1F00E),
				.b1(W1F01E),
				.b2(W1F02E),
				.b3(W1F10E),
				.b4(W1F11E),
				.b5(W1F12E),
				.b6(W1F20E),
				.b7(W1F21E),
				.b8(W1F22E),
				.c(c1E22F)
);

ninexnine_unit ninexnine_unit_3503(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1F00F),
				.b1(W1F01F),
				.b2(W1F02F),
				.b3(W1F10F),
				.b4(W1F11F),
				.b5(W1F12F),
				.b6(W1F20F),
				.b7(W1F21F),
				.b8(W1F22F),
				.c(c1F22F)
);

assign C122F=c1022F+c1122F+c1222F+c1322F+c1422F+c1522F+c1622F+c1722F+c1822F+c1922F+c1A22F+c1B22F+c1C22F+c1D22F+c1E22F+c1F22F;
assign A122F=(C122F>=0)?1:0;

assign P222F=A122F;

ninexnine_unit ninexnine_unit_3504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1000G)
);

ninexnine_unit ninexnine_unit_3505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1100G)
);

ninexnine_unit ninexnine_unit_3506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1200G)
);

ninexnine_unit ninexnine_unit_3507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1300G)
);

ninexnine_unit ninexnine_unit_3508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1400G)
);

ninexnine_unit ninexnine_unit_3509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1500G)
);

ninexnine_unit ninexnine_unit_3510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1600G)
);

ninexnine_unit ninexnine_unit_3511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1700G)
);

ninexnine_unit ninexnine_unit_3512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1800G)
);

ninexnine_unit ninexnine_unit_3513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1900G)
);

ninexnine_unit ninexnine_unit_3514(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A00G)
);

ninexnine_unit ninexnine_unit_3515(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B00G)
);

ninexnine_unit ninexnine_unit_3516(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C00G)
);

ninexnine_unit ninexnine_unit_3517(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D00G)
);

ninexnine_unit ninexnine_unit_3518(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E00G)
);

ninexnine_unit ninexnine_unit_3519(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F00G)
);

assign C100G=c1000G+c1100G+c1200G+c1300G+c1400G+c1500G+c1600G+c1700G+c1800G+c1900G+c1A00G+c1B00G+c1C00G+c1D00G+c1E00G+c1F00G;
assign A100G=(C100G>=0)?1:0;

assign P200G=A100G;

ninexnine_unit ninexnine_unit_3520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1001G)
);

ninexnine_unit ninexnine_unit_3521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1101G)
);

ninexnine_unit ninexnine_unit_3522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1201G)
);

ninexnine_unit ninexnine_unit_3523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1301G)
);

ninexnine_unit ninexnine_unit_3524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1401G)
);

ninexnine_unit ninexnine_unit_3525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1501G)
);

ninexnine_unit ninexnine_unit_3526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1601G)
);

ninexnine_unit ninexnine_unit_3527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1701G)
);

ninexnine_unit ninexnine_unit_3528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1801G)
);

ninexnine_unit ninexnine_unit_3529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1901G)
);

ninexnine_unit ninexnine_unit_3530(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A01G)
);

ninexnine_unit ninexnine_unit_3531(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B01G)
);

ninexnine_unit ninexnine_unit_3532(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C01G)
);

ninexnine_unit ninexnine_unit_3533(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D01G)
);

ninexnine_unit ninexnine_unit_3534(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E01G)
);

ninexnine_unit ninexnine_unit_3535(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F01G)
);

assign C101G=c1001G+c1101G+c1201G+c1301G+c1401G+c1501G+c1601G+c1701G+c1801G+c1901G+c1A01G+c1B01G+c1C01G+c1D01G+c1E01G+c1F01G;
assign A101G=(C101G>=0)?1:0;

assign P201G=A101G;

ninexnine_unit ninexnine_unit_3536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1002G)
);

ninexnine_unit ninexnine_unit_3537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1102G)
);

ninexnine_unit ninexnine_unit_3538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1202G)
);

ninexnine_unit ninexnine_unit_3539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1302G)
);

ninexnine_unit ninexnine_unit_3540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1402G)
);

ninexnine_unit ninexnine_unit_3541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1502G)
);

ninexnine_unit ninexnine_unit_3542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1602G)
);

ninexnine_unit ninexnine_unit_3543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1702G)
);

ninexnine_unit ninexnine_unit_3544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1802G)
);

ninexnine_unit ninexnine_unit_3545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1902G)
);

ninexnine_unit ninexnine_unit_3546(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A02G)
);

ninexnine_unit ninexnine_unit_3547(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B02G)
);

ninexnine_unit ninexnine_unit_3548(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C02G)
);

ninexnine_unit ninexnine_unit_3549(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D02G)
);

ninexnine_unit ninexnine_unit_3550(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E02G)
);

ninexnine_unit ninexnine_unit_3551(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F02G)
);

assign C102G=c1002G+c1102G+c1202G+c1302G+c1402G+c1502G+c1602G+c1702G+c1802G+c1902G+c1A02G+c1B02G+c1C02G+c1D02G+c1E02G+c1F02G;
assign A102G=(C102G>=0)?1:0;

assign P202G=A102G;

ninexnine_unit ninexnine_unit_3552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1010G)
);

ninexnine_unit ninexnine_unit_3553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1110G)
);

ninexnine_unit ninexnine_unit_3554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1210G)
);

ninexnine_unit ninexnine_unit_3555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1310G)
);

ninexnine_unit ninexnine_unit_3556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1410G)
);

ninexnine_unit ninexnine_unit_3557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1510G)
);

ninexnine_unit ninexnine_unit_3558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1610G)
);

ninexnine_unit ninexnine_unit_3559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1710G)
);

ninexnine_unit ninexnine_unit_3560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1810G)
);

ninexnine_unit ninexnine_unit_3561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1910G)
);

ninexnine_unit ninexnine_unit_3562(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A10G)
);

ninexnine_unit ninexnine_unit_3563(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B10G)
);

ninexnine_unit ninexnine_unit_3564(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C10G)
);

ninexnine_unit ninexnine_unit_3565(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D10G)
);

ninexnine_unit ninexnine_unit_3566(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E10G)
);

ninexnine_unit ninexnine_unit_3567(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F10G)
);

assign C110G=c1010G+c1110G+c1210G+c1310G+c1410G+c1510G+c1610G+c1710G+c1810G+c1910G+c1A10G+c1B10G+c1C10G+c1D10G+c1E10G+c1F10G;
assign A110G=(C110G>=0)?1:0;

assign P210G=A110G;

ninexnine_unit ninexnine_unit_3568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1011G)
);

ninexnine_unit ninexnine_unit_3569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1111G)
);

ninexnine_unit ninexnine_unit_3570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1211G)
);

ninexnine_unit ninexnine_unit_3571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1311G)
);

ninexnine_unit ninexnine_unit_3572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1411G)
);

ninexnine_unit ninexnine_unit_3573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1511G)
);

ninexnine_unit ninexnine_unit_3574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1611G)
);

ninexnine_unit ninexnine_unit_3575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1711G)
);

ninexnine_unit ninexnine_unit_3576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1811G)
);

ninexnine_unit ninexnine_unit_3577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1911G)
);

ninexnine_unit ninexnine_unit_3578(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A11G)
);

ninexnine_unit ninexnine_unit_3579(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B11G)
);

ninexnine_unit ninexnine_unit_3580(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C11G)
);

ninexnine_unit ninexnine_unit_3581(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D11G)
);

ninexnine_unit ninexnine_unit_3582(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E11G)
);

ninexnine_unit ninexnine_unit_3583(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F11G)
);

assign C111G=c1011G+c1111G+c1211G+c1311G+c1411G+c1511G+c1611G+c1711G+c1811G+c1911G+c1A11G+c1B11G+c1C11G+c1D11G+c1E11G+c1F11G;
assign A111G=(C111G>=0)?1:0;

assign P211G=A111G;

ninexnine_unit ninexnine_unit_3584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1012G)
);

ninexnine_unit ninexnine_unit_3585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1112G)
);

ninexnine_unit ninexnine_unit_3586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1212G)
);

ninexnine_unit ninexnine_unit_3587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1312G)
);

ninexnine_unit ninexnine_unit_3588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1412G)
);

ninexnine_unit ninexnine_unit_3589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1512G)
);

ninexnine_unit ninexnine_unit_3590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1612G)
);

ninexnine_unit ninexnine_unit_3591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1712G)
);

ninexnine_unit ninexnine_unit_3592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1812G)
);

ninexnine_unit ninexnine_unit_3593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1912G)
);

ninexnine_unit ninexnine_unit_3594(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A12G)
);

ninexnine_unit ninexnine_unit_3595(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B12G)
);

ninexnine_unit ninexnine_unit_3596(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C12G)
);

ninexnine_unit ninexnine_unit_3597(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D12G)
);

ninexnine_unit ninexnine_unit_3598(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E12G)
);

ninexnine_unit ninexnine_unit_3599(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F12G)
);

assign C112G=c1012G+c1112G+c1212G+c1312G+c1412G+c1512G+c1612G+c1712G+c1812G+c1912G+c1A12G+c1B12G+c1C12G+c1D12G+c1E12G+c1F12G;
assign A112G=(C112G>=0)?1:0;

assign P212G=A112G;

ninexnine_unit ninexnine_unit_3600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1020G)
);

ninexnine_unit ninexnine_unit_3601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1120G)
);

ninexnine_unit ninexnine_unit_3602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1220G)
);

ninexnine_unit ninexnine_unit_3603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1320G)
);

ninexnine_unit ninexnine_unit_3604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1420G)
);

ninexnine_unit ninexnine_unit_3605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1520G)
);

ninexnine_unit ninexnine_unit_3606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1620G)
);

ninexnine_unit ninexnine_unit_3607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1720G)
);

ninexnine_unit ninexnine_unit_3608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1820G)
);

ninexnine_unit ninexnine_unit_3609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1920G)
);

ninexnine_unit ninexnine_unit_3610(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A20G)
);

ninexnine_unit ninexnine_unit_3611(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B20G)
);

ninexnine_unit ninexnine_unit_3612(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C20G)
);

ninexnine_unit ninexnine_unit_3613(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D20G)
);

ninexnine_unit ninexnine_unit_3614(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E20G)
);

ninexnine_unit ninexnine_unit_3615(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F20G)
);

assign C120G=c1020G+c1120G+c1220G+c1320G+c1420G+c1520G+c1620G+c1720G+c1820G+c1920G+c1A20G+c1B20G+c1C20G+c1D20G+c1E20G+c1F20G;
assign A120G=(C120G>=0)?1:0;

assign P220G=A120G;

ninexnine_unit ninexnine_unit_3616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1021G)
);

ninexnine_unit ninexnine_unit_3617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1121G)
);

ninexnine_unit ninexnine_unit_3618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1221G)
);

ninexnine_unit ninexnine_unit_3619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1321G)
);

ninexnine_unit ninexnine_unit_3620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1421G)
);

ninexnine_unit ninexnine_unit_3621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1521G)
);

ninexnine_unit ninexnine_unit_3622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1621G)
);

ninexnine_unit ninexnine_unit_3623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1721G)
);

ninexnine_unit ninexnine_unit_3624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1821G)
);

ninexnine_unit ninexnine_unit_3625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1921G)
);

ninexnine_unit ninexnine_unit_3626(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A21G)
);

ninexnine_unit ninexnine_unit_3627(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B21G)
);

ninexnine_unit ninexnine_unit_3628(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C21G)
);

ninexnine_unit ninexnine_unit_3629(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D21G)
);

ninexnine_unit ninexnine_unit_3630(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E21G)
);

ninexnine_unit ninexnine_unit_3631(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F21G)
);

assign C121G=c1021G+c1121G+c1221G+c1321G+c1421G+c1521G+c1621G+c1721G+c1821G+c1921G+c1A21G+c1B21G+c1C21G+c1D21G+c1E21G+c1F21G;
assign A121G=(C121G>=0)?1:0;

assign P221G=A121G;

ninexnine_unit ninexnine_unit_3632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1G000),
				.b1(W1G010),
				.b2(W1G020),
				.b3(W1G100),
				.b4(W1G110),
				.b5(W1G120),
				.b6(W1G200),
				.b7(W1G210),
				.b8(W1G220),
				.c(c1022G)
);

ninexnine_unit ninexnine_unit_3633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1G001),
				.b1(W1G011),
				.b2(W1G021),
				.b3(W1G101),
				.b4(W1G111),
				.b5(W1G121),
				.b6(W1G201),
				.b7(W1G211),
				.b8(W1G221),
				.c(c1122G)
);

ninexnine_unit ninexnine_unit_3634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1G002),
				.b1(W1G012),
				.b2(W1G022),
				.b3(W1G102),
				.b4(W1G112),
				.b5(W1G122),
				.b6(W1G202),
				.b7(W1G212),
				.b8(W1G222),
				.c(c1222G)
);

ninexnine_unit ninexnine_unit_3635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1G003),
				.b1(W1G013),
				.b2(W1G023),
				.b3(W1G103),
				.b4(W1G113),
				.b5(W1G123),
				.b6(W1G203),
				.b7(W1G213),
				.b8(W1G223),
				.c(c1322G)
);

ninexnine_unit ninexnine_unit_3636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1G004),
				.b1(W1G014),
				.b2(W1G024),
				.b3(W1G104),
				.b4(W1G114),
				.b5(W1G124),
				.b6(W1G204),
				.b7(W1G214),
				.b8(W1G224),
				.c(c1422G)
);

ninexnine_unit ninexnine_unit_3637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1G005),
				.b1(W1G015),
				.b2(W1G025),
				.b3(W1G105),
				.b4(W1G115),
				.b5(W1G125),
				.b6(W1G205),
				.b7(W1G215),
				.b8(W1G225),
				.c(c1522G)
);

ninexnine_unit ninexnine_unit_3638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1G006),
				.b1(W1G016),
				.b2(W1G026),
				.b3(W1G106),
				.b4(W1G116),
				.b5(W1G126),
				.b6(W1G206),
				.b7(W1G216),
				.b8(W1G226),
				.c(c1622G)
);

ninexnine_unit ninexnine_unit_3639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1G007),
				.b1(W1G017),
				.b2(W1G027),
				.b3(W1G107),
				.b4(W1G117),
				.b5(W1G127),
				.b6(W1G207),
				.b7(W1G217),
				.b8(W1G227),
				.c(c1722G)
);

ninexnine_unit ninexnine_unit_3640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1G008),
				.b1(W1G018),
				.b2(W1G028),
				.b3(W1G108),
				.b4(W1G118),
				.b5(W1G128),
				.b6(W1G208),
				.b7(W1G218),
				.b8(W1G228),
				.c(c1822G)
);

ninexnine_unit ninexnine_unit_3641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1G009),
				.b1(W1G019),
				.b2(W1G029),
				.b3(W1G109),
				.b4(W1G119),
				.b5(W1G129),
				.b6(W1G209),
				.b7(W1G219),
				.b8(W1G229),
				.c(c1922G)
);

ninexnine_unit ninexnine_unit_3642(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1G00A),
				.b1(W1G01A),
				.b2(W1G02A),
				.b3(W1G10A),
				.b4(W1G11A),
				.b5(W1G12A),
				.b6(W1G20A),
				.b7(W1G21A),
				.b8(W1G22A),
				.c(c1A22G)
);

ninexnine_unit ninexnine_unit_3643(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1G00B),
				.b1(W1G01B),
				.b2(W1G02B),
				.b3(W1G10B),
				.b4(W1G11B),
				.b5(W1G12B),
				.b6(W1G20B),
				.b7(W1G21B),
				.b8(W1G22B),
				.c(c1B22G)
);

ninexnine_unit ninexnine_unit_3644(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1G00C),
				.b1(W1G01C),
				.b2(W1G02C),
				.b3(W1G10C),
				.b4(W1G11C),
				.b5(W1G12C),
				.b6(W1G20C),
				.b7(W1G21C),
				.b8(W1G22C),
				.c(c1C22G)
);

ninexnine_unit ninexnine_unit_3645(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1G00D),
				.b1(W1G01D),
				.b2(W1G02D),
				.b3(W1G10D),
				.b4(W1G11D),
				.b5(W1G12D),
				.b6(W1G20D),
				.b7(W1G21D),
				.b8(W1G22D),
				.c(c1D22G)
);

ninexnine_unit ninexnine_unit_3646(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1G00E),
				.b1(W1G01E),
				.b2(W1G02E),
				.b3(W1G10E),
				.b4(W1G11E),
				.b5(W1G12E),
				.b6(W1G20E),
				.b7(W1G21E),
				.b8(W1G22E),
				.c(c1E22G)
);

ninexnine_unit ninexnine_unit_3647(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1G00F),
				.b1(W1G01F),
				.b2(W1G02F),
				.b3(W1G10F),
				.b4(W1G11F),
				.b5(W1G12F),
				.b6(W1G20F),
				.b7(W1G21F),
				.b8(W1G22F),
				.c(c1F22G)
);

assign C122G=c1022G+c1122G+c1222G+c1322G+c1422G+c1522G+c1622G+c1722G+c1822G+c1922G+c1A22G+c1B22G+c1C22G+c1D22G+c1E22G+c1F22G;
assign A122G=(C122G>=0)?1:0;

assign P222G=A122G;

ninexnine_unit ninexnine_unit_3648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1000H)
);

ninexnine_unit ninexnine_unit_3649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1100H)
);

ninexnine_unit ninexnine_unit_3650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1200H)
);

ninexnine_unit ninexnine_unit_3651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1300H)
);

ninexnine_unit ninexnine_unit_3652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1400H)
);

ninexnine_unit ninexnine_unit_3653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1500H)
);

ninexnine_unit ninexnine_unit_3654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1600H)
);

ninexnine_unit ninexnine_unit_3655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1700H)
);

ninexnine_unit ninexnine_unit_3656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1800H)
);

ninexnine_unit ninexnine_unit_3657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1900H)
);

ninexnine_unit ninexnine_unit_3658(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A00H)
);

ninexnine_unit ninexnine_unit_3659(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B00H)
);

ninexnine_unit ninexnine_unit_3660(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C00H)
);

ninexnine_unit ninexnine_unit_3661(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D00H)
);

ninexnine_unit ninexnine_unit_3662(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E00H)
);

ninexnine_unit ninexnine_unit_3663(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F00H)
);

assign C100H=c1000H+c1100H+c1200H+c1300H+c1400H+c1500H+c1600H+c1700H+c1800H+c1900H+c1A00H+c1B00H+c1C00H+c1D00H+c1E00H+c1F00H;
assign A100H=(C100H>=0)?1:0;

assign P200H=A100H;

ninexnine_unit ninexnine_unit_3664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1001H)
);

ninexnine_unit ninexnine_unit_3665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1101H)
);

ninexnine_unit ninexnine_unit_3666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1201H)
);

ninexnine_unit ninexnine_unit_3667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1301H)
);

ninexnine_unit ninexnine_unit_3668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1401H)
);

ninexnine_unit ninexnine_unit_3669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1501H)
);

ninexnine_unit ninexnine_unit_3670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1601H)
);

ninexnine_unit ninexnine_unit_3671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1701H)
);

ninexnine_unit ninexnine_unit_3672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1801H)
);

ninexnine_unit ninexnine_unit_3673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1901H)
);

ninexnine_unit ninexnine_unit_3674(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A01H)
);

ninexnine_unit ninexnine_unit_3675(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B01H)
);

ninexnine_unit ninexnine_unit_3676(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C01H)
);

ninexnine_unit ninexnine_unit_3677(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D01H)
);

ninexnine_unit ninexnine_unit_3678(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E01H)
);

ninexnine_unit ninexnine_unit_3679(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F01H)
);

assign C101H=c1001H+c1101H+c1201H+c1301H+c1401H+c1501H+c1601H+c1701H+c1801H+c1901H+c1A01H+c1B01H+c1C01H+c1D01H+c1E01H+c1F01H;
assign A101H=(C101H>=0)?1:0;

assign P201H=A101H;

ninexnine_unit ninexnine_unit_3680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1002H)
);

ninexnine_unit ninexnine_unit_3681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1102H)
);

ninexnine_unit ninexnine_unit_3682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1202H)
);

ninexnine_unit ninexnine_unit_3683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1302H)
);

ninexnine_unit ninexnine_unit_3684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1402H)
);

ninexnine_unit ninexnine_unit_3685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1502H)
);

ninexnine_unit ninexnine_unit_3686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1602H)
);

ninexnine_unit ninexnine_unit_3687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1702H)
);

ninexnine_unit ninexnine_unit_3688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1802H)
);

ninexnine_unit ninexnine_unit_3689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1902H)
);

ninexnine_unit ninexnine_unit_3690(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A02H)
);

ninexnine_unit ninexnine_unit_3691(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B02H)
);

ninexnine_unit ninexnine_unit_3692(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C02H)
);

ninexnine_unit ninexnine_unit_3693(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D02H)
);

ninexnine_unit ninexnine_unit_3694(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E02H)
);

ninexnine_unit ninexnine_unit_3695(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F02H)
);

assign C102H=c1002H+c1102H+c1202H+c1302H+c1402H+c1502H+c1602H+c1702H+c1802H+c1902H+c1A02H+c1B02H+c1C02H+c1D02H+c1E02H+c1F02H;
assign A102H=(C102H>=0)?1:0;

assign P202H=A102H;

ninexnine_unit ninexnine_unit_3696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1010H)
);

ninexnine_unit ninexnine_unit_3697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1110H)
);

ninexnine_unit ninexnine_unit_3698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1210H)
);

ninexnine_unit ninexnine_unit_3699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1310H)
);

ninexnine_unit ninexnine_unit_3700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1410H)
);

ninexnine_unit ninexnine_unit_3701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1510H)
);

ninexnine_unit ninexnine_unit_3702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1610H)
);

ninexnine_unit ninexnine_unit_3703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1710H)
);

ninexnine_unit ninexnine_unit_3704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1810H)
);

ninexnine_unit ninexnine_unit_3705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1910H)
);

ninexnine_unit ninexnine_unit_3706(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A10H)
);

ninexnine_unit ninexnine_unit_3707(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B10H)
);

ninexnine_unit ninexnine_unit_3708(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C10H)
);

ninexnine_unit ninexnine_unit_3709(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D10H)
);

ninexnine_unit ninexnine_unit_3710(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E10H)
);

ninexnine_unit ninexnine_unit_3711(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F10H)
);

assign C110H=c1010H+c1110H+c1210H+c1310H+c1410H+c1510H+c1610H+c1710H+c1810H+c1910H+c1A10H+c1B10H+c1C10H+c1D10H+c1E10H+c1F10H;
assign A110H=(C110H>=0)?1:0;

assign P210H=A110H;

ninexnine_unit ninexnine_unit_3712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1011H)
);

ninexnine_unit ninexnine_unit_3713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1111H)
);

ninexnine_unit ninexnine_unit_3714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1211H)
);

ninexnine_unit ninexnine_unit_3715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1311H)
);

ninexnine_unit ninexnine_unit_3716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1411H)
);

ninexnine_unit ninexnine_unit_3717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1511H)
);

ninexnine_unit ninexnine_unit_3718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1611H)
);

ninexnine_unit ninexnine_unit_3719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1711H)
);

ninexnine_unit ninexnine_unit_3720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1811H)
);

ninexnine_unit ninexnine_unit_3721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1911H)
);

ninexnine_unit ninexnine_unit_3722(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A11H)
);

ninexnine_unit ninexnine_unit_3723(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B11H)
);

ninexnine_unit ninexnine_unit_3724(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C11H)
);

ninexnine_unit ninexnine_unit_3725(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D11H)
);

ninexnine_unit ninexnine_unit_3726(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E11H)
);

ninexnine_unit ninexnine_unit_3727(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F11H)
);

assign C111H=c1011H+c1111H+c1211H+c1311H+c1411H+c1511H+c1611H+c1711H+c1811H+c1911H+c1A11H+c1B11H+c1C11H+c1D11H+c1E11H+c1F11H;
assign A111H=(C111H>=0)?1:0;

assign P211H=A111H;

ninexnine_unit ninexnine_unit_3728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1012H)
);

ninexnine_unit ninexnine_unit_3729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1112H)
);

ninexnine_unit ninexnine_unit_3730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1212H)
);

ninexnine_unit ninexnine_unit_3731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1312H)
);

ninexnine_unit ninexnine_unit_3732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1412H)
);

ninexnine_unit ninexnine_unit_3733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1512H)
);

ninexnine_unit ninexnine_unit_3734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1612H)
);

ninexnine_unit ninexnine_unit_3735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1712H)
);

ninexnine_unit ninexnine_unit_3736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1812H)
);

ninexnine_unit ninexnine_unit_3737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1912H)
);

ninexnine_unit ninexnine_unit_3738(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A12H)
);

ninexnine_unit ninexnine_unit_3739(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B12H)
);

ninexnine_unit ninexnine_unit_3740(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C12H)
);

ninexnine_unit ninexnine_unit_3741(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D12H)
);

ninexnine_unit ninexnine_unit_3742(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E12H)
);

ninexnine_unit ninexnine_unit_3743(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F12H)
);

assign C112H=c1012H+c1112H+c1212H+c1312H+c1412H+c1512H+c1612H+c1712H+c1812H+c1912H+c1A12H+c1B12H+c1C12H+c1D12H+c1E12H+c1F12H;
assign A112H=(C112H>=0)?1:0;

assign P212H=A112H;

ninexnine_unit ninexnine_unit_3744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1020H)
);

ninexnine_unit ninexnine_unit_3745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1120H)
);

ninexnine_unit ninexnine_unit_3746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1220H)
);

ninexnine_unit ninexnine_unit_3747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1320H)
);

ninexnine_unit ninexnine_unit_3748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1420H)
);

ninexnine_unit ninexnine_unit_3749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1520H)
);

ninexnine_unit ninexnine_unit_3750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1620H)
);

ninexnine_unit ninexnine_unit_3751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1720H)
);

ninexnine_unit ninexnine_unit_3752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1820H)
);

ninexnine_unit ninexnine_unit_3753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1920H)
);

ninexnine_unit ninexnine_unit_3754(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A20H)
);

ninexnine_unit ninexnine_unit_3755(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B20H)
);

ninexnine_unit ninexnine_unit_3756(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C20H)
);

ninexnine_unit ninexnine_unit_3757(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D20H)
);

ninexnine_unit ninexnine_unit_3758(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E20H)
);

ninexnine_unit ninexnine_unit_3759(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F20H)
);

assign C120H=c1020H+c1120H+c1220H+c1320H+c1420H+c1520H+c1620H+c1720H+c1820H+c1920H+c1A20H+c1B20H+c1C20H+c1D20H+c1E20H+c1F20H;
assign A120H=(C120H>=0)?1:0;

assign P220H=A120H;

ninexnine_unit ninexnine_unit_3760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1021H)
);

ninexnine_unit ninexnine_unit_3761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1121H)
);

ninexnine_unit ninexnine_unit_3762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1221H)
);

ninexnine_unit ninexnine_unit_3763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1321H)
);

ninexnine_unit ninexnine_unit_3764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1421H)
);

ninexnine_unit ninexnine_unit_3765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1521H)
);

ninexnine_unit ninexnine_unit_3766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1621H)
);

ninexnine_unit ninexnine_unit_3767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1721H)
);

ninexnine_unit ninexnine_unit_3768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1821H)
);

ninexnine_unit ninexnine_unit_3769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1921H)
);

ninexnine_unit ninexnine_unit_3770(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A21H)
);

ninexnine_unit ninexnine_unit_3771(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B21H)
);

ninexnine_unit ninexnine_unit_3772(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C21H)
);

ninexnine_unit ninexnine_unit_3773(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D21H)
);

ninexnine_unit ninexnine_unit_3774(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E21H)
);

ninexnine_unit ninexnine_unit_3775(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F21H)
);

assign C121H=c1021H+c1121H+c1221H+c1321H+c1421H+c1521H+c1621H+c1721H+c1821H+c1921H+c1A21H+c1B21H+c1C21H+c1D21H+c1E21H+c1F21H;
assign A121H=(C121H>=0)?1:0;

assign P221H=A121H;

ninexnine_unit ninexnine_unit_3776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1H000),
				.b1(W1H010),
				.b2(W1H020),
				.b3(W1H100),
				.b4(W1H110),
				.b5(W1H120),
				.b6(W1H200),
				.b7(W1H210),
				.b8(W1H220),
				.c(c1022H)
);

ninexnine_unit ninexnine_unit_3777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1H001),
				.b1(W1H011),
				.b2(W1H021),
				.b3(W1H101),
				.b4(W1H111),
				.b5(W1H121),
				.b6(W1H201),
				.b7(W1H211),
				.b8(W1H221),
				.c(c1122H)
);

ninexnine_unit ninexnine_unit_3778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1H002),
				.b1(W1H012),
				.b2(W1H022),
				.b3(W1H102),
				.b4(W1H112),
				.b5(W1H122),
				.b6(W1H202),
				.b7(W1H212),
				.b8(W1H222),
				.c(c1222H)
);

ninexnine_unit ninexnine_unit_3779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1H003),
				.b1(W1H013),
				.b2(W1H023),
				.b3(W1H103),
				.b4(W1H113),
				.b5(W1H123),
				.b6(W1H203),
				.b7(W1H213),
				.b8(W1H223),
				.c(c1322H)
);

ninexnine_unit ninexnine_unit_3780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1H004),
				.b1(W1H014),
				.b2(W1H024),
				.b3(W1H104),
				.b4(W1H114),
				.b5(W1H124),
				.b6(W1H204),
				.b7(W1H214),
				.b8(W1H224),
				.c(c1422H)
);

ninexnine_unit ninexnine_unit_3781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1H005),
				.b1(W1H015),
				.b2(W1H025),
				.b3(W1H105),
				.b4(W1H115),
				.b5(W1H125),
				.b6(W1H205),
				.b7(W1H215),
				.b8(W1H225),
				.c(c1522H)
);

ninexnine_unit ninexnine_unit_3782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1H006),
				.b1(W1H016),
				.b2(W1H026),
				.b3(W1H106),
				.b4(W1H116),
				.b5(W1H126),
				.b6(W1H206),
				.b7(W1H216),
				.b8(W1H226),
				.c(c1622H)
);

ninexnine_unit ninexnine_unit_3783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1H007),
				.b1(W1H017),
				.b2(W1H027),
				.b3(W1H107),
				.b4(W1H117),
				.b5(W1H127),
				.b6(W1H207),
				.b7(W1H217),
				.b8(W1H227),
				.c(c1722H)
);

ninexnine_unit ninexnine_unit_3784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1H008),
				.b1(W1H018),
				.b2(W1H028),
				.b3(W1H108),
				.b4(W1H118),
				.b5(W1H128),
				.b6(W1H208),
				.b7(W1H218),
				.b8(W1H228),
				.c(c1822H)
);

ninexnine_unit ninexnine_unit_3785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1H009),
				.b1(W1H019),
				.b2(W1H029),
				.b3(W1H109),
				.b4(W1H119),
				.b5(W1H129),
				.b6(W1H209),
				.b7(W1H219),
				.b8(W1H229),
				.c(c1922H)
);

ninexnine_unit ninexnine_unit_3786(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1H00A),
				.b1(W1H01A),
				.b2(W1H02A),
				.b3(W1H10A),
				.b4(W1H11A),
				.b5(W1H12A),
				.b6(W1H20A),
				.b7(W1H21A),
				.b8(W1H22A),
				.c(c1A22H)
);

ninexnine_unit ninexnine_unit_3787(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1H00B),
				.b1(W1H01B),
				.b2(W1H02B),
				.b3(W1H10B),
				.b4(W1H11B),
				.b5(W1H12B),
				.b6(W1H20B),
				.b7(W1H21B),
				.b8(W1H22B),
				.c(c1B22H)
);

ninexnine_unit ninexnine_unit_3788(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1H00C),
				.b1(W1H01C),
				.b2(W1H02C),
				.b3(W1H10C),
				.b4(W1H11C),
				.b5(W1H12C),
				.b6(W1H20C),
				.b7(W1H21C),
				.b8(W1H22C),
				.c(c1C22H)
);

ninexnine_unit ninexnine_unit_3789(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1H00D),
				.b1(W1H01D),
				.b2(W1H02D),
				.b3(W1H10D),
				.b4(W1H11D),
				.b5(W1H12D),
				.b6(W1H20D),
				.b7(W1H21D),
				.b8(W1H22D),
				.c(c1D22H)
);

ninexnine_unit ninexnine_unit_3790(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1H00E),
				.b1(W1H01E),
				.b2(W1H02E),
				.b3(W1H10E),
				.b4(W1H11E),
				.b5(W1H12E),
				.b6(W1H20E),
				.b7(W1H21E),
				.b8(W1H22E),
				.c(c1E22H)
);

ninexnine_unit ninexnine_unit_3791(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1H00F),
				.b1(W1H01F),
				.b2(W1H02F),
				.b3(W1H10F),
				.b4(W1H11F),
				.b5(W1H12F),
				.b6(W1H20F),
				.b7(W1H21F),
				.b8(W1H22F),
				.c(c1F22H)
);

assign C122H=c1022H+c1122H+c1222H+c1322H+c1422H+c1522H+c1622H+c1722H+c1822H+c1922H+c1A22H+c1B22H+c1C22H+c1D22H+c1E22H+c1F22H;
assign A122H=(C122H>=0)?1:0;

assign P222H=A122H;

ninexnine_unit ninexnine_unit_3792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1000I)
);

ninexnine_unit ninexnine_unit_3793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1100I)
);

ninexnine_unit ninexnine_unit_3794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1200I)
);

ninexnine_unit ninexnine_unit_3795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1300I)
);

ninexnine_unit ninexnine_unit_3796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1400I)
);

ninexnine_unit ninexnine_unit_3797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1500I)
);

ninexnine_unit ninexnine_unit_3798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1600I)
);

ninexnine_unit ninexnine_unit_3799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1700I)
);

ninexnine_unit ninexnine_unit_3800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1800I)
);

ninexnine_unit ninexnine_unit_3801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1900I)
);

ninexnine_unit ninexnine_unit_3802(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A00I)
);

ninexnine_unit ninexnine_unit_3803(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B00I)
);

ninexnine_unit ninexnine_unit_3804(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C00I)
);

ninexnine_unit ninexnine_unit_3805(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D00I)
);

ninexnine_unit ninexnine_unit_3806(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E00I)
);

ninexnine_unit ninexnine_unit_3807(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F00I)
);

assign C100I=c1000I+c1100I+c1200I+c1300I+c1400I+c1500I+c1600I+c1700I+c1800I+c1900I+c1A00I+c1B00I+c1C00I+c1D00I+c1E00I+c1F00I;
assign A100I=(C100I>=0)?1:0;

assign P200I=A100I;

ninexnine_unit ninexnine_unit_3808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1001I)
);

ninexnine_unit ninexnine_unit_3809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1101I)
);

ninexnine_unit ninexnine_unit_3810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1201I)
);

ninexnine_unit ninexnine_unit_3811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1301I)
);

ninexnine_unit ninexnine_unit_3812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1401I)
);

ninexnine_unit ninexnine_unit_3813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1501I)
);

ninexnine_unit ninexnine_unit_3814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1601I)
);

ninexnine_unit ninexnine_unit_3815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1701I)
);

ninexnine_unit ninexnine_unit_3816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1801I)
);

ninexnine_unit ninexnine_unit_3817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1901I)
);

ninexnine_unit ninexnine_unit_3818(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A01I)
);

ninexnine_unit ninexnine_unit_3819(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B01I)
);

ninexnine_unit ninexnine_unit_3820(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C01I)
);

ninexnine_unit ninexnine_unit_3821(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D01I)
);

ninexnine_unit ninexnine_unit_3822(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E01I)
);

ninexnine_unit ninexnine_unit_3823(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F01I)
);

assign C101I=c1001I+c1101I+c1201I+c1301I+c1401I+c1501I+c1601I+c1701I+c1801I+c1901I+c1A01I+c1B01I+c1C01I+c1D01I+c1E01I+c1F01I;
assign A101I=(C101I>=0)?1:0;

assign P201I=A101I;

ninexnine_unit ninexnine_unit_3824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1002I)
);

ninexnine_unit ninexnine_unit_3825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1102I)
);

ninexnine_unit ninexnine_unit_3826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1202I)
);

ninexnine_unit ninexnine_unit_3827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1302I)
);

ninexnine_unit ninexnine_unit_3828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1402I)
);

ninexnine_unit ninexnine_unit_3829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1502I)
);

ninexnine_unit ninexnine_unit_3830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1602I)
);

ninexnine_unit ninexnine_unit_3831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1702I)
);

ninexnine_unit ninexnine_unit_3832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1802I)
);

ninexnine_unit ninexnine_unit_3833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1902I)
);

ninexnine_unit ninexnine_unit_3834(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A02I)
);

ninexnine_unit ninexnine_unit_3835(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B02I)
);

ninexnine_unit ninexnine_unit_3836(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C02I)
);

ninexnine_unit ninexnine_unit_3837(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D02I)
);

ninexnine_unit ninexnine_unit_3838(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E02I)
);

ninexnine_unit ninexnine_unit_3839(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F02I)
);

assign C102I=c1002I+c1102I+c1202I+c1302I+c1402I+c1502I+c1602I+c1702I+c1802I+c1902I+c1A02I+c1B02I+c1C02I+c1D02I+c1E02I+c1F02I;
assign A102I=(C102I>=0)?1:0;

assign P202I=A102I;

ninexnine_unit ninexnine_unit_3840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1010I)
);

ninexnine_unit ninexnine_unit_3841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1110I)
);

ninexnine_unit ninexnine_unit_3842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1210I)
);

ninexnine_unit ninexnine_unit_3843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1310I)
);

ninexnine_unit ninexnine_unit_3844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1410I)
);

ninexnine_unit ninexnine_unit_3845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1510I)
);

ninexnine_unit ninexnine_unit_3846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1610I)
);

ninexnine_unit ninexnine_unit_3847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1710I)
);

ninexnine_unit ninexnine_unit_3848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1810I)
);

ninexnine_unit ninexnine_unit_3849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1910I)
);

ninexnine_unit ninexnine_unit_3850(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A10I)
);

ninexnine_unit ninexnine_unit_3851(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B10I)
);

ninexnine_unit ninexnine_unit_3852(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C10I)
);

ninexnine_unit ninexnine_unit_3853(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D10I)
);

ninexnine_unit ninexnine_unit_3854(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E10I)
);

ninexnine_unit ninexnine_unit_3855(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F10I)
);

assign C110I=c1010I+c1110I+c1210I+c1310I+c1410I+c1510I+c1610I+c1710I+c1810I+c1910I+c1A10I+c1B10I+c1C10I+c1D10I+c1E10I+c1F10I;
assign A110I=(C110I>=0)?1:0;

assign P210I=A110I;

ninexnine_unit ninexnine_unit_3856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1011I)
);

ninexnine_unit ninexnine_unit_3857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1111I)
);

ninexnine_unit ninexnine_unit_3858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1211I)
);

ninexnine_unit ninexnine_unit_3859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1311I)
);

ninexnine_unit ninexnine_unit_3860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1411I)
);

ninexnine_unit ninexnine_unit_3861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1511I)
);

ninexnine_unit ninexnine_unit_3862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1611I)
);

ninexnine_unit ninexnine_unit_3863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1711I)
);

ninexnine_unit ninexnine_unit_3864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1811I)
);

ninexnine_unit ninexnine_unit_3865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1911I)
);

ninexnine_unit ninexnine_unit_3866(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A11I)
);

ninexnine_unit ninexnine_unit_3867(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B11I)
);

ninexnine_unit ninexnine_unit_3868(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C11I)
);

ninexnine_unit ninexnine_unit_3869(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D11I)
);

ninexnine_unit ninexnine_unit_3870(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E11I)
);

ninexnine_unit ninexnine_unit_3871(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F11I)
);

assign C111I=c1011I+c1111I+c1211I+c1311I+c1411I+c1511I+c1611I+c1711I+c1811I+c1911I+c1A11I+c1B11I+c1C11I+c1D11I+c1E11I+c1F11I;
assign A111I=(C111I>=0)?1:0;

assign P211I=A111I;

ninexnine_unit ninexnine_unit_3872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1012I)
);

ninexnine_unit ninexnine_unit_3873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1112I)
);

ninexnine_unit ninexnine_unit_3874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1212I)
);

ninexnine_unit ninexnine_unit_3875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1312I)
);

ninexnine_unit ninexnine_unit_3876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1412I)
);

ninexnine_unit ninexnine_unit_3877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1512I)
);

ninexnine_unit ninexnine_unit_3878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1612I)
);

ninexnine_unit ninexnine_unit_3879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1712I)
);

ninexnine_unit ninexnine_unit_3880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1812I)
);

ninexnine_unit ninexnine_unit_3881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1912I)
);

ninexnine_unit ninexnine_unit_3882(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A12I)
);

ninexnine_unit ninexnine_unit_3883(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B12I)
);

ninexnine_unit ninexnine_unit_3884(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C12I)
);

ninexnine_unit ninexnine_unit_3885(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D12I)
);

ninexnine_unit ninexnine_unit_3886(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E12I)
);

ninexnine_unit ninexnine_unit_3887(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F12I)
);

assign C112I=c1012I+c1112I+c1212I+c1312I+c1412I+c1512I+c1612I+c1712I+c1812I+c1912I+c1A12I+c1B12I+c1C12I+c1D12I+c1E12I+c1F12I;
assign A112I=(C112I>=0)?1:0;

assign P212I=A112I;

ninexnine_unit ninexnine_unit_3888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1020I)
);

ninexnine_unit ninexnine_unit_3889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1120I)
);

ninexnine_unit ninexnine_unit_3890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1220I)
);

ninexnine_unit ninexnine_unit_3891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1320I)
);

ninexnine_unit ninexnine_unit_3892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1420I)
);

ninexnine_unit ninexnine_unit_3893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1520I)
);

ninexnine_unit ninexnine_unit_3894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1620I)
);

ninexnine_unit ninexnine_unit_3895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1720I)
);

ninexnine_unit ninexnine_unit_3896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1820I)
);

ninexnine_unit ninexnine_unit_3897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1920I)
);

ninexnine_unit ninexnine_unit_3898(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A20I)
);

ninexnine_unit ninexnine_unit_3899(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B20I)
);

ninexnine_unit ninexnine_unit_3900(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C20I)
);

ninexnine_unit ninexnine_unit_3901(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D20I)
);

ninexnine_unit ninexnine_unit_3902(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E20I)
);

ninexnine_unit ninexnine_unit_3903(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F20I)
);

assign C120I=c1020I+c1120I+c1220I+c1320I+c1420I+c1520I+c1620I+c1720I+c1820I+c1920I+c1A20I+c1B20I+c1C20I+c1D20I+c1E20I+c1F20I;
assign A120I=(C120I>=0)?1:0;

assign P220I=A120I;

ninexnine_unit ninexnine_unit_3904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1021I)
);

ninexnine_unit ninexnine_unit_3905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1121I)
);

ninexnine_unit ninexnine_unit_3906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1221I)
);

ninexnine_unit ninexnine_unit_3907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1321I)
);

ninexnine_unit ninexnine_unit_3908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1421I)
);

ninexnine_unit ninexnine_unit_3909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1521I)
);

ninexnine_unit ninexnine_unit_3910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1621I)
);

ninexnine_unit ninexnine_unit_3911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1721I)
);

ninexnine_unit ninexnine_unit_3912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1821I)
);

ninexnine_unit ninexnine_unit_3913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1921I)
);

ninexnine_unit ninexnine_unit_3914(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A21I)
);

ninexnine_unit ninexnine_unit_3915(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B21I)
);

ninexnine_unit ninexnine_unit_3916(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C21I)
);

ninexnine_unit ninexnine_unit_3917(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D21I)
);

ninexnine_unit ninexnine_unit_3918(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E21I)
);

ninexnine_unit ninexnine_unit_3919(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F21I)
);

assign C121I=c1021I+c1121I+c1221I+c1321I+c1421I+c1521I+c1621I+c1721I+c1821I+c1921I+c1A21I+c1B21I+c1C21I+c1D21I+c1E21I+c1F21I;
assign A121I=(C121I>=0)?1:0;

assign P221I=A121I;

ninexnine_unit ninexnine_unit_3920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1I000),
				.b1(W1I010),
				.b2(W1I020),
				.b3(W1I100),
				.b4(W1I110),
				.b5(W1I120),
				.b6(W1I200),
				.b7(W1I210),
				.b8(W1I220),
				.c(c1022I)
);

ninexnine_unit ninexnine_unit_3921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1I001),
				.b1(W1I011),
				.b2(W1I021),
				.b3(W1I101),
				.b4(W1I111),
				.b5(W1I121),
				.b6(W1I201),
				.b7(W1I211),
				.b8(W1I221),
				.c(c1122I)
);

ninexnine_unit ninexnine_unit_3922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1I002),
				.b1(W1I012),
				.b2(W1I022),
				.b3(W1I102),
				.b4(W1I112),
				.b5(W1I122),
				.b6(W1I202),
				.b7(W1I212),
				.b8(W1I222),
				.c(c1222I)
);

ninexnine_unit ninexnine_unit_3923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1I003),
				.b1(W1I013),
				.b2(W1I023),
				.b3(W1I103),
				.b4(W1I113),
				.b5(W1I123),
				.b6(W1I203),
				.b7(W1I213),
				.b8(W1I223),
				.c(c1322I)
);

ninexnine_unit ninexnine_unit_3924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1I004),
				.b1(W1I014),
				.b2(W1I024),
				.b3(W1I104),
				.b4(W1I114),
				.b5(W1I124),
				.b6(W1I204),
				.b7(W1I214),
				.b8(W1I224),
				.c(c1422I)
);

ninexnine_unit ninexnine_unit_3925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1I005),
				.b1(W1I015),
				.b2(W1I025),
				.b3(W1I105),
				.b4(W1I115),
				.b5(W1I125),
				.b6(W1I205),
				.b7(W1I215),
				.b8(W1I225),
				.c(c1522I)
);

ninexnine_unit ninexnine_unit_3926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1I006),
				.b1(W1I016),
				.b2(W1I026),
				.b3(W1I106),
				.b4(W1I116),
				.b5(W1I126),
				.b6(W1I206),
				.b7(W1I216),
				.b8(W1I226),
				.c(c1622I)
);

ninexnine_unit ninexnine_unit_3927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1I007),
				.b1(W1I017),
				.b2(W1I027),
				.b3(W1I107),
				.b4(W1I117),
				.b5(W1I127),
				.b6(W1I207),
				.b7(W1I217),
				.b8(W1I227),
				.c(c1722I)
);

ninexnine_unit ninexnine_unit_3928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1I008),
				.b1(W1I018),
				.b2(W1I028),
				.b3(W1I108),
				.b4(W1I118),
				.b5(W1I128),
				.b6(W1I208),
				.b7(W1I218),
				.b8(W1I228),
				.c(c1822I)
);

ninexnine_unit ninexnine_unit_3929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1I009),
				.b1(W1I019),
				.b2(W1I029),
				.b3(W1I109),
				.b4(W1I119),
				.b5(W1I129),
				.b6(W1I209),
				.b7(W1I219),
				.b8(W1I229),
				.c(c1922I)
);

ninexnine_unit ninexnine_unit_3930(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1I00A),
				.b1(W1I01A),
				.b2(W1I02A),
				.b3(W1I10A),
				.b4(W1I11A),
				.b5(W1I12A),
				.b6(W1I20A),
				.b7(W1I21A),
				.b8(W1I22A),
				.c(c1A22I)
);

ninexnine_unit ninexnine_unit_3931(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1I00B),
				.b1(W1I01B),
				.b2(W1I02B),
				.b3(W1I10B),
				.b4(W1I11B),
				.b5(W1I12B),
				.b6(W1I20B),
				.b7(W1I21B),
				.b8(W1I22B),
				.c(c1B22I)
);

ninexnine_unit ninexnine_unit_3932(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1I00C),
				.b1(W1I01C),
				.b2(W1I02C),
				.b3(W1I10C),
				.b4(W1I11C),
				.b5(W1I12C),
				.b6(W1I20C),
				.b7(W1I21C),
				.b8(W1I22C),
				.c(c1C22I)
);

ninexnine_unit ninexnine_unit_3933(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1I00D),
				.b1(W1I01D),
				.b2(W1I02D),
				.b3(W1I10D),
				.b4(W1I11D),
				.b5(W1I12D),
				.b6(W1I20D),
				.b7(W1I21D),
				.b8(W1I22D),
				.c(c1D22I)
);

ninexnine_unit ninexnine_unit_3934(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1I00E),
				.b1(W1I01E),
				.b2(W1I02E),
				.b3(W1I10E),
				.b4(W1I11E),
				.b5(W1I12E),
				.b6(W1I20E),
				.b7(W1I21E),
				.b8(W1I22E),
				.c(c1E22I)
);

ninexnine_unit ninexnine_unit_3935(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1I00F),
				.b1(W1I01F),
				.b2(W1I02F),
				.b3(W1I10F),
				.b4(W1I11F),
				.b5(W1I12F),
				.b6(W1I20F),
				.b7(W1I21F),
				.b8(W1I22F),
				.c(c1F22I)
);

assign C122I=c1022I+c1122I+c1222I+c1322I+c1422I+c1522I+c1622I+c1722I+c1822I+c1922I+c1A22I+c1B22I+c1C22I+c1D22I+c1E22I+c1F22I;
assign A122I=(C122I>=0)?1:0;

assign P222I=A122I;

ninexnine_unit ninexnine_unit_3936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1000J)
);

ninexnine_unit ninexnine_unit_3937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1100J)
);

ninexnine_unit ninexnine_unit_3938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1200J)
);

ninexnine_unit ninexnine_unit_3939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1300J)
);

ninexnine_unit ninexnine_unit_3940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1400J)
);

ninexnine_unit ninexnine_unit_3941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1500J)
);

ninexnine_unit ninexnine_unit_3942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1600J)
);

ninexnine_unit ninexnine_unit_3943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1700J)
);

ninexnine_unit ninexnine_unit_3944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1800J)
);

ninexnine_unit ninexnine_unit_3945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1900J)
);

ninexnine_unit ninexnine_unit_3946(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A00J)
);

ninexnine_unit ninexnine_unit_3947(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B00J)
);

ninexnine_unit ninexnine_unit_3948(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C00J)
);

ninexnine_unit ninexnine_unit_3949(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D00J)
);

ninexnine_unit ninexnine_unit_3950(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E00J)
);

ninexnine_unit ninexnine_unit_3951(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F00J)
);

assign C100J=c1000J+c1100J+c1200J+c1300J+c1400J+c1500J+c1600J+c1700J+c1800J+c1900J+c1A00J+c1B00J+c1C00J+c1D00J+c1E00J+c1F00J;
assign A100J=(C100J>=0)?1:0;

assign P200J=A100J;

ninexnine_unit ninexnine_unit_3952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1001J)
);

ninexnine_unit ninexnine_unit_3953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1101J)
);

ninexnine_unit ninexnine_unit_3954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1201J)
);

ninexnine_unit ninexnine_unit_3955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1301J)
);

ninexnine_unit ninexnine_unit_3956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1401J)
);

ninexnine_unit ninexnine_unit_3957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1501J)
);

ninexnine_unit ninexnine_unit_3958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1601J)
);

ninexnine_unit ninexnine_unit_3959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1701J)
);

ninexnine_unit ninexnine_unit_3960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1801J)
);

ninexnine_unit ninexnine_unit_3961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1901J)
);

ninexnine_unit ninexnine_unit_3962(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A01J)
);

ninexnine_unit ninexnine_unit_3963(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B01J)
);

ninexnine_unit ninexnine_unit_3964(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C01J)
);

ninexnine_unit ninexnine_unit_3965(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D01J)
);

ninexnine_unit ninexnine_unit_3966(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E01J)
);

ninexnine_unit ninexnine_unit_3967(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F01J)
);

assign C101J=c1001J+c1101J+c1201J+c1301J+c1401J+c1501J+c1601J+c1701J+c1801J+c1901J+c1A01J+c1B01J+c1C01J+c1D01J+c1E01J+c1F01J;
assign A101J=(C101J>=0)?1:0;

assign P201J=A101J;

ninexnine_unit ninexnine_unit_3968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1002J)
);

ninexnine_unit ninexnine_unit_3969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1102J)
);

ninexnine_unit ninexnine_unit_3970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1202J)
);

ninexnine_unit ninexnine_unit_3971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1302J)
);

ninexnine_unit ninexnine_unit_3972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1402J)
);

ninexnine_unit ninexnine_unit_3973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1502J)
);

ninexnine_unit ninexnine_unit_3974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1602J)
);

ninexnine_unit ninexnine_unit_3975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1702J)
);

ninexnine_unit ninexnine_unit_3976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1802J)
);

ninexnine_unit ninexnine_unit_3977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1902J)
);

ninexnine_unit ninexnine_unit_3978(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A02J)
);

ninexnine_unit ninexnine_unit_3979(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B02J)
);

ninexnine_unit ninexnine_unit_3980(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C02J)
);

ninexnine_unit ninexnine_unit_3981(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D02J)
);

ninexnine_unit ninexnine_unit_3982(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E02J)
);

ninexnine_unit ninexnine_unit_3983(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F02J)
);

assign C102J=c1002J+c1102J+c1202J+c1302J+c1402J+c1502J+c1602J+c1702J+c1802J+c1902J+c1A02J+c1B02J+c1C02J+c1D02J+c1E02J+c1F02J;
assign A102J=(C102J>=0)?1:0;

assign P202J=A102J;

ninexnine_unit ninexnine_unit_3984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1010J)
);

ninexnine_unit ninexnine_unit_3985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1110J)
);

ninexnine_unit ninexnine_unit_3986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1210J)
);

ninexnine_unit ninexnine_unit_3987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1310J)
);

ninexnine_unit ninexnine_unit_3988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1410J)
);

ninexnine_unit ninexnine_unit_3989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1510J)
);

ninexnine_unit ninexnine_unit_3990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1610J)
);

ninexnine_unit ninexnine_unit_3991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1710J)
);

ninexnine_unit ninexnine_unit_3992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1810J)
);

ninexnine_unit ninexnine_unit_3993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1910J)
);

ninexnine_unit ninexnine_unit_3994(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A10J)
);

ninexnine_unit ninexnine_unit_3995(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B10J)
);

ninexnine_unit ninexnine_unit_3996(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C10J)
);

ninexnine_unit ninexnine_unit_3997(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D10J)
);

ninexnine_unit ninexnine_unit_3998(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E10J)
);

ninexnine_unit ninexnine_unit_3999(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F10J)
);

assign C110J=c1010J+c1110J+c1210J+c1310J+c1410J+c1510J+c1610J+c1710J+c1810J+c1910J+c1A10J+c1B10J+c1C10J+c1D10J+c1E10J+c1F10J;
assign A110J=(C110J>=0)?1:0;

assign P210J=A110J;

ninexnine_unit ninexnine_unit_4000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1011J)
);

ninexnine_unit ninexnine_unit_4001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1111J)
);

ninexnine_unit ninexnine_unit_4002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1211J)
);

ninexnine_unit ninexnine_unit_4003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1311J)
);

ninexnine_unit ninexnine_unit_4004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1411J)
);

ninexnine_unit ninexnine_unit_4005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1511J)
);

ninexnine_unit ninexnine_unit_4006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1611J)
);

ninexnine_unit ninexnine_unit_4007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1711J)
);

ninexnine_unit ninexnine_unit_4008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1811J)
);

ninexnine_unit ninexnine_unit_4009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1911J)
);

ninexnine_unit ninexnine_unit_4010(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A11J)
);

ninexnine_unit ninexnine_unit_4011(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B11J)
);

ninexnine_unit ninexnine_unit_4012(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C11J)
);

ninexnine_unit ninexnine_unit_4013(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D11J)
);

ninexnine_unit ninexnine_unit_4014(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E11J)
);

ninexnine_unit ninexnine_unit_4015(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F11J)
);

assign C111J=c1011J+c1111J+c1211J+c1311J+c1411J+c1511J+c1611J+c1711J+c1811J+c1911J+c1A11J+c1B11J+c1C11J+c1D11J+c1E11J+c1F11J;
assign A111J=(C111J>=0)?1:0;

assign P211J=A111J;

ninexnine_unit ninexnine_unit_4016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1012J)
);

ninexnine_unit ninexnine_unit_4017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1112J)
);

ninexnine_unit ninexnine_unit_4018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1212J)
);

ninexnine_unit ninexnine_unit_4019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1312J)
);

ninexnine_unit ninexnine_unit_4020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1412J)
);

ninexnine_unit ninexnine_unit_4021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1512J)
);

ninexnine_unit ninexnine_unit_4022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1612J)
);

ninexnine_unit ninexnine_unit_4023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1712J)
);

ninexnine_unit ninexnine_unit_4024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1812J)
);

ninexnine_unit ninexnine_unit_4025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1912J)
);

ninexnine_unit ninexnine_unit_4026(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A12J)
);

ninexnine_unit ninexnine_unit_4027(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B12J)
);

ninexnine_unit ninexnine_unit_4028(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C12J)
);

ninexnine_unit ninexnine_unit_4029(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D12J)
);

ninexnine_unit ninexnine_unit_4030(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E12J)
);

ninexnine_unit ninexnine_unit_4031(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F12J)
);

assign C112J=c1012J+c1112J+c1212J+c1312J+c1412J+c1512J+c1612J+c1712J+c1812J+c1912J+c1A12J+c1B12J+c1C12J+c1D12J+c1E12J+c1F12J;
assign A112J=(C112J>=0)?1:0;

assign P212J=A112J;

ninexnine_unit ninexnine_unit_4032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1020J)
);

ninexnine_unit ninexnine_unit_4033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1120J)
);

ninexnine_unit ninexnine_unit_4034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1220J)
);

ninexnine_unit ninexnine_unit_4035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1320J)
);

ninexnine_unit ninexnine_unit_4036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1420J)
);

ninexnine_unit ninexnine_unit_4037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1520J)
);

ninexnine_unit ninexnine_unit_4038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1620J)
);

ninexnine_unit ninexnine_unit_4039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1720J)
);

ninexnine_unit ninexnine_unit_4040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1820J)
);

ninexnine_unit ninexnine_unit_4041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1920J)
);

ninexnine_unit ninexnine_unit_4042(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A20J)
);

ninexnine_unit ninexnine_unit_4043(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B20J)
);

ninexnine_unit ninexnine_unit_4044(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C20J)
);

ninexnine_unit ninexnine_unit_4045(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D20J)
);

ninexnine_unit ninexnine_unit_4046(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E20J)
);

ninexnine_unit ninexnine_unit_4047(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F20J)
);

assign C120J=c1020J+c1120J+c1220J+c1320J+c1420J+c1520J+c1620J+c1720J+c1820J+c1920J+c1A20J+c1B20J+c1C20J+c1D20J+c1E20J+c1F20J;
assign A120J=(C120J>=0)?1:0;

assign P220J=A120J;

ninexnine_unit ninexnine_unit_4048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1021J)
);

ninexnine_unit ninexnine_unit_4049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1121J)
);

ninexnine_unit ninexnine_unit_4050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1221J)
);

ninexnine_unit ninexnine_unit_4051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1321J)
);

ninexnine_unit ninexnine_unit_4052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1421J)
);

ninexnine_unit ninexnine_unit_4053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1521J)
);

ninexnine_unit ninexnine_unit_4054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1621J)
);

ninexnine_unit ninexnine_unit_4055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1721J)
);

ninexnine_unit ninexnine_unit_4056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1821J)
);

ninexnine_unit ninexnine_unit_4057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1921J)
);

ninexnine_unit ninexnine_unit_4058(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A21J)
);

ninexnine_unit ninexnine_unit_4059(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B21J)
);

ninexnine_unit ninexnine_unit_4060(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C21J)
);

ninexnine_unit ninexnine_unit_4061(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D21J)
);

ninexnine_unit ninexnine_unit_4062(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E21J)
);

ninexnine_unit ninexnine_unit_4063(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F21J)
);

assign C121J=c1021J+c1121J+c1221J+c1321J+c1421J+c1521J+c1621J+c1721J+c1821J+c1921J+c1A21J+c1B21J+c1C21J+c1D21J+c1E21J+c1F21J;
assign A121J=(C121J>=0)?1:0;

assign P221J=A121J;

ninexnine_unit ninexnine_unit_4064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1J000),
				.b1(W1J010),
				.b2(W1J020),
				.b3(W1J100),
				.b4(W1J110),
				.b5(W1J120),
				.b6(W1J200),
				.b7(W1J210),
				.b8(W1J220),
				.c(c1022J)
);

ninexnine_unit ninexnine_unit_4065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1J001),
				.b1(W1J011),
				.b2(W1J021),
				.b3(W1J101),
				.b4(W1J111),
				.b5(W1J121),
				.b6(W1J201),
				.b7(W1J211),
				.b8(W1J221),
				.c(c1122J)
);

ninexnine_unit ninexnine_unit_4066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1J002),
				.b1(W1J012),
				.b2(W1J022),
				.b3(W1J102),
				.b4(W1J112),
				.b5(W1J122),
				.b6(W1J202),
				.b7(W1J212),
				.b8(W1J222),
				.c(c1222J)
);

ninexnine_unit ninexnine_unit_4067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1J003),
				.b1(W1J013),
				.b2(W1J023),
				.b3(W1J103),
				.b4(W1J113),
				.b5(W1J123),
				.b6(W1J203),
				.b7(W1J213),
				.b8(W1J223),
				.c(c1322J)
);

ninexnine_unit ninexnine_unit_4068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1J004),
				.b1(W1J014),
				.b2(W1J024),
				.b3(W1J104),
				.b4(W1J114),
				.b5(W1J124),
				.b6(W1J204),
				.b7(W1J214),
				.b8(W1J224),
				.c(c1422J)
);

ninexnine_unit ninexnine_unit_4069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1J005),
				.b1(W1J015),
				.b2(W1J025),
				.b3(W1J105),
				.b4(W1J115),
				.b5(W1J125),
				.b6(W1J205),
				.b7(W1J215),
				.b8(W1J225),
				.c(c1522J)
);

ninexnine_unit ninexnine_unit_4070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1J006),
				.b1(W1J016),
				.b2(W1J026),
				.b3(W1J106),
				.b4(W1J116),
				.b5(W1J126),
				.b6(W1J206),
				.b7(W1J216),
				.b8(W1J226),
				.c(c1622J)
);

ninexnine_unit ninexnine_unit_4071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1J007),
				.b1(W1J017),
				.b2(W1J027),
				.b3(W1J107),
				.b4(W1J117),
				.b5(W1J127),
				.b6(W1J207),
				.b7(W1J217),
				.b8(W1J227),
				.c(c1722J)
);

ninexnine_unit ninexnine_unit_4072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1J008),
				.b1(W1J018),
				.b2(W1J028),
				.b3(W1J108),
				.b4(W1J118),
				.b5(W1J128),
				.b6(W1J208),
				.b7(W1J218),
				.b8(W1J228),
				.c(c1822J)
);

ninexnine_unit ninexnine_unit_4073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1J009),
				.b1(W1J019),
				.b2(W1J029),
				.b3(W1J109),
				.b4(W1J119),
				.b5(W1J129),
				.b6(W1J209),
				.b7(W1J219),
				.b8(W1J229),
				.c(c1922J)
);

ninexnine_unit ninexnine_unit_4074(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1J00A),
				.b1(W1J01A),
				.b2(W1J02A),
				.b3(W1J10A),
				.b4(W1J11A),
				.b5(W1J12A),
				.b6(W1J20A),
				.b7(W1J21A),
				.b8(W1J22A),
				.c(c1A22J)
);

ninexnine_unit ninexnine_unit_4075(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1J00B),
				.b1(W1J01B),
				.b2(W1J02B),
				.b3(W1J10B),
				.b4(W1J11B),
				.b5(W1J12B),
				.b6(W1J20B),
				.b7(W1J21B),
				.b8(W1J22B),
				.c(c1B22J)
);

ninexnine_unit ninexnine_unit_4076(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1J00C),
				.b1(W1J01C),
				.b2(W1J02C),
				.b3(W1J10C),
				.b4(W1J11C),
				.b5(W1J12C),
				.b6(W1J20C),
				.b7(W1J21C),
				.b8(W1J22C),
				.c(c1C22J)
);

ninexnine_unit ninexnine_unit_4077(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1J00D),
				.b1(W1J01D),
				.b2(W1J02D),
				.b3(W1J10D),
				.b4(W1J11D),
				.b5(W1J12D),
				.b6(W1J20D),
				.b7(W1J21D),
				.b8(W1J22D),
				.c(c1D22J)
);

ninexnine_unit ninexnine_unit_4078(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1J00E),
				.b1(W1J01E),
				.b2(W1J02E),
				.b3(W1J10E),
				.b4(W1J11E),
				.b5(W1J12E),
				.b6(W1J20E),
				.b7(W1J21E),
				.b8(W1J22E),
				.c(c1E22J)
);

ninexnine_unit ninexnine_unit_4079(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1J00F),
				.b1(W1J01F),
				.b2(W1J02F),
				.b3(W1J10F),
				.b4(W1J11F),
				.b5(W1J12F),
				.b6(W1J20F),
				.b7(W1J21F),
				.b8(W1J22F),
				.c(c1F22J)
);

assign C122J=c1022J+c1122J+c1222J+c1322J+c1422J+c1522J+c1622J+c1722J+c1822J+c1922J+c1A22J+c1B22J+c1C22J+c1D22J+c1E22J+c1F22J;
assign A122J=(C122J>=0)?1:0;

assign P222J=A122J;

ninexnine_unit ninexnine_unit_4080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1000K)
);

ninexnine_unit ninexnine_unit_4081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1100K)
);

ninexnine_unit ninexnine_unit_4082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1200K)
);

ninexnine_unit ninexnine_unit_4083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1300K)
);

ninexnine_unit ninexnine_unit_4084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1400K)
);

ninexnine_unit ninexnine_unit_4085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1500K)
);

ninexnine_unit ninexnine_unit_4086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1600K)
);

ninexnine_unit ninexnine_unit_4087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1700K)
);

ninexnine_unit ninexnine_unit_4088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1800K)
);

ninexnine_unit ninexnine_unit_4089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1900K)
);

ninexnine_unit ninexnine_unit_4090(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A00K)
);

ninexnine_unit ninexnine_unit_4091(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B00K)
);

ninexnine_unit ninexnine_unit_4092(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C00K)
);

ninexnine_unit ninexnine_unit_4093(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D00K)
);

ninexnine_unit ninexnine_unit_4094(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E00K)
);

ninexnine_unit ninexnine_unit_4095(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F00K)
);

assign C100K=c1000K+c1100K+c1200K+c1300K+c1400K+c1500K+c1600K+c1700K+c1800K+c1900K+c1A00K+c1B00K+c1C00K+c1D00K+c1E00K+c1F00K;
assign A100K=(C100K>=0)?1:0;

assign P200K=A100K;

ninexnine_unit ninexnine_unit_4096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1001K)
);

ninexnine_unit ninexnine_unit_4097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1101K)
);

ninexnine_unit ninexnine_unit_4098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1201K)
);

ninexnine_unit ninexnine_unit_4099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1301K)
);

ninexnine_unit ninexnine_unit_4100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1401K)
);

ninexnine_unit ninexnine_unit_4101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1501K)
);

ninexnine_unit ninexnine_unit_4102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1601K)
);

ninexnine_unit ninexnine_unit_4103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1701K)
);

ninexnine_unit ninexnine_unit_4104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1801K)
);

ninexnine_unit ninexnine_unit_4105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1901K)
);

ninexnine_unit ninexnine_unit_4106(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A01K)
);

ninexnine_unit ninexnine_unit_4107(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B01K)
);

ninexnine_unit ninexnine_unit_4108(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C01K)
);

ninexnine_unit ninexnine_unit_4109(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D01K)
);

ninexnine_unit ninexnine_unit_4110(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E01K)
);

ninexnine_unit ninexnine_unit_4111(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F01K)
);

assign C101K=c1001K+c1101K+c1201K+c1301K+c1401K+c1501K+c1601K+c1701K+c1801K+c1901K+c1A01K+c1B01K+c1C01K+c1D01K+c1E01K+c1F01K;
assign A101K=(C101K>=0)?1:0;

assign P201K=A101K;

ninexnine_unit ninexnine_unit_4112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1002K)
);

ninexnine_unit ninexnine_unit_4113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1102K)
);

ninexnine_unit ninexnine_unit_4114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1202K)
);

ninexnine_unit ninexnine_unit_4115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1302K)
);

ninexnine_unit ninexnine_unit_4116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1402K)
);

ninexnine_unit ninexnine_unit_4117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1502K)
);

ninexnine_unit ninexnine_unit_4118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1602K)
);

ninexnine_unit ninexnine_unit_4119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1702K)
);

ninexnine_unit ninexnine_unit_4120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1802K)
);

ninexnine_unit ninexnine_unit_4121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1902K)
);

ninexnine_unit ninexnine_unit_4122(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A02K)
);

ninexnine_unit ninexnine_unit_4123(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B02K)
);

ninexnine_unit ninexnine_unit_4124(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C02K)
);

ninexnine_unit ninexnine_unit_4125(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D02K)
);

ninexnine_unit ninexnine_unit_4126(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E02K)
);

ninexnine_unit ninexnine_unit_4127(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F02K)
);

assign C102K=c1002K+c1102K+c1202K+c1302K+c1402K+c1502K+c1602K+c1702K+c1802K+c1902K+c1A02K+c1B02K+c1C02K+c1D02K+c1E02K+c1F02K;
assign A102K=(C102K>=0)?1:0;

assign P202K=A102K;

ninexnine_unit ninexnine_unit_4128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1010K)
);

ninexnine_unit ninexnine_unit_4129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1110K)
);

ninexnine_unit ninexnine_unit_4130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1210K)
);

ninexnine_unit ninexnine_unit_4131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1310K)
);

ninexnine_unit ninexnine_unit_4132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1410K)
);

ninexnine_unit ninexnine_unit_4133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1510K)
);

ninexnine_unit ninexnine_unit_4134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1610K)
);

ninexnine_unit ninexnine_unit_4135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1710K)
);

ninexnine_unit ninexnine_unit_4136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1810K)
);

ninexnine_unit ninexnine_unit_4137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1910K)
);

ninexnine_unit ninexnine_unit_4138(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A10K)
);

ninexnine_unit ninexnine_unit_4139(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B10K)
);

ninexnine_unit ninexnine_unit_4140(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C10K)
);

ninexnine_unit ninexnine_unit_4141(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D10K)
);

ninexnine_unit ninexnine_unit_4142(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E10K)
);

ninexnine_unit ninexnine_unit_4143(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F10K)
);

assign C110K=c1010K+c1110K+c1210K+c1310K+c1410K+c1510K+c1610K+c1710K+c1810K+c1910K+c1A10K+c1B10K+c1C10K+c1D10K+c1E10K+c1F10K;
assign A110K=(C110K>=0)?1:0;

assign P210K=A110K;

ninexnine_unit ninexnine_unit_4144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1011K)
);

ninexnine_unit ninexnine_unit_4145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1111K)
);

ninexnine_unit ninexnine_unit_4146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1211K)
);

ninexnine_unit ninexnine_unit_4147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1311K)
);

ninexnine_unit ninexnine_unit_4148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1411K)
);

ninexnine_unit ninexnine_unit_4149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1511K)
);

ninexnine_unit ninexnine_unit_4150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1611K)
);

ninexnine_unit ninexnine_unit_4151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1711K)
);

ninexnine_unit ninexnine_unit_4152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1811K)
);

ninexnine_unit ninexnine_unit_4153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1911K)
);

ninexnine_unit ninexnine_unit_4154(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A11K)
);

ninexnine_unit ninexnine_unit_4155(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B11K)
);

ninexnine_unit ninexnine_unit_4156(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C11K)
);

ninexnine_unit ninexnine_unit_4157(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D11K)
);

ninexnine_unit ninexnine_unit_4158(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E11K)
);

ninexnine_unit ninexnine_unit_4159(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F11K)
);

assign C111K=c1011K+c1111K+c1211K+c1311K+c1411K+c1511K+c1611K+c1711K+c1811K+c1911K+c1A11K+c1B11K+c1C11K+c1D11K+c1E11K+c1F11K;
assign A111K=(C111K>=0)?1:0;

assign P211K=A111K;

ninexnine_unit ninexnine_unit_4160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1012K)
);

ninexnine_unit ninexnine_unit_4161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1112K)
);

ninexnine_unit ninexnine_unit_4162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1212K)
);

ninexnine_unit ninexnine_unit_4163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1312K)
);

ninexnine_unit ninexnine_unit_4164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1412K)
);

ninexnine_unit ninexnine_unit_4165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1512K)
);

ninexnine_unit ninexnine_unit_4166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1612K)
);

ninexnine_unit ninexnine_unit_4167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1712K)
);

ninexnine_unit ninexnine_unit_4168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1812K)
);

ninexnine_unit ninexnine_unit_4169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1912K)
);

ninexnine_unit ninexnine_unit_4170(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A12K)
);

ninexnine_unit ninexnine_unit_4171(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B12K)
);

ninexnine_unit ninexnine_unit_4172(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C12K)
);

ninexnine_unit ninexnine_unit_4173(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D12K)
);

ninexnine_unit ninexnine_unit_4174(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E12K)
);

ninexnine_unit ninexnine_unit_4175(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F12K)
);

assign C112K=c1012K+c1112K+c1212K+c1312K+c1412K+c1512K+c1612K+c1712K+c1812K+c1912K+c1A12K+c1B12K+c1C12K+c1D12K+c1E12K+c1F12K;
assign A112K=(C112K>=0)?1:0;

assign P212K=A112K;

ninexnine_unit ninexnine_unit_4176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1020K)
);

ninexnine_unit ninexnine_unit_4177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1120K)
);

ninexnine_unit ninexnine_unit_4178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1220K)
);

ninexnine_unit ninexnine_unit_4179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1320K)
);

ninexnine_unit ninexnine_unit_4180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1420K)
);

ninexnine_unit ninexnine_unit_4181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1520K)
);

ninexnine_unit ninexnine_unit_4182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1620K)
);

ninexnine_unit ninexnine_unit_4183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1720K)
);

ninexnine_unit ninexnine_unit_4184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1820K)
);

ninexnine_unit ninexnine_unit_4185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1920K)
);

ninexnine_unit ninexnine_unit_4186(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A20K)
);

ninexnine_unit ninexnine_unit_4187(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B20K)
);

ninexnine_unit ninexnine_unit_4188(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C20K)
);

ninexnine_unit ninexnine_unit_4189(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D20K)
);

ninexnine_unit ninexnine_unit_4190(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E20K)
);

ninexnine_unit ninexnine_unit_4191(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F20K)
);

assign C120K=c1020K+c1120K+c1220K+c1320K+c1420K+c1520K+c1620K+c1720K+c1820K+c1920K+c1A20K+c1B20K+c1C20K+c1D20K+c1E20K+c1F20K;
assign A120K=(C120K>=0)?1:0;

assign P220K=A120K;

ninexnine_unit ninexnine_unit_4192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1021K)
);

ninexnine_unit ninexnine_unit_4193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1121K)
);

ninexnine_unit ninexnine_unit_4194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1221K)
);

ninexnine_unit ninexnine_unit_4195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1321K)
);

ninexnine_unit ninexnine_unit_4196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1421K)
);

ninexnine_unit ninexnine_unit_4197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1521K)
);

ninexnine_unit ninexnine_unit_4198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1621K)
);

ninexnine_unit ninexnine_unit_4199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1721K)
);

ninexnine_unit ninexnine_unit_4200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1821K)
);

ninexnine_unit ninexnine_unit_4201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1921K)
);

ninexnine_unit ninexnine_unit_4202(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A21K)
);

ninexnine_unit ninexnine_unit_4203(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B21K)
);

ninexnine_unit ninexnine_unit_4204(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C21K)
);

ninexnine_unit ninexnine_unit_4205(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D21K)
);

ninexnine_unit ninexnine_unit_4206(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E21K)
);

ninexnine_unit ninexnine_unit_4207(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F21K)
);

assign C121K=c1021K+c1121K+c1221K+c1321K+c1421K+c1521K+c1621K+c1721K+c1821K+c1921K+c1A21K+c1B21K+c1C21K+c1D21K+c1E21K+c1F21K;
assign A121K=(C121K>=0)?1:0;

assign P221K=A121K;

ninexnine_unit ninexnine_unit_4208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1K000),
				.b1(W1K010),
				.b2(W1K020),
				.b3(W1K100),
				.b4(W1K110),
				.b5(W1K120),
				.b6(W1K200),
				.b7(W1K210),
				.b8(W1K220),
				.c(c1022K)
);

ninexnine_unit ninexnine_unit_4209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1K001),
				.b1(W1K011),
				.b2(W1K021),
				.b3(W1K101),
				.b4(W1K111),
				.b5(W1K121),
				.b6(W1K201),
				.b7(W1K211),
				.b8(W1K221),
				.c(c1122K)
);

ninexnine_unit ninexnine_unit_4210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1K002),
				.b1(W1K012),
				.b2(W1K022),
				.b3(W1K102),
				.b4(W1K112),
				.b5(W1K122),
				.b6(W1K202),
				.b7(W1K212),
				.b8(W1K222),
				.c(c1222K)
);

ninexnine_unit ninexnine_unit_4211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1K003),
				.b1(W1K013),
				.b2(W1K023),
				.b3(W1K103),
				.b4(W1K113),
				.b5(W1K123),
				.b6(W1K203),
				.b7(W1K213),
				.b8(W1K223),
				.c(c1322K)
);

ninexnine_unit ninexnine_unit_4212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1K004),
				.b1(W1K014),
				.b2(W1K024),
				.b3(W1K104),
				.b4(W1K114),
				.b5(W1K124),
				.b6(W1K204),
				.b7(W1K214),
				.b8(W1K224),
				.c(c1422K)
);

ninexnine_unit ninexnine_unit_4213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1K005),
				.b1(W1K015),
				.b2(W1K025),
				.b3(W1K105),
				.b4(W1K115),
				.b5(W1K125),
				.b6(W1K205),
				.b7(W1K215),
				.b8(W1K225),
				.c(c1522K)
);

ninexnine_unit ninexnine_unit_4214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1K006),
				.b1(W1K016),
				.b2(W1K026),
				.b3(W1K106),
				.b4(W1K116),
				.b5(W1K126),
				.b6(W1K206),
				.b7(W1K216),
				.b8(W1K226),
				.c(c1622K)
);

ninexnine_unit ninexnine_unit_4215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1K007),
				.b1(W1K017),
				.b2(W1K027),
				.b3(W1K107),
				.b4(W1K117),
				.b5(W1K127),
				.b6(W1K207),
				.b7(W1K217),
				.b8(W1K227),
				.c(c1722K)
);

ninexnine_unit ninexnine_unit_4216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1K008),
				.b1(W1K018),
				.b2(W1K028),
				.b3(W1K108),
				.b4(W1K118),
				.b5(W1K128),
				.b6(W1K208),
				.b7(W1K218),
				.b8(W1K228),
				.c(c1822K)
);

ninexnine_unit ninexnine_unit_4217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1K009),
				.b1(W1K019),
				.b2(W1K029),
				.b3(W1K109),
				.b4(W1K119),
				.b5(W1K129),
				.b6(W1K209),
				.b7(W1K219),
				.b8(W1K229),
				.c(c1922K)
);

ninexnine_unit ninexnine_unit_4218(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1K00A),
				.b1(W1K01A),
				.b2(W1K02A),
				.b3(W1K10A),
				.b4(W1K11A),
				.b5(W1K12A),
				.b6(W1K20A),
				.b7(W1K21A),
				.b8(W1K22A),
				.c(c1A22K)
);

ninexnine_unit ninexnine_unit_4219(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1K00B),
				.b1(W1K01B),
				.b2(W1K02B),
				.b3(W1K10B),
				.b4(W1K11B),
				.b5(W1K12B),
				.b6(W1K20B),
				.b7(W1K21B),
				.b8(W1K22B),
				.c(c1B22K)
);

ninexnine_unit ninexnine_unit_4220(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1K00C),
				.b1(W1K01C),
				.b2(W1K02C),
				.b3(W1K10C),
				.b4(W1K11C),
				.b5(W1K12C),
				.b6(W1K20C),
				.b7(W1K21C),
				.b8(W1K22C),
				.c(c1C22K)
);

ninexnine_unit ninexnine_unit_4221(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1K00D),
				.b1(W1K01D),
				.b2(W1K02D),
				.b3(W1K10D),
				.b4(W1K11D),
				.b5(W1K12D),
				.b6(W1K20D),
				.b7(W1K21D),
				.b8(W1K22D),
				.c(c1D22K)
);

ninexnine_unit ninexnine_unit_4222(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1K00E),
				.b1(W1K01E),
				.b2(W1K02E),
				.b3(W1K10E),
				.b4(W1K11E),
				.b5(W1K12E),
				.b6(W1K20E),
				.b7(W1K21E),
				.b8(W1K22E),
				.c(c1E22K)
);

ninexnine_unit ninexnine_unit_4223(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1K00F),
				.b1(W1K01F),
				.b2(W1K02F),
				.b3(W1K10F),
				.b4(W1K11F),
				.b5(W1K12F),
				.b6(W1K20F),
				.b7(W1K21F),
				.b8(W1K22F),
				.c(c1F22K)
);

assign C122K=c1022K+c1122K+c1222K+c1322K+c1422K+c1522K+c1622K+c1722K+c1822K+c1922K+c1A22K+c1B22K+c1C22K+c1D22K+c1E22K+c1F22K;
assign A122K=(C122K>=0)?1:0;

assign P222K=A122K;

ninexnine_unit ninexnine_unit_4224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1000L)
);

ninexnine_unit ninexnine_unit_4225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1100L)
);

ninexnine_unit ninexnine_unit_4226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1200L)
);

ninexnine_unit ninexnine_unit_4227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1300L)
);

ninexnine_unit ninexnine_unit_4228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1400L)
);

ninexnine_unit ninexnine_unit_4229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1500L)
);

ninexnine_unit ninexnine_unit_4230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1600L)
);

ninexnine_unit ninexnine_unit_4231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1700L)
);

ninexnine_unit ninexnine_unit_4232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1800L)
);

ninexnine_unit ninexnine_unit_4233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1900L)
);

ninexnine_unit ninexnine_unit_4234(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A00L)
);

ninexnine_unit ninexnine_unit_4235(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B00L)
);

ninexnine_unit ninexnine_unit_4236(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C00L)
);

ninexnine_unit ninexnine_unit_4237(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D00L)
);

ninexnine_unit ninexnine_unit_4238(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E00L)
);

ninexnine_unit ninexnine_unit_4239(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F00L)
);

assign C100L=c1000L+c1100L+c1200L+c1300L+c1400L+c1500L+c1600L+c1700L+c1800L+c1900L+c1A00L+c1B00L+c1C00L+c1D00L+c1E00L+c1F00L;
assign A100L=(C100L>=0)?1:0;

assign P200L=A100L;

ninexnine_unit ninexnine_unit_4240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1001L)
);

ninexnine_unit ninexnine_unit_4241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1101L)
);

ninexnine_unit ninexnine_unit_4242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1201L)
);

ninexnine_unit ninexnine_unit_4243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1301L)
);

ninexnine_unit ninexnine_unit_4244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1401L)
);

ninexnine_unit ninexnine_unit_4245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1501L)
);

ninexnine_unit ninexnine_unit_4246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1601L)
);

ninexnine_unit ninexnine_unit_4247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1701L)
);

ninexnine_unit ninexnine_unit_4248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1801L)
);

ninexnine_unit ninexnine_unit_4249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1901L)
);

ninexnine_unit ninexnine_unit_4250(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A01L)
);

ninexnine_unit ninexnine_unit_4251(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B01L)
);

ninexnine_unit ninexnine_unit_4252(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C01L)
);

ninexnine_unit ninexnine_unit_4253(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D01L)
);

ninexnine_unit ninexnine_unit_4254(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E01L)
);

ninexnine_unit ninexnine_unit_4255(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F01L)
);

assign C101L=c1001L+c1101L+c1201L+c1301L+c1401L+c1501L+c1601L+c1701L+c1801L+c1901L+c1A01L+c1B01L+c1C01L+c1D01L+c1E01L+c1F01L;
assign A101L=(C101L>=0)?1:0;

assign P201L=A101L;

ninexnine_unit ninexnine_unit_4256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1002L)
);

ninexnine_unit ninexnine_unit_4257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1102L)
);

ninexnine_unit ninexnine_unit_4258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1202L)
);

ninexnine_unit ninexnine_unit_4259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1302L)
);

ninexnine_unit ninexnine_unit_4260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1402L)
);

ninexnine_unit ninexnine_unit_4261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1502L)
);

ninexnine_unit ninexnine_unit_4262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1602L)
);

ninexnine_unit ninexnine_unit_4263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1702L)
);

ninexnine_unit ninexnine_unit_4264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1802L)
);

ninexnine_unit ninexnine_unit_4265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1902L)
);

ninexnine_unit ninexnine_unit_4266(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A02L)
);

ninexnine_unit ninexnine_unit_4267(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B02L)
);

ninexnine_unit ninexnine_unit_4268(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C02L)
);

ninexnine_unit ninexnine_unit_4269(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D02L)
);

ninexnine_unit ninexnine_unit_4270(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E02L)
);

ninexnine_unit ninexnine_unit_4271(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F02L)
);

assign C102L=c1002L+c1102L+c1202L+c1302L+c1402L+c1502L+c1602L+c1702L+c1802L+c1902L+c1A02L+c1B02L+c1C02L+c1D02L+c1E02L+c1F02L;
assign A102L=(C102L>=0)?1:0;

assign P202L=A102L;

ninexnine_unit ninexnine_unit_4272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1010L)
);

ninexnine_unit ninexnine_unit_4273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1110L)
);

ninexnine_unit ninexnine_unit_4274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1210L)
);

ninexnine_unit ninexnine_unit_4275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1310L)
);

ninexnine_unit ninexnine_unit_4276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1410L)
);

ninexnine_unit ninexnine_unit_4277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1510L)
);

ninexnine_unit ninexnine_unit_4278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1610L)
);

ninexnine_unit ninexnine_unit_4279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1710L)
);

ninexnine_unit ninexnine_unit_4280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1810L)
);

ninexnine_unit ninexnine_unit_4281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1910L)
);

ninexnine_unit ninexnine_unit_4282(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A10L)
);

ninexnine_unit ninexnine_unit_4283(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B10L)
);

ninexnine_unit ninexnine_unit_4284(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C10L)
);

ninexnine_unit ninexnine_unit_4285(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D10L)
);

ninexnine_unit ninexnine_unit_4286(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E10L)
);

ninexnine_unit ninexnine_unit_4287(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F10L)
);

assign C110L=c1010L+c1110L+c1210L+c1310L+c1410L+c1510L+c1610L+c1710L+c1810L+c1910L+c1A10L+c1B10L+c1C10L+c1D10L+c1E10L+c1F10L;
assign A110L=(C110L>=0)?1:0;

assign P210L=A110L;

ninexnine_unit ninexnine_unit_4288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1011L)
);

ninexnine_unit ninexnine_unit_4289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1111L)
);

ninexnine_unit ninexnine_unit_4290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1211L)
);

ninexnine_unit ninexnine_unit_4291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1311L)
);

ninexnine_unit ninexnine_unit_4292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1411L)
);

ninexnine_unit ninexnine_unit_4293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1511L)
);

ninexnine_unit ninexnine_unit_4294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1611L)
);

ninexnine_unit ninexnine_unit_4295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1711L)
);

ninexnine_unit ninexnine_unit_4296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1811L)
);

ninexnine_unit ninexnine_unit_4297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1911L)
);

ninexnine_unit ninexnine_unit_4298(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A11L)
);

ninexnine_unit ninexnine_unit_4299(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B11L)
);

ninexnine_unit ninexnine_unit_4300(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C11L)
);

ninexnine_unit ninexnine_unit_4301(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D11L)
);

ninexnine_unit ninexnine_unit_4302(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E11L)
);

ninexnine_unit ninexnine_unit_4303(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F11L)
);

assign C111L=c1011L+c1111L+c1211L+c1311L+c1411L+c1511L+c1611L+c1711L+c1811L+c1911L+c1A11L+c1B11L+c1C11L+c1D11L+c1E11L+c1F11L;
assign A111L=(C111L>=0)?1:0;

assign P211L=A111L;

ninexnine_unit ninexnine_unit_4304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1012L)
);

ninexnine_unit ninexnine_unit_4305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1112L)
);

ninexnine_unit ninexnine_unit_4306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1212L)
);

ninexnine_unit ninexnine_unit_4307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1312L)
);

ninexnine_unit ninexnine_unit_4308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1412L)
);

ninexnine_unit ninexnine_unit_4309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1512L)
);

ninexnine_unit ninexnine_unit_4310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1612L)
);

ninexnine_unit ninexnine_unit_4311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1712L)
);

ninexnine_unit ninexnine_unit_4312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1812L)
);

ninexnine_unit ninexnine_unit_4313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1912L)
);

ninexnine_unit ninexnine_unit_4314(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A12L)
);

ninexnine_unit ninexnine_unit_4315(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B12L)
);

ninexnine_unit ninexnine_unit_4316(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C12L)
);

ninexnine_unit ninexnine_unit_4317(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D12L)
);

ninexnine_unit ninexnine_unit_4318(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E12L)
);

ninexnine_unit ninexnine_unit_4319(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F12L)
);

assign C112L=c1012L+c1112L+c1212L+c1312L+c1412L+c1512L+c1612L+c1712L+c1812L+c1912L+c1A12L+c1B12L+c1C12L+c1D12L+c1E12L+c1F12L;
assign A112L=(C112L>=0)?1:0;

assign P212L=A112L;

ninexnine_unit ninexnine_unit_4320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1020L)
);

ninexnine_unit ninexnine_unit_4321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1120L)
);

ninexnine_unit ninexnine_unit_4322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1220L)
);

ninexnine_unit ninexnine_unit_4323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1320L)
);

ninexnine_unit ninexnine_unit_4324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1420L)
);

ninexnine_unit ninexnine_unit_4325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1520L)
);

ninexnine_unit ninexnine_unit_4326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1620L)
);

ninexnine_unit ninexnine_unit_4327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1720L)
);

ninexnine_unit ninexnine_unit_4328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1820L)
);

ninexnine_unit ninexnine_unit_4329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1920L)
);

ninexnine_unit ninexnine_unit_4330(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A20L)
);

ninexnine_unit ninexnine_unit_4331(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B20L)
);

ninexnine_unit ninexnine_unit_4332(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C20L)
);

ninexnine_unit ninexnine_unit_4333(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D20L)
);

ninexnine_unit ninexnine_unit_4334(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E20L)
);

ninexnine_unit ninexnine_unit_4335(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F20L)
);

assign C120L=c1020L+c1120L+c1220L+c1320L+c1420L+c1520L+c1620L+c1720L+c1820L+c1920L+c1A20L+c1B20L+c1C20L+c1D20L+c1E20L+c1F20L;
assign A120L=(C120L>=0)?1:0;

assign P220L=A120L;

ninexnine_unit ninexnine_unit_4336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1021L)
);

ninexnine_unit ninexnine_unit_4337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1121L)
);

ninexnine_unit ninexnine_unit_4338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1221L)
);

ninexnine_unit ninexnine_unit_4339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1321L)
);

ninexnine_unit ninexnine_unit_4340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1421L)
);

ninexnine_unit ninexnine_unit_4341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1521L)
);

ninexnine_unit ninexnine_unit_4342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1621L)
);

ninexnine_unit ninexnine_unit_4343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1721L)
);

ninexnine_unit ninexnine_unit_4344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1821L)
);

ninexnine_unit ninexnine_unit_4345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1921L)
);

ninexnine_unit ninexnine_unit_4346(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A21L)
);

ninexnine_unit ninexnine_unit_4347(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B21L)
);

ninexnine_unit ninexnine_unit_4348(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C21L)
);

ninexnine_unit ninexnine_unit_4349(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D21L)
);

ninexnine_unit ninexnine_unit_4350(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E21L)
);

ninexnine_unit ninexnine_unit_4351(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F21L)
);

assign C121L=c1021L+c1121L+c1221L+c1321L+c1421L+c1521L+c1621L+c1721L+c1821L+c1921L+c1A21L+c1B21L+c1C21L+c1D21L+c1E21L+c1F21L;
assign A121L=(C121L>=0)?1:0;

assign P221L=A121L;

ninexnine_unit ninexnine_unit_4352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1L000),
				.b1(W1L010),
				.b2(W1L020),
				.b3(W1L100),
				.b4(W1L110),
				.b5(W1L120),
				.b6(W1L200),
				.b7(W1L210),
				.b8(W1L220),
				.c(c1022L)
);

ninexnine_unit ninexnine_unit_4353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1L001),
				.b1(W1L011),
				.b2(W1L021),
				.b3(W1L101),
				.b4(W1L111),
				.b5(W1L121),
				.b6(W1L201),
				.b7(W1L211),
				.b8(W1L221),
				.c(c1122L)
);

ninexnine_unit ninexnine_unit_4354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1L002),
				.b1(W1L012),
				.b2(W1L022),
				.b3(W1L102),
				.b4(W1L112),
				.b5(W1L122),
				.b6(W1L202),
				.b7(W1L212),
				.b8(W1L222),
				.c(c1222L)
);

ninexnine_unit ninexnine_unit_4355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1L003),
				.b1(W1L013),
				.b2(W1L023),
				.b3(W1L103),
				.b4(W1L113),
				.b5(W1L123),
				.b6(W1L203),
				.b7(W1L213),
				.b8(W1L223),
				.c(c1322L)
);

ninexnine_unit ninexnine_unit_4356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1L004),
				.b1(W1L014),
				.b2(W1L024),
				.b3(W1L104),
				.b4(W1L114),
				.b5(W1L124),
				.b6(W1L204),
				.b7(W1L214),
				.b8(W1L224),
				.c(c1422L)
);

ninexnine_unit ninexnine_unit_4357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1L005),
				.b1(W1L015),
				.b2(W1L025),
				.b3(W1L105),
				.b4(W1L115),
				.b5(W1L125),
				.b6(W1L205),
				.b7(W1L215),
				.b8(W1L225),
				.c(c1522L)
);

ninexnine_unit ninexnine_unit_4358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1L006),
				.b1(W1L016),
				.b2(W1L026),
				.b3(W1L106),
				.b4(W1L116),
				.b5(W1L126),
				.b6(W1L206),
				.b7(W1L216),
				.b8(W1L226),
				.c(c1622L)
);

ninexnine_unit ninexnine_unit_4359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1L007),
				.b1(W1L017),
				.b2(W1L027),
				.b3(W1L107),
				.b4(W1L117),
				.b5(W1L127),
				.b6(W1L207),
				.b7(W1L217),
				.b8(W1L227),
				.c(c1722L)
);

ninexnine_unit ninexnine_unit_4360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1L008),
				.b1(W1L018),
				.b2(W1L028),
				.b3(W1L108),
				.b4(W1L118),
				.b5(W1L128),
				.b6(W1L208),
				.b7(W1L218),
				.b8(W1L228),
				.c(c1822L)
);

ninexnine_unit ninexnine_unit_4361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1L009),
				.b1(W1L019),
				.b2(W1L029),
				.b3(W1L109),
				.b4(W1L119),
				.b5(W1L129),
				.b6(W1L209),
				.b7(W1L219),
				.b8(W1L229),
				.c(c1922L)
);

ninexnine_unit ninexnine_unit_4362(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1L00A),
				.b1(W1L01A),
				.b2(W1L02A),
				.b3(W1L10A),
				.b4(W1L11A),
				.b5(W1L12A),
				.b6(W1L20A),
				.b7(W1L21A),
				.b8(W1L22A),
				.c(c1A22L)
);

ninexnine_unit ninexnine_unit_4363(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1L00B),
				.b1(W1L01B),
				.b2(W1L02B),
				.b3(W1L10B),
				.b4(W1L11B),
				.b5(W1L12B),
				.b6(W1L20B),
				.b7(W1L21B),
				.b8(W1L22B),
				.c(c1B22L)
);

ninexnine_unit ninexnine_unit_4364(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1L00C),
				.b1(W1L01C),
				.b2(W1L02C),
				.b3(W1L10C),
				.b4(W1L11C),
				.b5(W1L12C),
				.b6(W1L20C),
				.b7(W1L21C),
				.b8(W1L22C),
				.c(c1C22L)
);

ninexnine_unit ninexnine_unit_4365(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1L00D),
				.b1(W1L01D),
				.b2(W1L02D),
				.b3(W1L10D),
				.b4(W1L11D),
				.b5(W1L12D),
				.b6(W1L20D),
				.b7(W1L21D),
				.b8(W1L22D),
				.c(c1D22L)
);

ninexnine_unit ninexnine_unit_4366(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1L00E),
				.b1(W1L01E),
				.b2(W1L02E),
				.b3(W1L10E),
				.b4(W1L11E),
				.b5(W1L12E),
				.b6(W1L20E),
				.b7(W1L21E),
				.b8(W1L22E),
				.c(c1E22L)
);

ninexnine_unit ninexnine_unit_4367(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1L00F),
				.b1(W1L01F),
				.b2(W1L02F),
				.b3(W1L10F),
				.b4(W1L11F),
				.b5(W1L12F),
				.b6(W1L20F),
				.b7(W1L21F),
				.b8(W1L22F),
				.c(c1F22L)
);

assign C122L=c1022L+c1122L+c1222L+c1322L+c1422L+c1522L+c1622L+c1722L+c1822L+c1922L+c1A22L+c1B22L+c1C22L+c1D22L+c1E22L+c1F22L;
assign A122L=(C122L>=0)?1:0;

assign P222L=A122L;

ninexnine_unit ninexnine_unit_4368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1000M)
);

ninexnine_unit ninexnine_unit_4369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1100M)
);

ninexnine_unit ninexnine_unit_4370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1200M)
);

ninexnine_unit ninexnine_unit_4371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1300M)
);

ninexnine_unit ninexnine_unit_4372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1004),
				.a1(P1014),
				.a2(P1024),
				.a3(P1104),
				.a4(P1114),
				.a5(P1124),
				.a6(P1204),
				.a7(P1214),
				.a8(P1224),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1400M)
);

ninexnine_unit ninexnine_unit_4373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1005),
				.a1(P1015),
				.a2(P1025),
				.a3(P1105),
				.a4(P1115),
				.a5(P1125),
				.a6(P1205),
				.a7(P1215),
				.a8(P1225),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1500M)
);

ninexnine_unit ninexnine_unit_4374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1006),
				.a1(P1016),
				.a2(P1026),
				.a3(P1106),
				.a4(P1116),
				.a5(P1126),
				.a6(P1206),
				.a7(P1216),
				.a8(P1226),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1600M)
);

ninexnine_unit ninexnine_unit_4375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1007),
				.a1(P1017),
				.a2(P1027),
				.a3(P1107),
				.a4(P1117),
				.a5(P1127),
				.a6(P1207),
				.a7(P1217),
				.a8(P1227),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1700M)
);

ninexnine_unit ninexnine_unit_4376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1008),
				.a1(P1018),
				.a2(P1028),
				.a3(P1108),
				.a4(P1118),
				.a5(P1128),
				.a6(P1208),
				.a7(P1218),
				.a8(P1228),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1800M)
);

ninexnine_unit ninexnine_unit_4377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1009),
				.a1(P1019),
				.a2(P1029),
				.a3(P1109),
				.a4(P1119),
				.a5(P1129),
				.a6(P1209),
				.a7(P1219),
				.a8(P1229),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1900M)
);

ninexnine_unit ninexnine_unit_4378(
				.clk(clk),
				.rstn(rstn),
				.a0(P100A),
				.a1(P101A),
				.a2(P102A),
				.a3(P110A),
				.a4(P111A),
				.a5(P112A),
				.a6(P120A),
				.a7(P121A),
				.a8(P122A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A00M)
);

ninexnine_unit ninexnine_unit_4379(
				.clk(clk),
				.rstn(rstn),
				.a0(P100B),
				.a1(P101B),
				.a2(P102B),
				.a3(P110B),
				.a4(P111B),
				.a5(P112B),
				.a6(P120B),
				.a7(P121B),
				.a8(P122B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B00M)
);

ninexnine_unit ninexnine_unit_4380(
				.clk(clk),
				.rstn(rstn),
				.a0(P100C),
				.a1(P101C),
				.a2(P102C),
				.a3(P110C),
				.a4(P111C),
				.a5(P112C),
				.a6(P120C),
				.a7(P121C),
				.a8(P122C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C00M)
);

ninexnine_unit ninexnine_unit_4381(
				.clk(clk),
				.rstn(rstn),
				.a0(P100D),
				.a1(P101D),
				.a2(P102D),
				.a3(P110D),
				.a4(P111D),
				.a5(P112D),
				.a6(P120D),
				.a7(P121D),
				.a8(P122D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D00M)
);

ninexnine_unit ninexnine_unit_4382(
				.clk(clk),
				.rstn(rstn),
				.a0(P100E),
				.a1(P101E),
				.a2(P102E),
				.a3(P110E),
				.a4(P111E),
				.a5(P112E),
				.a6(P120E),
				.a7(P121E),
				.a8(P122E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E00M)
);

ninexnine_unit ninexnine_unit_4383(
				.clk(clk),
				.rstn(rstn),
				.a0(P100F),
				.a1(P101F),
				.a2(P102F),
				.a3(P110F),
				.a4(P111F),
				.a5(P112F),
				.a6(P120F),
				.a7(P121F),
				.a8(P122F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F00M)
);

assign C100M=c1000M+c1100M+c1200M+c1300M+c1400M+c1500M+c1600M+c1700M+c1800M+c1900M+c1A00M+c1B00M+c1C00M+c1D00M+c1E00M+c1F00M;
assign A100M=(C100M>=0)?1:0;

assign P200M=A100M;

ninexnine_unit ninexnine_unit_4384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1001M)
);

ninexnine_unit ninexnine_unit_4385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1101M)
);

ninexnine_unit ninexnine_unit_4386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1201M)
);

ninexnine_unit ninexnine_unit_4387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1301M)
);

ninexnine_unit ninexnine_unit_4388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1014),
				.a1(P1024),
				.a2(P1034),
				.a3(P1114),
				.a4(P1124),
				.a5(P1134),
				.a6(P1214),
				.a7(P1224),
				.a8(P1234),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1401M)
);

ninexnine_unit ninexnine_unit_4389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1015),
				.a1(P1025),
				.a2(P1035),
				.a3(P1115),
				.a4(P1125),
				.a5(P1135),
				.a6(P1215),
				.a7(P1225),
				.a8(P1235),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1501M)
);

ninexnine_unit ninexnine_unit_4390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1016),
				.a1(P1026),
				.a2(P1036),
				.a3(P1116),
				.a4(P1126),
				.a5(P1136),
				.a6(P1216),
				.a7(P1226),
				.a8(P1236),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1601M)
);

ninexnine_unit ninexnine_unit_4391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1017),
				.a1(P1027),
				.a2(P1037),
				.a3(P1117),
				.a4(P1127),
				.a5(P1137),
				.a6(P1217),
				.a7(P1227),
				.a8(P1237),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1701M)
);

ninexnine_unit ninexnine_unit_4392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1018),
				.a1(P1028),
				.a2(P1038),
				.a3(P1118),
				.a4(P1128),
				.a5(P1138),
				.a6(P1218),
				.a7(P1228),
				.a8(P1238),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1801M)
);

ninexnine_unit ninexnine_unit_4393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1019),
				.a1(P1029),
				.a2(P1039),
				.a3(P1119),
				.a4(P1129),
				.a5(P1139),
				.a6(P1219),
				.a7(P1229),
				.a8(P1239),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1901M)
);

ninexnine_unit ninexnine_unit_4394(
				.clk(clk),
				.rstn(rstn),
				.a0(P101A),
				.a1(P102A),
				.a2(P103A),
				.a3(P111A),
				.a4(P112A),
				.a5(P113A),
				.a6(P121A),
				.a7(P122A),
				.a8(P123A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A01M)
);

ninexnine_unit ninexnine_unit_4395(
				.clk(clk),
				.rstn(rstn),
				.a0(P101B),
				.a1(P102B),
				.a2(P103B),
				.a3(P111B),
				.a4(P112B),
				.a5(P113B),
				.a6(P121B),
				.a7(P122B),
				.a8(P123B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B01M)
);

ninexnine_unit ninexnine_unit_4396(
				.clk(clk),
				.rstn(rstn),
				.a0(P101C),
				.a1(P102C),
				.a2(P103C),
				.a3(P111C),
				.a4(P112C),
				.a5(P113C),
				.a6(P121C),
				.a7(P122C),
				.a8(P123C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C01M)
);

ninexnine_unit ninexnine_unit_4397(
				.clk(clk),
				.rstn(rstn),
				.a0(P101D),
				.a1(P102D),
				.a2(P103D),
				.a3(P111D),
				.a4(P112D),
				.a5(P113D),
				.a6(P121D),
				.a7(P122D),
				.a8(P123D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D01M)
);

ninexnine_unit ninexnine_unit_4398(
				.clk(clk),
				.rstn(rstn),
				.a0(P101E),
				.a1(P102E),
				.a2(P103E),
				.a3(P111E),
				.a4(P112E),
				.a5(P113E),
				.a6(P121E),
				.a7(P122E),
				.a8(P123E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E01M)
);

ninexnine_unit ninexnine_unit_4399(
				.clk(clk),
				.rstn(rstn),
				.a0(P101F),
				.a1(P102F),
				.a2(P103F),
				.a3(P111F),
				.a4(P112F),
				.a5(P113F),
				.a6(P121F),
				.a7(P122F),
				.a8(P123F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F01M)
);

assign C101M=c1001M+c1101M+c1201M+c1301M+c1401M+c1501M+c1601M+c1701M+c1801M+c1901M+c1A01M+c1B01M+c1C01M+c1D01M+c1E01M+c1F01M;
assign A101M=(C101M>=0)?1:0;

assign P201M=A101M;

ninexnine_unit ninexnine_unit_4400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1002M)
);

ninexnine_unit ninexnine_unit_4401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1102M)
);

ninexnine_unit ninexnine_unit_4402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1202M)
);

ninexnine_unit ninexnine_unit_4403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1023),
				.a1(P1033),
				.a2(P1043),
				.a3(P1123),
				.a4(P1133),
				.a5(P1143),
				.a6(P1223),
				.a7(P1233),
				.a8(P1243),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1302M)
);

ninexnine_unit ninexnine_unit_4404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1024),
				.a1(P1034),
				.a2(P1044),
				.a3(P1124),
				.a4(P1134),
				.a5(P1144),
				.a6(P1224),
				.a7(P1234),
				.a8(P1244),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1402M)
);

ninexnine_unit ninexnine_unit_4405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1025),
				.a1(P1035),
				.a2(P1045),
				.a3(P1125),
				.a4(P1135),
				.a5(P1145),
				.a6(P1225),
				.a7(P1235),
				.a8(P1245),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1502M)
);

ninexnine_unit ninexnine_unit_4406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1026),
				.a1(P1036),
				.a2(P1046),
				.a3(P1126),
				.a4(P1136),
				.a5(P1146),
				.a6(P1226),
				.a7(P1236),
				.a8(P1246),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1602M)
);

ninexnine_unit ninexnine_unit_4407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1027),
				.a1(P1037),
				.a2(P1047),
				.a3(P1127),
				.a4(P1137),
				.a5(P1147),
				.a6(P1227),
				.a7(P1237),
				.a8(P1247),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1702M)
);

ninexnine_unit ninexnine_unit_4408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1028),
				.a1(P1038),
				.a2(P1048),
				.a3(P1128),
				.a4(P1138),
				.a5(P1148),
				.a6(P1228),
				.a7(P1238),
				.a8(P1248),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1802M)
);

ninexnine_unit ninexnine_unit_4409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1029),
				.a1(P1039),
				.a2(P1049),
				.a3(P1129),
				.a4(P1139),
				.a5(P1149),
				.a6(P1229),
				.a7(P1239),
				.a8(P1249),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1902M)
);

ninexnine_unit ninexnine_unit_4410(
				.clk(clk),
				.rstn(rstn),
				.a0(P102A),
				.a1(P103A),
				.a2(P104A),
				.a3(P112A),
				.a4(P113A),
				.a5(P114A),
				.a6(P122A),
				.a7(P123A),
				.a8(P124A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A02M)
);

ninexnine_unit ninexnine_unit_4411(
				.clk(clk),
				.rstn(rstn),
				.a0(P102B),
				.a1(P103B),
				.a2(P104B),
				.a3(P112B),
				.a4(P113B),
				.a5(P114B),
				.a6(P122B),
				.a7(P123B),
				.a8(P124B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B02M)
);

ninexnine_unit ninexnine_unit_4412(
				.clk(clk),
				.rstn(rstn),
				.a0(P102C),
				.a1(P103C),
				.a2(P104C),
				.a3(P112C),
				.a4(P113C),
				.a5(P114C),
				.a6(P122C),
				.a7(P123C),
				.a8(P124C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C02M)
);

ninexnine_unit ninexnine_unit_4413(
				.clk(clk),
				.rstn(rstn),
				.a0(P102D),
				.a1(P103D),
				.a2(P104D),
				.a3(P112D),
				.a4(P113D),
				.a5(P114D),
				.a6(P122D),
				.a7(P123D),
				.a8(P124D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D02M)
);

ninexnine_unit ninexnine_unit_4414(
				.clk(clk),
				.rstn(rstn),
				.a0(P102E),
				.a1(P103E),
				.a2(P104E),
				.a3(P112E),
				.a4(P113E),
				.a5(P114E),
				.a6(P122E),
				.a7(P123E),
				.a8(P124E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E02M)
);

ninexnine_unit ninexnine_unit_4415(
				.clk(clk),
				.rstn(rstn),
				.a0(P102F),
				.a1(P103F),
				.a2(P104F),
				.a3(P112F),
				.a4(P113F),
				.a5(P114F),
				.a6(P122F),
				.a7(P123F),
				.a8(P124F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F02M)
);

assign C102M=c1002M+c1102M+c1202M+c1302M+c1402M+c1502M+c1602M+c1702M+c1802M+c1902M+c1A02M+c1B02M+c1C02M+c1D02M+c1E02M+c1F02M;
assign A102M=(C102M>=0)?1:0;

assign P202M=A102M;

ninexnine_unit ninexnine_unit_4416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1010M)
);

ninexnine_unit ninexnine_unit_4417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1110M)
);

ninexnine_unit ninexnine_unit_4418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1210M)
);

ninexnine_unit ninexnine_unit_4419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1310M)
);

ninexnine_unit ninexnine_unit_4420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1104),
				.a1(P1114),
				.a2(P1124),
				.a3(P1204),
				.a4(P1214),
				.a5(P1224),
				.a6(P1304),
				.a7(P1314),
				.a8(P1324),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1410M)
);

ninexnine_unit ninexnine_unit_4421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1105),
				.a1(P1115),
				.a2(P1125),
				.a3(P1205),
				.a4(P1215),
				.a5(P1225),
				.a6(P1305),
				.a7(P1315),
				.a8(P1325),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1510M)
);

ninexnine_unit ninexnine_unit_4422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1106),
				.a1(P1116),
				.a2(P1126),
				.a3(P1206),
				.a4(P1216),
				.a5(P1226),
				.a6(P1306),
				.a7(P1316),
				.a8(P1326),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1610M)
);

ninexnine_unit ninexnine_unit_4423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1107),
				.a1(P1117),
				.a2(P1127),
				.a3(P1207),
				.a4(P1217),
				.a5(P1227),
				.a6(P1307),
				.a7(P1317),
				.a8(P1327),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1710M)
);

ninexnine_unit ninexnine_unit_4424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1108),
				.a1(P1118),
				.a2(P1128),
				.a3(P1208),
				.a4(P1218),
				.a5(P1228),
				.a6(P1308),
				.a7(P1318),
				.a8(P1328),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1810M)
);

ninexnine_unit ninexnine_unit_4425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1109),
				.a1(P1119),
				.a2(P1129),
				.a3(P1209),
				.a4(P1219),
				.a5(P1229),
				.a6(P1309),
				.a7(P1319),
				.a8(P1329),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1910M)
);

ninexnine_unit ninexnine_unit_4426(
				.clk(clk),
				.rstn(rstn),
				.a0(P110A),
				.a1(P111A),
				.a2(P112A),
				.a3(P120A),
				.a4(P121A),
				.a5(P122A),
				.a6(P130A),
				.a7(P131A),
				.a8(P132A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A10M)
);

ninexnine_unit ninexnine_unit_4427(
				.clk(clk),
				.rstn(rstn),
				.a0(P110B),
				.a1(P111B),
				.a2(P112B),
				.a3(P120B),
				.a4(P121B),
				.a5(P122B),
				.a6(P130B),
				.a7(P131B),
				.a8(P132B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B10M)
);

ninexnine_unit ninexnine_unit_4428(
				.clk(clk),
				.rstn(rstn),
				.a0(P110C),
				.a1(P111C),
				.a2(P112C),
				.a3(P120C),
				.a4(P121C),
				.a5(P122C),
				.a6(P130C),
				.a7(P131C),
				.a8(P132C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C10M)
);

ninexnine_unit ninexnine_unit_4429(
				.clk(clk),
				.rstn(rstn),
				.a0(P110D),
				.a1(P111D),
				.a2(P112D),
				.a3(P120D),
				.a4(P121D),
				.a5(P122D),
				.a6(P130D),
				.a7(P131D),
				.a8(P132D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D10M)
);

ninexnine_unit ninexnine_unit_4430(
				.clk(clk),
				.rstn(rstn),
				.a0(P110E),
				.a1(P111E),
				.a2(P112E),
				.a3(P120E),
				.a4(P121E),
				.a5(P122E),
				.a6(P130E),
				.a7(P131E),
				.a8(P132E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E10M)
);

ninexnine_unit ninexnine_unit_4431(
				.clk(clk),
				.rstn(rstn),
				.a0(P110F),
				.a1(P111F),
				.a2(P112F),
				.a3(P120F),
				.a4(P121F),
				.a5(P122F),
				.a6(P130F),
				.a7(P131F),
				.a8(P132F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F10M)
);

assign C110M=c1010M+c1110M+c1210M+c1310M+c1410M+c1510M+c1610M+c1710M+c1810M+c1910M+c1A10M+c1B10M+c1C10M+c1D10M+c1E10M+c1F10M;
assign A110M=(C110M>=0)?1:0;

assign P210M=A110M;

ninexnine_unit ninexnine_unit_4432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1011M)
);

ninexnine_unit ninexnine_unit_4433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1111M)
);

ninexnine_unit ninexnine_unit_4434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1211M)
);

ninexnine_unit ninexnine_unit_4435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1311M)
);

ninexnine_unit ninexnine_unit_4436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1114),
				.a1(P1124),
				.a2(P1134),
				.a3(P1214),
				.a4(P1224),
				.a5(P1234),
				.a6(P1314),
				.a7(P1324),
				.a8(P1334),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1411M)
);

ninexnine_unit ninexnine_unit_4437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1115),
				.a1(P1125),
				.a2(P1135),
				.a3(P1215),
				.a4(P1225),
				.a5(P1235),
				.a6(P1315),
				.a7(P1325),
				.a8(P1335),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1511M)
);

ninexnine_unit ninexnine_unit_4438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1116),
				.a1(P1126),
				.a2(P1136),
				.a3(P1216),
				.a4(P1226),
				.a5(P1236),
				.a6(P1316),
				.a7(P1326),
				.a8(P1336),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1611M)
);

ninexnine_unit ninexnine_unit_4439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1117),
				.a1(P1127),
				.a2(P1137),
				.a3(P1217),
				.a4(P1227),
				.a5(P1237),
				.a6(P1317),
				.a7(P1327),
				.a8(P1337),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1711M)
);

ninexnine_unit ninexnine_unit_4440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1118),
				.a1(P1128),
				.a2(P1138),
				.a3(P1218),
				.a4(P1228),
				.a5(P1238),
				.a6(P1318),
				.a7(P1328),
				.a8(P1338),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1811M)
);

ninexnine_unit ninexnine_unit_4441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1119),
				.a1(P1129),
				.a2(P1139),
				.a3(P1219),
				.a4(P1229),
				.a5(P1239),
				.a6(P1319),
				.a7(P1329),
				.a8(P1339),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1911M)
);

ninexnine_unit ninexnine_unit_4442(
				.clk(clk),
				.rstn(rstn),
				.a0(P111A),
				.a1(P112A),
				.a2(P113A),
				.a3(P121A),
				.a4(P122A),
				.a5(P123A),
				.a6(P131A),
				.a7(P132A),
				.a8(P133A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A11M)
);

ninexnine_unit ninexnine_unit_4443(
				.clk(clk),
				.rstn(rstn),
				.a0(P111B),
				.a1(P112B),
				.a2(P113B),
				.a3(P121B),
				.a4(P122B),
				.a5(P123B),
				.a6(P131B),
				.a7(P132B),
				.a8(P133B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B11M)
);

ninexnine_unit ninexnine_unit_4444(
				.clk(clk),
				.rstn(rstn),
				.a0(P111C),
				.a1(P112C),
				.a2(P113C),
				.a3(P121C),
				.a4(P122C),
				.a5(P123C),
				.a6(P131C),
				.a7(P132C),
				.a8(P133C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C11M)
);

ninexnine_unit ninexnine_unit_4445(
				.clk(clk),
				.rstn(rstn),
				.a0(P111D),
				.a1(P112D),
				.a2(P113D),
				.a3(P121D),
				.a4(P122D),
				.a5(P123D),
				.a6(P131D),
				.a7(P132D),
				.a8(P133D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D11M)
);

ninexnine_unit ninexnine_unit_4446(
				.clk(clk),
				.rstn(rstn),
				.a0(P111E),
				.a1(P112E),
				.a2(P113E),
				.a3(P121E),
				.a4(P122E),
				.a5(P123E),
				.a6(P131E),
				.a7(P132E),
				.a8(P133E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E11M)
);

ninexnine_unit ninexnine_unit_4447(
				.clk(clk),
				.rstn(rstn),
				.a0(P111F),
				.a1(P112F),
				.a2(P113F),
				.a3(P121F),
				.a4(P122F),
				.a5(P123F),
				.a6(P131F),
				.a7(P132F),
				.a8(P133F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F11M)
);

assign C111M=c1011M+c1111M+c1211M+c1311M+c1411M+c1511M+c1611M+c1711M+c1811M+c1911M+c1A11M+c1B11M+c1C11M+c1D11M+c1E11M+c1F11M;
assign A111M=(C111M>=0)?1:0;

assign P211M=A111M;

ninexnine_unit ninexnine_unit_4448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1012M)
);

ninexnine_unit ninexnine_unit_4449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1112M)
);

ninexnine_unit ninexnine_unit_4450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1212M)
);

ninexnine_unit ninexnine_unit_4451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1123),
				.a1(P1133),
				.a2(P1143),
				.a3(P1223),
				.a4(P1233),
				.a5(P1243),
				.a6(P1323),
				.a7(P1333),
				.a8(P1343),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1312M)
);

ninexnine_unit ninexnine_unit_4452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1124),
				.a1(P1134),
				.a2(P1144),
				.a3(P1224),
				.a4(P1234),
				.a5(P1244),
				.a6(P1324),
				.a7(P1334),
				.a8(P1344),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1412M)
);

ninexnine_unit ninexnine_unit_4453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1125),
				.a1(P1135),
				.a2(P1145),
				.a3(P1225),
				.a4(P1235),
				.a5(P1245),
				.a6(P1325),
				.a7(P1335),
				.a8(P1345),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1512M)
);

ninexnine_unit ninexnine_unit_4454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1126),
				.a1(P1136),
				.a2(P1146),
				.a3(P1226),
				.a4(P1236),
				.a5(P1246),
				.a6(P1326),
				.a7(P1336),
				.a8(P1346),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1612M)
);

ninexnine_unit ninexnine_unit_4455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1127),
				.a1(P1137),
				.a2(P1147),
				.a3(P1227),
				.a4(P1237),
				.a5(P1247),
				.a6(P1327),
				.a7(P1337),
				.a8(P1347),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1712M)
);

ninexnine_unit ninexnine_unit_4456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1128),
				.a1(P1138),
				.a2(P1148),
				.a3(P1228),
				.a4(P1238),
				.a5(P1248),
				.a6(P1328),
				.a7(P1338),
				.a8(P1348),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1812M)
);

ninexnine_unit ninexnine_unit_4457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1129),
				.a1(P1139),
				.a2(P1149),
				.a3(P1229),
				.a4(P1239),
				.a5(P1249),
				.a6(P1329),
				.a7(P1339),
				.a8(P1349),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1912M)
);

ninexnine_unit ninexnine_unit_4458(
				.clk(clk),
				.rstn(rstn),
				.a0(P112A),
				.a1(P113A),
				.a2(P114A),
				.a3(P122A),
				.a4(P123A),
				.a5(P124A),
				.a6(P132A),
				.a7(P133A),
				.a8(P134A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A12M)
);

ninexnine_unit ninexnine_unit_4459(
				.clk(clk),
				.rstn(rstn),
				.a0(P112B),
				.a1(P113B),
				.a2(P114B),
				.a3(P122B),
				.a4(P123B),
				.a5(P124B),
				.a6(P132B),
				.a7(P133B),
				.a8(P134B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B12M)
);

ninexnine_unit ninexnine_unit_4460(
				.clk(clk),
				.rstn(rstn),
				.a0(P112C),
				.a1(P113C),
				.a2(P114C),
				.a3(P122C),
				.a4(P123C),
				.a5(P124C),
				.a6(P132C),
				.a7(P133C),
				.a8(P134C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C12M)
);

ninexnine_unit ninexnine_unit_4461(
				.clk(clk),
				.rstn(rstn),
				.a0(P112D),
				.a1(P113D),
				.a2(P114D),
				.a3(P122D),
				.a4(P123D),
				.a5(P124D),
				.a6(P132D),
				.a7(P133D),
				.a8(P134D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D12M)
);

ninexnine_unit ninexnine_unit_4462(
				.clk(clk),
				.rstn(rstn),
				.a0(P112E),
				.a1(P113E),
				.a2(P114E),
				.a3(P122E),
				.a4(P123E),
				.a5(P124E),
				.a6(P132E),
				.a7(P133E),
				.a8(P134E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E12M)
);

ninexnine_unit ninexnine_unit_4463(
				.clk(clk),
				.rstn(rstn),
				.a0(P112F),
				.a1(P113F),
				.a2(P114F),
				.a3(P122F),
				.a4(P123F),
				.a5(P124F),
				.a6(P132F),
				.a7(P133F),
				.a8(P134F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F12M)
);

assign C112M=c1012M+c1112M+c1212M+c1312M+c1412M+c1512M+c1612M+c1712M+c1812M+c1912M+c1A12M+c1B12M+c1C12M+c1D12M+c1E12M+c1F12M;
assign A112M=(C112M>=0)?1:0;

assign P212M=A112M;

ninexnine_unit ninexnine_unit_4464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1020M)
);

ninexnine_unit ninexnine_unit_4465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1120M)
);

ninexnine_unit ninexnine_unit_4466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1220M)
);

ninexnine_unit ninexnine_unit_4467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1203),
				.a1(P1213),
				.a2(P1223),
				.a3(P1303),
				.a4(P1313),
				.a5(P1323),
				.a6(P1403),
				.a7(P1413),
				.a8(P1423),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1320M)
);

ninexnine_unit ninexnine_unit_4468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1204),
				.a1(P1214),
				.a2(P1224),
				.a3(P1304),
				.a4(P1314),
				.a5(P1324),
				.a6(P1404),
				.a7(P1414),
				.a8(P1424),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1420M)
);

ninexnine_unit ninexnine_unit_4469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1205),
				.a1(P1215),
				.a2(P1225),
				.a3(P1305),
				.a4(P1315),
				.a5(P1325),
				.a6(P1405),
				.a7(P1415),
				.a8(P1425),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1520M)
);

ninexnine_unit ninexnine_unit_4470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1206),
				.a1(P1216),
				.a2(P1226),
				.a3(P1306),
				.a4(P1316),
				.a5(P1326),
				.a6(P1406),
				.a7(P1416),
				.a8(P1426),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1620M)
);

ninexnine_unit ninexnine_unit_4471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1207),
				.a1(P1217),
				.a2(P1227),
				.a3(P1307),
				.a4(P1317),
				.a5(P1327),
				.a6(P1407),
				.a7(P1417),
				.a8(P1427),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1720M)
);

ninexnine_unit ninexnine_unit_4472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1208),
				.a1(P1218),
				.a2(P1228),
				.a3(P1308),
				.a4(P1318),
				.a5(P1328),
				.a6(P1408),
				.a7(P1418),
				.a8(P1428),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1820M)
);

ninexnine_unit ninexnine_unit_4473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1209),
				.a1(P1219),
				.a2(P1229),
				.a3(P1309),
				.a4(P1319),
				.a5(P1329),
				.a6(P1409),
				.a7(P1419),
				.a8(P1429),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1920M)
);

ninexnine_unit ninexnine_unit_4474(
				.clk(clk),
				.rstn(rstn),
				.a0(P120A),
				.a1(P121A),
				.a2(P122A),
				.a3(P130A),
				.a4(P131A),
				.a5(P132A),
				.a6(P140A),
				.a7(P141A),
				.a8(P142A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A20M)
);

ninexnine_unit ninexnine_unit_4475(
				.clk(clk),
				.rstn(rstn),
				.a0(P120B),
				.a1(P121B),
				.a2(P122B),
				.a3(P130B),
				.a4(P131B),
				.a5(P132B),
				.a6(P140B),
				.a7(P141B),
				.a8(P142B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B20M)
);

ninexnine_unit ninexnine_unit_4476(
				.clk(clk),
				.rstn(rstn),
				.a0(P120C),
				.a1(P121C),
				.a2(P122C),
				.a3(P130C),
				.a4(P131C),
				.a5(P132C),
				.a6(P140C),
				.a7(P141C),
				.a8(P142C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C20M)
);

ninexnine_unit ninexnine_unit_4477(
				.clk(clk),
				.rstn(rstn),
				.a0(P120D),
				.a1(P121D),
				.a2(P122D),
				.a3(P130D),
				.a4(P131D),
				.a5(P132D),
				.a6(P140D),
				.a7(P141D),
				.a8(P142D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D20M)
);

ninexnine_unit ninexnine_unit_4478(
				.clk(clk),
				.rstn(rstn),
				.a0(P120E),
				.a1(P121E),
				.a2(P122E),
				.a3(P130E),
				.a4(P131E),
				.a5(P132E),
				.a6(P140E),
				.a7(P141E),
				.a8(P142E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E20M)
);

ninexnine_unit ninexnine_unit_4479(
				.clk(clk),
				.rstn(rstn),
				.a0(P120F),
				.a1(P121F),
				.a2(P122F),
				.a3(P130F),
				.a4(P131F),
				.a5(P132F),
				.a6(P140F),
				.a7(P141F),
				.a8(P142F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F20M)
);

assign C120M=c1020M+c1120M+c1220M+c1320M+c1420M+c1520M+c1620M+c1720M+c1820M+c1920M+c1A20M+c1B20M+c1C20M+c1D20M+c1E20M+c1F20M;
assign A120M=(C120M>=0)?1:0;

assign P220M=A120M;

ninexnine_unit ninexnine_unit_4480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1021M)
);

ninexnine_unit ninexnine_unit_4481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1121M)
);

ninexnine_unit ninexnine_unit_4482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1221M)
);

ninexnine_unit ninexnine_unit_4483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1213),
				.a1(P1223),
				.a2(P1233),
				.a3(P1313),
				.a4(P1323),
				.a5(P1333),
				.a6(P1413),
				.a7(P1423),
				.a8(P1433),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1321M)
);

ninexnine_unit ninexnine_unit_4484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1214),
				.a1(P1224),
				.a2(P1234),
				.a3(P1314),
				.a4(P1324),
				.a5(P1334),
				.a6(P1414),
				.a7(P1424),
				.a8(P1434),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1421M)
);

ninexnine_unit ninexnine_unit_4485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1215),
				.a1(P1225),
				.a2(P1235),
				.a3(P1315),
				.a4(P1325),
				.a5(P1335),
				.a6(P1415),
				.a7(P1425),
				.a8(P1435),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1521M)
);

ninexnine_unit ninexnine_unit_4486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1216),
				.a1(P1226),
				.a2(P1236),
				.a3(P1316),
				.a4(P1326),
				.a5(P1336),
				.a6(P1416),
				.a7(P1426),
				.a8(P1436),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1621M)
);

ninexnine_unit ninexnine_unit_4487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1217),
				.a1(P1227),
				.a2(P1237),
				.a3(P1317),
				.a4(P1327),
				.a5(P1337),
				.a6(P1417),
				.a7(P1427),
				.a8(P1437),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1721M)
);

ninexnine_unit ninexnine_unit_4488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1218),
				.a1(P1228),
				.a2(P1238),
				.a3(P1318),
				.a4(P1328),
				.a5(P1338),
				.a6(P1418),
				.a7(P1428),
				.a8(P1438),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1821M)
);

ninexnine_unit ninexnine_unit_4489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1219),
				.a1(P1229),
				.a2(P1239),
				.a3(P1319),
				.a4(P1329),
				.a5(P1339),
				.a6(P1419),
				.a7(P1429),
				.a8(P1439),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1921M)
);

ninexnine_unit ninexnine_unit_4490(
				.clk(clk),
				.rstn(rstn),
				.a0(P121A),
				.a1(P122A),
				.a2(P123A),
				.a3(P131A),
				.a4(P132A),
				.a5(P133A),
				.a6(P141A),
				.a7(P142A),
				.a8(P143A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A21M)
);

ninexnine_unit ninexnine_unit_4491(
				.clk(clk),
				.rstn(rstn),
				.a0(P121B),
				.a1(P122B),
				.a2(P123B),
				.a3(P131B),
				.a4(P132B),
				.a5(P133B),
				.a6(P141B),
				.a7(P142B),
				.a8(P143B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B21M)
);

ninexnine_unit ninexnine_unit_4492(
				.clk(clk),
				.rstn(rstn),
				.a0(P121C),
				.a1(P122C),
				.a2(P123C),
				.a3(P131C),
				.a4(P132C),
				.a5(P133C),
				.a6(P141C),
				.a7(P142C),
				.a8(P143C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C21M)
);

ninexnine_unit ninexnine_unit_4493(
				.clk(clk),
				.rstn(rstn),
				.a0(P121D),
				.a1(P122D),
				.a2(P123D),
				.a3(P131D),
				.a4(P132D),
				.a5(P133D),
				.a6(P141D),
				.a7(P142D),
				.a8(P143D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D21M)
);

ninexnine_unit ninexnine_unit_4494(
				.clk(clk),
				.rstn(rstn),
				.a0(P121E),
				.a1(P122E),
				.a2(P123E),
				.a3(P131E),
				.a4(P132E),
				.a5(P133E),
				.a6(P141E),
				.a7(P142E),
				.a8(P143E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E21M)
);

ninexnine_unit ninexnine_unit_4495(
				.clk(clk),
				.rstn(rstn),
				.a0(P121F),
				.a1(P122F),
				.a2(P123F),
				.a3(P131F),
				.a4(P132F),
				.a5(P133F),
				.a6(P141F),
				.a7(P142F),
				.a8(P143F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F21M)
);

assign C121M=c1021M+c1121M+c1221M+c1321M+c1421M+c1521M+c1621M+c1721M+c1821M+c1921M+c1A21M+c1B21M+c1C21M+c1D21M+c1E21M+c1F21M;
assign A121M=(C121M>=0)?1:0;

assign P221M=A121M;

ninexnine_unit ninexnine_unit_4496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1M000),
				.b1(W1M010),
				.b2(W1M020),
				.b3(W1M100),
				.b4(W1M110),
				.b5(W1M120),
				.b6(W1M200),
				.b7(W1M210),
				.b8(W1M220),
				.c(c1022M)
);

ninexnine_unit ninexnine_unit_4497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1M001),
				.b1(W1M011),
				.b2(W1M021),
				.b3(W1M101),
				.b4(W1M111),
				.b5(W1M121),
				.b6(W1M201),
				.b7(W1M211),
				.b8(W1M221),
				.c(c1122M)
);

ninexnine_unit ninexnine_unit_4498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1M002),
				.b1(W1M012),
				.b2(W1M022),
				.b3(W1M102),
				.b4(W1M112),
				.b5(W1M122),
				.b6(W1M202),
				.b7(W1M212),
				.b8(W1M222),
				.c(c1222M)
);

ninexnine_unit ninexnine_unit_4499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1223),
				.a1(P1233),
				.a2(P1243),
				.a3(P1323),
				.a4(P1333),
				.a5(P1343),
				.a6(P1423),
				.a7(P1433),
				.a8(P1443),
				.b0(W1M003),
				.b1(W1M013),
				.b2(W1M023),
				.b3(W1M103),
				.b4(W1M113),
				.b5(W1M123),
				.b6(W1M203),
				.b7(W1M213),
				.b8(W1M223),
				.c(c1322M)
);

ninexnine_unit ninexnine_unit_4500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1224),
				.a1(P1234),
				.a2(P1244),
				.a3(P1324),
				.a4(P1334),
				.a5(P1344),
				.a6(P1424),
				.a7(P1434),
				.a8(P1444),
				.b0(W1M004),
				.b1(W1M014),
				.b2(W1M024),
				.b3(W1M104),
				.b4(W1M114),
				.b5(W1M124),
				.b6(W1M204),
				.b7(W1M214),
				.b8(W1M224),
				.c(c1422M)
);

ninexnine_unit ninexnine_unit_4501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1225),
				.a1(P1235),
				.a2(P1245),
				.a3(P1325),
				.a4(P1335),
				.a5(P1345),
				.a6(P1425),
				.a7(P1435),
				.a8(P1445),
				.b0(W1M005),
				.b1(W1M015),
				.b2(W1M025),
				.b3(W1M105),
				.b4(W1M115),
				.b5(W1M125),
				.b6(W1M205),
				.b7(W1M215),
				.b8(W1M225),
				.c(c1522M)
);

ninexnine_unit ninexnine_unit_4502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1226),
				.a1(P1236),
				.a2(P1246),
				.a3(P1326),
				.a4(P1336),
				.a5(P1346),
				.a6(P1426),
				.a7(P1436),
				.a8(P1446),
				.b0(W1M006),
				.b1(W1M016),
				.b2(W1M026),
				.b3(W1M106),
				.b4(W1M116),
				.b5(W1M126),
				.b6(W1M206),
				.b7(W1M216),
				.b8(W1M226),
				.c(c1622M)
);

ninexnine_unit ninexnine_unit_4503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1227),
				.a1(P1237),
				.a2(P1247),
				.a3(P1327),
				.a4(P1337),
				.a5(P1347),
				.a6(P1427),
				.a7(P1437),
				.a8(P1447),
				.b0(W1M007),
				.b1(W1M017),
				.b2(W1M027),
				.b3(W1M107),
				.b4(W1M117),
				.b5(W1M127),
				.b6(W1M207),
				.b7(W1M217),
				.b8(W1M227),
				.c(c1722M)
);

ninexnine_unit ninexnine_unit_4504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1228),
				.a1(P1238),
				.a2(P1248),
				.a3(P1328),
				.a4(P1338),
				.a5(P1348),
				.a6(P1428),
				.a7(P1438),
				.a8(P1448),
				.b0(W1M008),
				.b1(W1M018),
				.b2(W1M028),
				.b3(W1M108),
				.b4(W1M118),
				.b5(W1M128),
				.b6(W1M208),
				.b7(W1M218),
				.b8(W1M228),
				.c(c1822M)
);

ninexnine_unit ninexnine_unit_4505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1229),
				.a1(P1239),
				.a2(P1249),
				.a3(P1329),
				.a4(P1339),
				.a5(P1349),
				.a6(P1429),
				.a7(P1439),
				.a8(P1449),
				.b0(W1M009),
				.b1(W1M019),
				.b2(W1M029),
				.b3(W1M109),
				.b4(W1M119),
				.b5(W1M129),
				.b6(W1M209),
				.b7(W1M219),
				.b8(W1M229),
				.c(c1922M)
);

ninexnine_unit ninexnine_unit_4506(
				.clk(clk),
				.rstn(rstn),
				.a0(P122A),
				.a1(P123A),
				.a2(P124A),
				.a3(P132A),
				.a4(P133A),
				.a5(P134A),
				.a6(P142A),
				.a7(P143A),
				.a8(P144A),
				.b0(W1M00A),
				.b1(W1M01A),
				.b2(W1M02A),
				.b3(W1M10A),
				.b4(W1M11A),
				.b5(W1M12A),
				.b6(W1M20A),
				.b7(W1M21A),
				.b8(W1M22A),
				.c(c1A22M)
);

ninexnine_unit ninexnine_unit_4507(
				.clk(clk),
				.rstn(rstn),
				.a0(P122B),
				.a1(P123B),
				.a2(P124B),
				.a3(P132B),
				.a4(P133B),
				.a5(P134B),
				.a6(P142B),
				.a7(P143B),
				.a8(P144B),
				.b0(W1M00B),
				.b1(W1M01B),
				.b2(W1M02B),
				.b3(W1M10B),
				.b4(W1M11B),
				.b5(W1M12B),
				.b6(W1M20B),
				.b7(W1M21B),
				.b8(W1M22B),
				.c(c1B22M)
);

ninexnine_unit ninexnine_unit_4508(
				.clk(clk),
				.rstn(rstn),
				.a0(P122C),
				.a1(P123C),
				.a2(P124C),
				.a3(P132C),
				.a4(P133C),
				.a5(P134C),
				.a6(P142C),
				.a7(P143C),
				.a8(P144C),
				.b0(W1M00C),
				.b1(W1M01C),
				.b2(W1M02C),
				.b3(W1M10C),
				.b4(W1M11C),
				.b5(W1M12C),
				.b6(W1M20C),
				.b7(W1M21C),
				.b8(W1M22C),
				.c(c1C22M)
);

ninexnine_unit ninexnine_unit_4509(
				.clk(clk),
				.rstn(rstn),
				.a0(P122D),
				.a1(P123D),
				.a2(P124D),
				.a3(P132D),
				.a4(P133D),
				.a5(P134D),
				.a6(P142D),
				.a7(P143D),
				.a8(P144D),
				.b0(W1M00D),
				.b1(W1M01D),
				.b2(W1M02D),
				.b3(W1M10D),
				.b4(W1M11D),
				.b5(W1M12D),
				.b6(W1M20D),
				.b7(W1M21D),
				.b8(W1M22D),
				.c(c1D22M)
);

ninexnine_unit ninexnine_unit_4510(
				.clk(clk),
				.rstn(rstn),
				.a0(P122E),
				.a1(P123E),
				.a2(P124E),
				.a3(P132E),
				.a4(P133E),
				.a5(P134E),
				.a6(P142E),
				.a7(P143E),
				.a8(P144E),
				.b0(W1M00E),
				.b1(W1M01E),
				.b2(W1M02E),
				.b3(W1M10E),
				.b4(W1M11E),
				.b5(W1M12E),
				.b6(W1M20E),
				.b7(W1M21E),
				.b8(W1M22E),
				.c(c1E22M)
);

ninexnine_unit ninexnine_unit_4511(
				.clk(clk),
				.rstn(rstn),
				.a0(P122F),
				.a1(P123F),
				.a2(P124F),
				.a3(P132F),
				.a4(P133F),
				.a5(P134F),
				.a6(P142F),
				.a7(P143F),
				.a8(P144F),
				.b0(W1M00F),
				.b1(W1M01F),
				.b2(W1M02F),
				.b3(W1M10F),
				.b4(W1M11F),
				.b5(W1M12F),
				.b6(W1M20F),
				.b7(W1M21F),
				.b8(W1M22F),
				.c(c1F22M)
);

assign C122M=c1022M+c1122M+c1222M+c1322M+c1422M+c1522M+c1622M+c1722M+c1822M+c1922M+c1A22M+c1B22M+c1C22M+c1D22M+c1E22M+c1F22M;
assign A122M=(C122M>=0)?1:0;

assign P222M=A122M;

//layer3 done, begain next layer
wire P3000;
wire P3001;
wire W20000,W20010,W20020,W20100,W20110,W20120,W20200,W20210,W20220;
wire W20001,W20011,W20021,W20101,W20111,W20121,W20201,W20211,W20221;
wire W20002,W20012,W20022,W20102,W20112,W20122,W20202,W20212,W20222;
wire W20003,W20013,W20023,W20103,W20113,W20123,W20203,W20213,W20223;
wire W20004,W20014,W20024,W20104,W20114,W20124,W20204,W20214,W20224;
wire W20005,W20015,W20025,W20105,W20115,W20125,W20205,W20215,W20225;
wire W20006,W20016,W20026,W20106,W20116,W20126,W20206,W20216,W20226;
wire W20007,W20017,W20027,W20107,W20117,W20127,W20207,W20217,W20227;
wire W20008,W20018,W20028,W20108,W20118,W20128,W20208,W20218,W20228;
wire W20009,W20019,W20029,W20109,W20119,W20129,W20209,W20219,W20229;
wire W2000A,W2001A,W2002A,W2010A,W2011A,W2012A,W2020A,W2021A,W2022A;
wire W2000B,W2001B,W2002B,W2010B,W2011B,W2012B,W2020B,W2021B,W2022B;
wire W2000C,W2001C,W2002C,W2010C,W2011C,W2012C,W2020C,W2021C,W2022C;
wire W2000D,W2001D,W2002D,W2010D,W2011D,W2012D,W2020D,W2021D,W2022D;
wire W2000E,W2001E,W2002E,W2010E,W2011E,W2012E,W2020E,W2021E,W2022E;
wire W2000F,W2001F,W2002F,W2010F,W2011F,W2012F,W2020F,W2021F,W2022F;
wire W2000G,W2001G,W2002G,W2010G,W2011G,W2012G,W2020G,W2021G,W2022G;
wire W2000H,W2001H,W2002H,W2010H,W2011H,W2012H,W2020H,W2021H,W2022H;
wire W2000I,W2001I,W2002I,W2010I,W2011I,W2012I,W2020I,W2021I,W2022I;
wire W2000J,W2001J,W2002J,W2010J,W2011J,W2012J,W2020J,W2021J,W2022J;
wire W2000K,W2001K,W2002K,W2010K,W2011K,W2012K,W2020K,W2021K,W2022K;
wire W2000L,W2001L,W2002L,W2010L,W2011L,W2012L,W2020L,W2021L,W2022L;
wire W2000M,W2001M,W2002M,W2010M,W2011M,W2012M,W2020M,W2021M,W2022M;
wire W21000,W21010,W21020,W21100,W21110,W21120,W21200,W21210,W21220;
wire W21001,W21011,W21021,W21101,W21111,W21121,W21201,W21211,W21221;
wire W21002,W21012,W21022,W21102,W21112,W21122,W21202,W21212,W21222;
wire W21003,W21013,W21023,W21103,W21113,W21123,W21203,W21213,W21223;
wire W21004,W21014,W21024,W21104,W21114,W21124,W21204,W21214,W21224;
wire W21005,W21015,W21025,W21105,W21115,W21125,W21205,W21215,W21225;
wire W21006,W21016,W21026,W21106,W21116,W21126,W21206,W21216,W21226;
wire W21007,W21017,W21027,W21107,W21117,W21127,W21207,W21217,W21227;
wire W21008,W21018,W21028,W21108,W21118,W21128,W21208,W21218,W21228;
wire W21009,W21019,W21029,W21109,W21119,W21129,W21209,W21219,W21229;
wire W2100A,W2101A,W2102A,W2110A,W2111A,W2112A,W2120A,W2121A,W2122A;
wire W2100B,W2101B,W2102B,W2110B,W2111B,W2112B,W2120B,W2121B,W2122B;
wire W2100C,W2101C,W2102C,W2110C,W2111C,W2112C,W2120C,W2121C,W2122C;
wire W2100D,W2101D,W2102D,W2110D,W2111D,W2112D,W2120D,W2121D,W2122D;
wire W2100E,W2101E,W2102E,W2110E,W2111E,W2112E,W2120E,W2121E,W2122E;
wire W2100F,W2101F,W2102F,W2110F,W2111F,W2112F,W2120F,W2121F,W2122F;
wire W2100G,W2101G,W2102G,W2110G,W2111G,W2112G,W2120G,W2121G,W2122G;
wire W2100H,W2101H,W2102H,W2110H,W2111H,W2112H,W2120H,W2121H,W2122H;
wire W2100I,W2101I,W2102I,W2110I,W2111I,W2112I,W2120I,W2121I,W2122I;
wire W2100J,W2101J,W2102J,W2110J,W2111J,W2112J,W2120J,W2121J,W2122J;
wire W2100K,W2101K,W2102K,W2110K,W2111K,W2112K,W2120K,W2121K,W2122K;
wire W2100L,W2101L,W2102L,W2110L,W2111L,W2112L,W2120L,W2121L,W2122L;
wire W2100M,W2101M,W2102M,W2110M,W2111M,W2112M,W2120M,W2121M,W2122M;
wire signed [4:0] c20000,c21000,c22000,c23000,c24000,c25000,c26000,c27000,c28000,c29000,c2A000,c2B000,c2C000,c2D000,c2E000,c2F000,c2G000,c2H000,c2I000,c2J000,c2K000,c2L000,c2M000;
wire signed [4:0] c20001,c21001,c22001,c23001,c24001,c25001,c26001,c27001,c28001,c29001,c2A001,c2B001,c2C001,c2D001,c2E001,c2F001,c2G001,c2H001,c2I001,c2J001,c2K001,c2L001,c2M001;
wire signed [9:0] C2000;
wire A2000;
wire signed [9:0] C2001;
wire A2001;
DFF_save_fm DFF_W3744(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20000));
DFF_save_fm DFF_W3745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20010));
DFF_save_fm DFF_W3746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20020));
DFF_save_fm DFF_W3747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20100));
DFF_save_fm DFF_W3748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20110));
DFF_save_fm DFF_W3749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20120));
DFF_save_fm DFF_W3750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20200));
DFF_save_fm DFF_W3751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20210));
DFF_save_fm DFF_W3752(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20220));
DFF_save_fm DFF_W3753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20001));
DFF_save_fm DFF_W3754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20011));
DFF_save_fm DFF_W3755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20021));
DFF_save_fm DFF_W3756(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20101));
DFF_save_fm DFF_W3757(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20111));
DFF_save_fm DFF_W3758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20121));
DFF_save_fm DFF_W3759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20201));
DFF_save_fm DFF_W3760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20211));
DFF_save_fm DFF_W3761(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20221));
DFF_save_fm DFF_W3762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20002));
DFF_save_fm DFF_W3763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20012));
DFF_save_fm DFF_W3764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20022));
DFF_save_fm DFF_W3765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20102));
DFF_save_fm DFF_W3766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20112));
DFF_save_fm DFF_W3767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20122));
DFF_save_fm DFF_W3768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20202));
DFF_save_fm DFF_W3769(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20212));
DFF_save_fm DFF_W3770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20222));
DFF_save_fm DFF_W3771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20003));
DFF_save_fm DFF_W3772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20013));
DFF_save_fm DFF_W3773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20023));
DFF_save_fm DFF_W3774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20103));
DFF_save_fm DFF_W3775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20113));
DFF_save_fm DFF_W3776(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20123));
DFF_save_fm DFF_W3777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20203));
DFF_save_fm DFF_W3778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20213));
DFF_save_fm DFF_W3779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20223));
DFF_save_fm DFF_W3780(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20004));
DFF_save_fm DFF_W3781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20014));
DFF_save_fm DFF_W3782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20024));
DFF_save_fm DFF_W3783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20104));
DFF_save_fm DFF_W3784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20114));
DFF_save_fm DFF_W3785(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20124));
DFF_save_fm DFF_W3786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20204));
DFF_save_fm DFF_W3787(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20214));
DFF_save_fm DFF_W3788(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20224));
DFF_save_fm DFF_W3789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20005));
DFF_save_fm DFF_W3790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20015));
DFF_save_fm DFF_W3791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20025));
DFF_save_fm DFF_W3792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20105));
DFF_save_fm DFF_W3793(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20115));
DFF_save_fm DFF_W3794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20125));
DFF_save_fm DFF_W3795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20205));
DFF_save_fm DFF_W3796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20215));
DFF_save_fm DFF_W3797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20225));
DFF_save_fm DFF_W3798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20006));
DFF_save_fm DFF_W3799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20016));
DFF_save_fm DFF_W3800(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20026));
DFF_save_fm DFF_W3801(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20106));
DFF_save_fm DFF_W3802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20116));
DFF_save_fm DFF_W3803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20126));
DFF_save_fm DFF_W3804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20206));
DFF_save_fm DFF_W3805(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20216));
DFF_save_fm DFF_W3806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20226));
DFF_save_fm DFF_W3807(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20007));
DFF_save_fm DFF_W3808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20017));
DFF_save_fm DFF_W3809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20027));
DFF_save_fm DFF_W3810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20107));
DFF_save_fm DFF_W3811(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20117));
DFF_save_fm DFF_W3812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20127));
DFF_save_fm DFF_W3813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20207));
DFF_save_fm DFF_W3814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20217));
DFF_save_fm DFF_W3815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20227));
DFF_save_fm DFF_W3816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20008));
DFF_save_fm DFF_W3817(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20018));
DFF_save_fm DFF_W3818(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20028));
DFF_save_fm DFF_W3819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20108));
DFF_save_fm DFF_W3820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20118));
DFF_save_fm DFF_W3821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20128));
DFF_save_fm DFF_W3822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20208));
DFF_save_fm DFF_W3823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20218));
DFF_save_fm DFF_W3824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20228));
DFF_save_fm DFF_W3825(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20009));
DFF_save_fm DFF_W3826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20019));
DFF_save_fm DFF_W3827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20029));
DFF_save_fm DFF_W3828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20109));
DFF_save_fm DFF_W3829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20119));
DFF_save_fm DFF_W3830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20129));
DFF_save_fm DFF_W3831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20209));
DFF_save_fm DFF_W3832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20219));
DFF_save_fm DFF_W3833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20229));
DFF_save_fm DFF_W3834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000A));
DFF_save_fm DFF_W3835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001A));
DFF_save_fm DFF_W3836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002A));
DFF_save_fm DFF_W3837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010A));
DFF_save_fm DFF_W3838(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011A));
DFF_save_fm DFF_W3839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012A));
DFF_save_fm DFF_W3840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020A));
DFF_save_fm DFF_W3841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021A));
DFF_save_fm DFF_W3842(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2022A));
DFF_save_fm DFF_W3843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000B));
DFF_save_fm DFF_W3844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001B));
DFF_save_fm DFF_W3845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002B));
DFF_save_fm DFF_W3846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010B));
DFF_save_fm DFF_W3847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011B));
DFF_save_fm DFF_W3848(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012B));
DFF_save_fm DFF_W3849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020B));
DFF_save_fm DFF_W3850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021B));
DFF_save_fm DFF_W3851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022B));
DFF_save_fm DFF_W3852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000C));
DFF_save_fm DFF_W3853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001C));
DFF_save_fm DFF_W3854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002C));
DFF_save_fm DFF_W3855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010C));
DFF_save_fm DFF_W3856(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011C));
DFF_save_fm DFF_W3857(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012C));
DFF_save_fm DFF_W3858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020C));
DFF_save_fm DFF_W3859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021C));
DFF_save_fm DFF_W3860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2022C));
DFF_save_fm DFF_W3861(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000D));
DFF_save_fm DFF_W3862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001D));
DFF_save_fm DFF_W3863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002D));
DFF_save_fm DFF_W3864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010D));
DFF_save_fm DFF_W3865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011D));
DFF_save_fm DFF_W3866(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012D));
DFF_save_fm DFF_W3867(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020D));
DFF_save_fm DFF_W3868(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021D));
DFF_save_fm DFF_W3869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022D));
DFF_save_fm DFF_W3870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000E));
DFF_save_fm DFF_W3871(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001E));
DFF_save_fm DFF_W3872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002E));
DFF_save_fm DFF_W3873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010E));
DFF_save_fm DFF_W3874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011E));
DFF_save_fm DFF_W3875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012E));
DFF_save_fm DFF_W3876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020E));
DFF_save_fm DFF_W3877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021E));
DFF_save_fm DFF_W3878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022E));
DFF_save_fm DFF_W3879(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000F));
DFF_save_fm DFF_W3880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001F));
DFF_save_fm DFF_W3881(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002F));
DFF_save_fm DFF_W3882(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010F));
DFF_save_fm DFF_W3883(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011F));
DFF_save_fm DFF_W3884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012F));
DFF_save_fm DFF_W3885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020F));
DFF_save_fm DFF_W3886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021F));
DFF_save_fm DFF_W3887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022F));
DFF_save_fm DFF_W3888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000G));
DFF_save_fm DFF_W3889(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001G));
DFF_save_fm DFF_W3890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002G));
DFF_save_fm DFF_W3891(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010G));
DFF_save_fm DFF_W3892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011G));
DFF_save_fm DFF_W3893(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012G));
DFF_save_fm DFF_W3894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020G));
DFF_save_fm DFF_W3895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021G));
DFF_save_fm DFF_W3896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022G));
DFF_save_fm DFF_W3897(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000H));
DFF_save_fm DFF_W3898(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001H));
DFF_save_fm DFF_W3899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002H));
DFF_save_fm DFF_W3900(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010H));
DFF_save_fm DFF_W3901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011H));
DFF_save_fm DFF_W3902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012H));
DFF_save_fm DFF_W3903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020H));
DFF_save_fm DFF_W3904(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021H));
DFF_save_fm DFF_W3905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022H));
DFF_save_fm DFF_W3906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000I));
DFF_save_fm DFF_W3907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001I));
DFF_save_fm DFF_W3908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002I));
DFF_save_fm DFF_W3909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010I));
DFF_save_fm DFF_W3910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011I));
DFF_save_fm DFF_W3911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012I));
DFF_save_fm DFF_W3912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020I));
DFF_save_fm DFF_W3913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021I));
DFF_save_fm DFF_W3914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2022I));
DFF_save_fm DFF_W3915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000J));
DFF_save_fm DFF_W3916(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001J));
DFF_save_fm DFF_W3917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002J));
DFF_save_fm DFF_W3918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010J));
DFF_save_fm DFF_W3919(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011J));
DFF_save_fm DFF_W3920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012J));
DFF_save_fm DFF_W3921(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020J));
DFF_save_fm DFF_W3922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021J));
DFF_save_fm DFF_W3923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022J));
DFF_save_fm DFF_W3924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000K));
DFF_save_fm DFF_W3925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001K));
DFF_save_fm DFF_W3926(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002K));
DFF_save_fm DFF_W3927(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010K));
DFF_save_fm DFF_W3928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011K));
DFF_save_fm DFF_W3929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012K));
DFF_save_fm DFF_W3930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020K));
DFF_save_fm DFF_W3931(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021K));
DFF_save_fm DFF_W3932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022K));
DFF_save_fm DFF_W3933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000L));
DFF_save_fm DFF_W3934(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001L));
DFF_save_fm DFF_W3935(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002L));
DFF_save_fm DFF_W3936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010L));
DFF_save_fm DFF_W3937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011L));
DFF_save_fm DFF_W3938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012L));
DFF_save_fm DFF_W3939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020L));
DFF_save_fm DFF_W3940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021L));
DFF_save_fm DFF_W3941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022L));
DFF_save_fm DFF_W3942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000M));
DFF_save_fm DFF_W3943(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001M));
DFF_save_fm DFF_W3944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002M));
DFF_save_fm DFF_W3945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010M));
DFF_save_fm DFF_W3946(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011M));
DFF_save_fm DFF_W3947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012M));
DFF_save_fm DFF_W3948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020M));
DFF_save_fm DFF_W3949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021M));
DFF_save_fm DFF_W3950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022M));
DFF_save_fm DFF_W3951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21000));
DFF_save_fm DFF_W3952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21010));
DFF_save_fm DFF_W3953(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21020));
DFF_save_fm DFF_W3954(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21100));
DFF_save_fm DFF_W3955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21110));
DFF_save_fm DFF_W3956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21120));
DFF_save_fm DFF_W3957(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21200));
DFF_save_fm DFF_W3958(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21210));
DFF_save_fm DFF_W3959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21220));
DFF_save_fm DFF_W3960(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21001));
DFF_save_fm DFF_W3961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21011));
DFF_save_fm DFF_W3962(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21021));
DFF_save_fm DFF_W3963(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21101));
DFF_save_fm DFF_W3964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21111));
DFF_save_fm DFF_W3965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21121));
DFF_save_fm DFF_W3966(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21201));
DFF_save_fm DFF_W3967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21211));
DFF_save_fm DFF_W3968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21221));
DFF_save_fm DFF_W3969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21002));
DFF_save_fm DFF_W3970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21012));
DFF_save_fm DFF_W3971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21022));
DFF_save_fm DFF_W3972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21102));
DFF_save_fm DFF_W3973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21112));
DFF_save_fm DFF_W3974(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21122));
DFF_save_fm DFF_W3975(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21202));
DFF_save_fm DFF_W3976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21212));
DFF_save_fm DFF_W3977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21222));
DFF_save_fm DFF_W3978(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21003));
DFF_save_fm DFF_W3979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21013));
DFF_save_fm DFF_W3980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21023));
DFF_save_fm DFF_W3981(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21103));
DFF_save_fm DFF_W3982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21113));
DFF_save_fm DFF_W3983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21123));
DFF_save_fm DFF_W3984(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21203));
DFF_save_fm DFF_W3985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21213));
DFF_save_fm DFF_W3986(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21223));
DFF_save_fm DFF_W3987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21004));
DFF_save_fm DFF_W3988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21014));
DFF_save_fm DFF_W3989(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21024));
DFF_save_fm DFF_W3990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21104));
DFF_save_fm DFF_W3991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21114));
DFF_save_fm DFF_W3992(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21124));
DFF_save_fm DFF_W3993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21204));
DFF_save_fm DFF_W3994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21214));
DFF_save_fm DFF_W3995(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21224));
DFF_save_fm DFF_W3996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21005));
DFF_save_fm DFF_W3997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21015));
DFF_save_fm DFF_W3998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21025));
DFF_save_fm DFF_W3999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21105));
DFF_save_fm DFF_W4000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21115));
DFF_save_fm DFF_W4001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21125));
DFF_save_fm DFF_W4002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21205));
DFF_save_fm DFF_W4003(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21215));
DFF_save_fm DFF_W4004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21225));
DFF_save_fm DFF_W4005(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21006));
DFF_save_fm DFF_W4006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21016));
DFF_save_fm DFF_W4007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21026));
DFF_save_fm DFF_W4008(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21106));
DFF_save_fm DFF_W4009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21116));
DFF_save_fm DFF_W4010(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21126));
DFF_save_fm DFF_W4011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21206));
DFF_save_fm DFF_W4012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21216));
DFF_save_fm DFF_W4013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21226));
DFF_save_fm DFF_W4014(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21007));
DFF_save_fm DFF_W4015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21017));
DFF_save_fm DFF_W4016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21027));
DFF_save_fm DFF_W4017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21107));
DFF_save_fm DFF_W4018(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21117));
DFF_save_fm DFF_W4019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21127));
DFF_save_fm DFF_W4020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21207));
DFF_save_fm DFF_W4021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21217));
DFF_save_fm DFF_W4022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21227));
DFF_save_fm DFF_W4023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21008));
DFF_save_fm DFF_W4024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21018));
DFF_save_fm DFF_W4025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21028));
DFF_save_fm DFF_W4026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21108));
DFF_save_fm DFF_W4027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21118));
DFF_save_fm DFF_W4028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21128));
DFF_save_fm DFF_W4029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21208));
DFF_save_fm DFF_W4030(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21218));
DFF_save_fm DFF_W4031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21228));
DFF_save_fm DFF_W4032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21009));
DFF_save_fm DFF_W4033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21019));
DFF_save_fm DFF_W4034(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21029));
DFF_save_fm DFF_W4035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21109));
DFF_save_fm DFF_W4036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21119));
DFF_save_fm DFF_W4037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21129));
DFF_save_fm DFF_W4038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21209));
DFF_save_fm DFF_W4039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21219));
DFF_save_fm DFF_W4040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21229));
DFF_save_fm DFF_W4041(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100A));
DFF_save_fm DFF_W4042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101A));
DFF_save_fm DFF_W4043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102A));
DFF_save_fm DFF_W4044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110A));
DFF_save_fm DFF_W4045(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111A));
DFF_save_fm DFF_W4046(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112A));
DFF_save_fm DFF_W4047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120A));
DFF_save_fm DFF_W4048(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121A));
DFF_save_fm DFF_W4049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122A));
DFF_save_fm DFF_W4050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100B));
DFF_save_fm DFF_W4051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101B));
DFF_save_fm DFF_W4052(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102B));
DFF_save_fm DFF_W4053(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110B));
DFF_save_fm DFF_W4054(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111B));
DFF_save_fm DFF_W4055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112B));
DFF_save_fm DFF_W4056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120B));
DFF_save_fm DFF_W4057(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121B));
DFF_save_fm DFF_W4058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122B));
DFF_save_fm DFF_W4059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100C));
DFF_save_fm DFF_W4060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101C));
DFF_save_fm DFF_W4061(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102C));
DFF_save_fm DFF_W4062(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110C));
DFF_save_fm DFF_W4063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111C));
DFF_save_fm DFF_W4064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112C));
DFF_save_fm DFF_W4065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120C));
DFF_save_fm DFF_W4066(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121C));
DFF_save_fm DFF_W4067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122C));
DFF_save_fm DFF_W4068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100D));
DFF_save_fm DFF_W4069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101D));
DFF_save_fm DFF_W4070(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102D));
DFF_save_fm DFF_W4071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110D));
DFF_save_fm DFF_W4072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111D));
DFF_save_fm DFF_W4073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112D));
DFF_save_fm DFF_W4074(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120D));
DFF_save_fm DFF_W4075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121D));
DFF_save_fm DFF_W4076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122D));
DFF_save_fm DFF_W4077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100E));
DFF_save_fm DFF_W4078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101E));
DFF_save_fm DFF_W4079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102E));
DFF_save_fm DFF_W4080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110E));
DFF_save_fm DFF_W4081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111E));
DFF_save_fm DFF_W4082(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112E));
DFF_save_fm DFF_W4083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120E));
DFF_save_fm DFF_W4084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121E));
DFF_save_fm DFF_W4085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122E));
DFF_save_fm DFF_W4086(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100F));
DFF_save_fm DFF_W4087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101F));
DFF_save_fm DFF_W4088(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102F));
DFF_save_fm DFF_W4089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110F));
DFF_save_fm DFF_W4090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111F));
DFF_save_fm DFF_W4091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112F));
DFF_save_fm DFF_W4092(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120F));
DFF_save_fm DFF_W4093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121F));
DFF_save_fm DFF_W4094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122F));
DFF_save_fm DFF_W4095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100G));
DFF_save_fm DFF_W4096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101G));
DFF_save_fm DFF_W4097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102G));
DFF_save_fm DFF_W4098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110G));
DFF_save_fm DFF_W4099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111G));
DFF_save_fm DFF_W4100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112G));
DFF_save_fm DFF_W4101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120G));
DFF_save_fm DFF_W4102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121G));
DFF_save_fm DFF_W4103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122G));
DFF_save_fm DFF_W4104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100H));
DFF_save_fm DFF_W4105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101H));
DFF_save_fm DFF_W4106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102H));
DFF_save_fm DFF_W4107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110H));
DFF_save_fm DFF_W4108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111H));
DFF_save_fm DFF_W4109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112H));
DFF_save_fm DFF_W4110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120H));
DFF_save_fm DFF_W4111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121H));
DFF_save_fm DFF_W4112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122H));
DFF_save_fm DFF_W4113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100I));
DFF_save_fm DFF_W4114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101I));
DFF_save_fm DFF_W4115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102I));
DFF_save_fm DFF_W4116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110I));
DFF_save_fm DFF_W4117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111I));
DFF_save_fm DFF_W4118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112I));
DFF_save_fm DFF_W4119(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120I));
DFF_save_fm DFF_W4120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121I));
DFF_save_fm DFF_W4121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122I));
DFF_save_fm DFF_W4122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100J));
DFF_save_fm DFF_W4123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101J));
DFF_save_fm DFF_W4124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102J));
DFF_save_fm DFF_W4125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110J));
DFF_save_fm DFF_W4126(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111J));
DFF_save_fm DFF_W4127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112J));
DFF_save_fm DFF_W4128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120J));
DFF_save_fm DFF_W4129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121J));
DFF_save_fm DFF_W4130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122J));
DFF_save_fm DFF_W4131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100K));
DFF_save_fm DFF_W4132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101K));
DFF_save_fm DFF_W4133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102K));
DFF_save_fm DFF_W4134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110K));
DFF_save_fm DFF_W4135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111K));
DFF_save_fm DFF_W4136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112K));
DFF_save_fm DFF_W4137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120K));
DFF_save_fm DFF_W4138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121K));
DFF_save_fm DFF_W4139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122K));
DFF_save_fm DFF_W4140(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100L));
DFF_save_fm DFF_W4141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101L));
DFF_save_fm DFF_W4142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102L));
DFF_save_fm DFF_W4143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110L));
DFF_save_fm DFF_W4144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111L));
DFF_save_fm DFF_W4145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112L));
DFF_save_fm DFF_W4146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120L));
DFF_save_fm DFF_W4147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121L));
DFF_save_fm DFF_W4148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122L));
DFF_save_fm DFF_W4149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100M));
DFF_save_fm DFF_W4150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101M));
DFF_save_fm DFF_W4151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102M));
DFF_save_fm DFF_W4152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110M));
DFF_save_fm DFF_W4153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111M));
DFF_save_fm DFF_W4154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112M));
DFF_save_fm DFF_W4155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120M));
DFF_save_fm DFF_W4156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121M));
DFF_save_fm DFF_W4157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122M));
ninexnine_unit ninexnine_unit_4512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20000)
);

ninexnine_unit ninexnine_unit_4513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21000)
);

ninexnine_unit ninexnine_unit_4514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22000)
);

ninexnine_unit ninexnine_unit_4515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23000)
);

ninexnine_unit ninexnine_unit_4516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24000)
);

ninexnine_unit ninexnine_unit_4517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25000)
);

ninexnine_unit ninexnine_unit_4518(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26000)
);

ninexnine_unit ninexnine_unit_4519(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27000)
);

ninexnine_unit ninexnine_unit_4520(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28000)
);

ninexnine_unit ninexnine_unit_4521(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29000)
);

ninexnine_unit ninexnine_unit_4522(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A000)
);

ninexnine_unit ninexnine_unit_4523(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B000)
);

ninexnine_unit ninexnine_unit_4524(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C000)
);

ninexnine_unit ninexnine_unit_4525(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D000)
);

ninexnine_unit ninexnine_unit_4526(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E000)
);

ninexnine_unit ninexnine_unit_4527(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F000)
);

ninexnine_unit ninexnine_unit_4528(
				.clk(clk),
				.rstn(rstn),
				.a0(P200G),
				.a1(P201G),
				.a2(P202G),
				.a3(P210G),
				.a4(P211G),
				.a5(P212G),
				.a6(P220G),
				.a7(P221G),
				.a8(P222G),
				.b0(W2000G),
				.b1(W2001G),
				.b2(W2002G),
				.b3(W2010G),
				.b4(W2011G),
				.b5(W2012G),
				.b6(W2020G),
				.b7(W2021G),
				.b8(W2022G),
				.c(c2G000)
);

ninexnine_unit ninexnine_unit_4529(
				.clk(clk),
				.rstn(rstn),
				.a0(P200H),
				.a1(P201H),
				.a2(P202H),
				.a3(P210H),
				.a4(P211H),
				.a5(P212H),
				.a6(P220H),
				.a7(P221H),
				.a8(P222H),
				.b0(W2000H),
				.b1(W2001H),
				.b2(W2002H),
				.b3(W2010H),
				.b4(W2011H),
				.b5(W2012H),
				.b6(W2020H),
				.b7(W2021H),
				.b8(W2022H),
				.c(c2H000)
);

ninexnine_unit ninexnine_unit_4530(
				.clk(clk),
				.rstn(rstn),
				.a0(P200I),
				.a1(P201I),
				.a2(P202I),
				.a3(P210I),
				.a4(P211I),
				.a5(P212I),
				.a6(P220I),
				.a7(P221I),
				.a8(P222I),
				.b0(W2000I),
				.b1(W2001I),
				.b2(W2002I),
				.b3(W2010I),
				.b4(W2011I),
				.b5(W2012I),
				.b6(W2020I),
				.b7(W2021I),
				.b8(W2022I),
				.c(c2I000)
);

ninexnine_unit ninexnine_unit_4531(
				.clk(clk),
				.rstn(rstn),
				.a0(P200J),
				.a1(P201J),
				.a2(P202J),
				.a3(P210J),
				.a4(P211J),
				.a5(P212J),
				.a6(P220J),
				.a7(P221J),
				.a8(P222J),
				.b0(W2000J),
				.b1(W2001J),
				.b2(W2002J),
				.b3(W2010J),
				.b4(W2011J),
				.b5(W2012J),
				.b6(W2020J),
				.b7(W2021J),
				.b8(W2022J),
				.c(c2J000)
);

ninexnine_unit ninexnine_unit_4532(
				.clk(clk),
				.rstn(rstn),
				.a0(P200K),
				.a1(P201K),
				.a2(P202K),
				.a3(P210K),
				.a4(P211K),
				.a5(P212K),
				.a6(P220K),
				.a7(P221K),
				.a8(P222K),
				.b0(W2000K),
				.b1(W2001K),
				.b2(W2002K),
				.b3(W2010K),
				.b4(W2011K),
				.b5(W2012K),
				.b6(W2020K),
				.b7(W2021K),
				.b8(W2022K),
				.c(c2K000)
);

ninexnine_unit ninexnine_unit_4533(
				.clk(clk),
				.rstn(rstn),
				.a0(P200L),
				.a1(P201L),
				.a2(P202L),
				.a3(P210L),
				.a4(P211L),
				.a5(P212L),
				.a6(P220L),
				.a7(P221L),
				.a8(P222L),
				.b0(W2000L),
				.b1(W2001L),
				.b2(W2002L),
				.b3(W2010L),
				.b4(W2011L),
				.b5(W2012L),
				.b6(W2020L),
				.b7(W2021L),
				.b8(W2022L),
				.c(c2L000)
);

ninexnine_unit ninexnine_unit_4534(
				.clk(clk),
				.rstn(rstn),
				.a0(P200M),
				.a1(P201M),
				.a2(P202M),
				.a3(P210M),
				.a4(P211M),
				.a5(P212M),
				.a6(P220M),
				.a7(P221M),
				.a8(P222M),
				.b0(W2000M),
				.b1(W2001M),
				.b2(W2002M),
				.b3(W2010M),
				.b4(W2011M),
				.b5(W2012M),
				.b6(W2020M),
				.b7(W2021M),
				.b8(W2022M),
				.c(c2M000)
);

assign C2000=c20000+c21000+c22000+c23000+c24000+c25000+c26000+c27000+c28000+c29000+c2A000+c2B000+c2C000+c2D000+c2E000+c2F000+c2G000+c2H000+c2I000+c2J000+c2K000+c2L000+c2M000;
assign A2000=(C2000>=0)?1:0;

assign P3000=A2000;

ninexnine_unit ninexnine_unit_4535(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20001)
);

ninexnine_unit ninexnine_unit_4536(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21001)
);

ninexnine_unit ninexnine_unit_4537(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22001)
);

ninexnine_unit ninexnine_unit_4538(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23001)
);

ninexnine_unit ninexnine_unit_4539(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24001)
);

ninexnine_unit ninexnine_unit_4540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25001)
);

ninexnine_unit ninexnine_unit_4541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26001)
);

ninexnine_unit ninexnine_unit_4542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27001)
);

ninexnine_unit ninexnine_unit_4543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28001)
);

ninexnine_unit ninexnine_unit_4544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29001)
);

ninexnine_unit ninexnine_unit_4545(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A001)
);

ninexnine_unit ninexnine_unit_4546(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B001)
);

ninexnine_unit ninexnine_unit_4547(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C001)
);

ninexnine_unit ninexnine_unit_4548(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D001)
);

ninexnine_unit ninexnine_unit_4549(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E001)
);

ninexnine_unit ninexnine_unit_4550(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F001)
);

ninexnine_unit ninexnine_unit_4551(
				.clk(clk),
				.rstn(rstn),
				.a0(P200G),
				.a1(P201G),
				.a2(P202G),
				.a3(P210G),
				.a4(P211G),
				.a5(P212G),
				.a6(P220G),
				.a7(P221G),
				.a8(P222G),
				.b0(W2100G),
				.b1(W2101G),
				.b2(W2102G),
				.b3(W2110G),
				.b4(W2111G),
				.b5(W2112G),
				.b6(W2120G),
				.b7(W2121G),
				.b8(W2122G),
				.c(c2G001)
);

ninexnine_unit ninexnine_unit_4552(
				.clk(clk),
				.rstn(rstn),
				.a0(P200H),
				.a1(P201H),
				.a2(P202H),
				.a3(P210H),
				.a4(P211H),
				.a5(P212H),
				.a6(P220H),
				.a7(P221H),
				.a8(P222H),
				.b0(W2100H),
				.b1(W2101H),
				.b2(W2102H),
				.b3(W2110H),
				.b4(W2111H),
				.b5(W2112H),
				.b6(W2120H),
				.b7(W2121H),
				.b8(W2122H),
				.c(c2H001)
);

ninexnine_unit ninexnine_unit_4553(
				.clk(clk),
				.rstn(rstn),
				.a0(P200I),
				.a1(P201I),
				.a2(P202I),
				.a3(P210I),
				.a4(P211I),
				.a5(P212I),
				.a6(P220I),
				.a7(P221I),
				.a8(P222I),
				.b0(W2100I),
				.b1(W2101I),
				.b2(W2102I),
				.b3(W2110I),
				.b4(W2111I),
				.b5(W2112I),
				.b6(W2120I),
				.b7(W2121I),
				.b8(W2122I),
				.c(c2I001)
);

ninexnine_unit ninexnine_unit_4554(
				.clk(clk),
				.rstn(rstn),
				.a0(P200J),
				.a1(P201J),
				.a2(P202J),
				.a3(P210J),
				.a4(P211J),
				.a5(P212J),
				.a6(P220J),
				.a7(P221J),
				.a8(P222J),
				.b0(W2100J),
				.b1(W2101J),
				.b2(W2102J),
				.b3(W2110J),
				.b4(W2111J),
				.b5(W2112J),
				.b6(W2120J),
				.b7(W2121J),
				.b8(W2122J),
				.c(c2J001)
);

ninexnine_unit ninexnine_unit_4555(
				.clk(clk),
				.rstn(rstn),
				.a0(P200K),
				.a1(P201K),
				.a2(P202K),
				.a3(P210K),
				.a4(P211K),
				.a5(P212K),
				.a6(P220K),
				.a7(P221K),
				.a8(P222K),
				.b0(W2100K),
				.b1(W2101K),
				.b2(W2102K),
				.b3(W2110K),
				.b4(W2111K),
				.b5(W2112K),
				.b6(W2120K),
				.b7(W2121K),
				.b8(W2122K),
				.c(c2K001)
);

ninexnine_unit ninexnine_unit_4556(
				.clk(clk),
				.rstn(rstn),
				.a0(P200L),
				.a1(P201L),
				.a2(P202L),
				.a3(P210L),
				.a4(P211L),
				.a5(P212L),
				.a6(P220L),
				.a7(P221L),
				.a8(P222L),
				.b0(W2100L),
				.b1(W2101L),
				.b2(W2102L),
				.b3(W2110L),
				.b4(W2111L),
				.b5(W2112L),
				.b6(W2120L),
				.b7(W2121L),
				.b8(W2122L),
				.c(c2L001)
);

ninexnine_unit ninexnine_unit_4557(
				.clk(clk),
				.rstn(rstn),
				.a0(P200M),
				.a1(P201M),
				.a2(P202M),
				.a3(P210M),
				.a4(P211M),
				.a5(P212M),
				.a6(P220M),
				.a7(P221M),
				.a8(P222M),
				.b0(W2100M),
				.b1(W2101M),
				.b2(W2102M),
				.b3(W2110M),
				.b4(W2111M),
				.b5(W2112M),
				.b6(W2120M),
				.b7(W2121M),
				.b8(W2122M),
				.c(c2M001)
);

assign C2001=c20001+c21001+c22001+c23001+c24001+c25001+c26001+c27001+c28001+c29001+c2A001+c2B001+c2C001+c2D001+c2E001+c2F001+c2G001+c2H001+c2I001+c2J001+c2K001+c2L001+c2M001;
assign A2001=(C2001>=0)?1:0;

assign P3001=A2001;

endmodule
//layer4 done, begain next layer
