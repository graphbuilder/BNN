module test_layer_all(
clk, 
rstn
);
input clk;
input rstn;

(*DONT_TOUCH="true"*) wire P0000;
(*DONT_TOUCH="true"*) wire P0010;
(*DONT_TOUCH="true"*) wire P0020;
(*DONT_TOUCH="true"*) wire P0030;
(*DONT_TOUCH="true"*) wire P0040;
(*DONT_TOUCH="true"*) wire P0050;
(*DONT_TOUCH="true"*) wire P0060;
(*DONT_TOUCH="true"*) wire P0070;
(*DONT_TOUCH="true"*) wire P0100;
(*DONT_TOUCH="true"*) wire P0110;
(*DONT_TOUCH="true"*) wire P0120;
(*DONT_TOUCH="true"*) wire P0130;
(*DONT_TOUCH="true"*) wire P0140;
(*DONT_TOUCH="true"*) wire P0150;
(*DONT_TOUCH="true"*) wire P0160;
(*DONT_TOUCH="true"*) wire P0170;
(*DONT_TOUCH="true"*) wire P0200;
(*DONT_TOUCH="true"*) wire P0210;
(*DONT_TOUCH="true"*) wire P0220;
(*DONT_TOUCH="true"*) wire P0230;
(*DONT_TOUCH="true"*) wire P0240;
(*DONT_TOUCH="true"*) wire P0250;
(*DONT_TOUCH="true"*) wire P0260;
(*DONT_TOUCH="true"*) wire P0270;
(*DONT_TOUCH="true"*) wire P0300;
(*DONT_TOUCH="true"*) wire P0310;
(*DONT_TOUCH="true"*) wire P0320;
(*DONT_TOUCH="true"*) wire P0330;
(*DONT_TOUCH="true"*) wire P0340;
(*DONT_TOUCH="true"*) wire P0350;
(*DONT_TOUCH="true"*) wire P0360;
(*DONT_TOUCH="true"*) wire P0370;
(*DONT_TOUCH="true"*) wire P0400;
(*DONT_TOUCH="true"*) wire P0410;
(*DONT_TOUCH="true"*) wire P0420;
(*DONT_TOUCH="true"*) wire P0430;
(*DONT_TOUCH="true"*) wire P0440;
(*DONT_TOUCH="true"*) wire P0450;
(*DONT_TOUCH="true"*) wire P0460;
(*DONT_TOUCH="true"*) wire P0470;
(*DONT_TOUCH="true"*) wire P0500;
(*DONT_TOUCH="true"*) wire P0510;
(*DONT_TOUCH="true"*) wire P0520;
(*DONT_TOUCH="true"*) wire P0530;
(*DONT_TOUCH="true"*) wire P0540;
(*DONT_TOUCH="true"*) wire P0550;
(*DONT_TOUCH="true"*) wire P0560;
(*DONT_TOUCH="true"*) wire P0570;
(*DONT_TOUCH="true"*) wire P0600;
(*DONT_TOUCH="true"*) wire P0610;
(*DONT_TOUCH="true"*) wire P0620;
(*DONT_TOUCH="true"*) wire P0630;
(*DONT_TOUCH="true"*) wire P0640;
(*DONT_TOUCH="true"*) wire P0650;
(*DONT_TOUCH="true"*) wire P0660;
(*DONT_TOUCH="true"*) wire P0670;
(*DONT_TOUCH="true"*) wire P0700;
(*DONT_TOUCH="true"*) wire P0710;
(*DONT_TOUCH="true"*) wire P0720;
(*DONT_TOUCH="true"*) wire P0730;
(*DONT_TOUCH="true"*) wire P0740;
(*DONT_TOUCH="true"*) wire P0750;
(*DONT_TOUCH="true"*) wire P0760;
(*DONT_TOUCH="true"*) wire P0770;
(*DONT_TOUCH="true"*) wire P0001;
(*DONT_TOUCH="true"*) wire P0011;
(*DONT_TOUCH="true"*) wire P0021;
(*DONT_TOUCH="true"*) wire P0031;
(*DONT_TOUCH="true"*) wire P0041;
(*DONT_TOUCH="true"*) wire P0051;
(*DONT_TOUCH="true"*) wire P0061;
(*DONT_TOUCH="true"*) wire P0071;
(*DONT_TOUCH="true"*) wire P0101;
(*DONT_TOUCH="true"*) wire P0111;
(*DONT_TOUCH="true"*) wire P0121;
(*DONT_TOUCH="true"*) wire P0131;
(*DONT_TOUCH="true"*) wire P0141;
(*DONT_TOUCH="true"*) wire P0151;
(*DONT_TOUCH="true"*) wire P0161;
(*DONT_TOUCH="true"*) wire P0171;
(*DONT_TOUCH="true"*) wire P0201;
(*DONT_TOUCH="true"*) wire P0211;
(*DONT_TOUCH="true"*) wire P0221;
(*DONT_TOUCH="true"*) wire P0231;
(*DONT_TOUCH="true"*) wire P0241;
(*DONT_TOUCH="true"*) wire P0251;
(*DONT_TOUCH="true"*) wire P0261;
(*DONT_TOUCH="true"*) wire P0271;
(*DONT_TOUCH="true"*) wire P0301;
(*DONT_TOUCH="true"*) wire P0311;
(*DONT_TOUCH="true"*) wire P0321;
(*DONT_TOUCH="true"*) wire P0331;
(*DONT_TOUCH="true"*) wire P0341;
(*DONT_TOUCH="true"*) wire P0351;
(*DONT_TOUCH="true"*) wire P0361;
(*DONT_TOUCH="true"*) wire P0371;
(*DONT_TOUCH="true"*) wire P0401;
(*DONT_TOUCH="true"*) wire P0411;
(*DONT_TOUCH="true"*) wire P0421;
(*DONT_TOUCH="true"*) wire P0431;
(*DONT_TOUCH="true"*) wire P0441;
(*DONT_TOUCH="true"*) wire P0451;
(*DONT_TOUCH="true"*) wire P0461;
(*DONT_TOUCH="true"*) wire P0471;
(*DONT_TOUCH="true"*) wire P0501;
(*DONT_TOUCH="true"*) wire P0511;
(*DONT_TOUCH="true"*) wire P0521;
(*DONT_TOUCH="true"*) wire P0531;
(*DONT_TOUCH="true"*) wire P0541;
(*DONT_TOUCH="true"*) wire P0551;
(*DONT_TOUCH="true"*) wire P0561;
(*DONT_TOUCH="true"*) wire P0571;
(*DONT_TOUCH="true"*) wire P0601;
(*DONT_TOUCH="true"*) wire P0611;
(*DONT_TOUCH="true"*) wire P0621;
(*DONT_TOUCH="true"*) wire P0631;
(*DONT_TOUCH="true"*) wire P0641;
(*DONT_TOUCH="true"*) wire P0651;
(*DONT_TOUCH="true"*) wire P0661;
(*DONT_TOUCH="true"*) wire P0671;
(*DONT_TOUCH="true"*) wire P0701;
(*DONT_TOUCH="true"*) wire P0711;
(*DONT_TOUCH="true"*) wire P0721;
(*DONT_TOUCH="true"*) wire P0731;
(*DONT_TOUCH="true"*) wire P0741;
(*DONT_TOUCH="true"*) wire P0751;
(*DONT_TOUCH="true"*) wire P0761;
(*DONT_TOUCH="true"*) wire P0771;
(*DONT_TOUCH="true"*) wire P0002;
(*DONT_TOUCH="true"*) wire P0012;
(*DONT_TOUCH="true"*) wire P0022;
(*DONT_TOUCH="true"*) wire P0032;
(*DONT_TOUCH="true"*) wire P0042;
(*DONT_TOUCH="true"*) wire P0052;
(*DONT_TOUCH="true"*) wire P0062;
(*DONT_TOUCH="true"*) wire P0072;
(*DONT_TOUCH="true"*) wire P0102;
(*DONT_TOUCH="true"*) wire P0112;
(*DONT_TOUCH="true"*) wire P0122;
(*DONT_TOUCH="true"*) wire P0132;
(*DONT_TOUCH="true"*) wire P0142;
(*DONT_TOUCH="true"*) wire P0152;
(*DONT_TOUCH="true"*) wire P0162;
(*DONT_TOUCH="true"*) wire P0172;
(*DONT_TOUCH="true"*) wire P0202;
(*DONT_TOUCH="true"*) wire P0212;
(*DONT_TOUCH="true"*) wire P0222;
(*DONT_TOUCH="true"*) wire P0232;
(*DONT_TOUCH="true"*) wire P0242;
(*DONT_TOUCH="true"*) wire P0252;
(*DONT_TOUCH="true"*) wire P0262;
(*DONT_TOUCH="true"*) wire P0272;
(*DONT_TOUCH="true"*) wire P0302;
(*DONT_TOUCH="true"*) wire P0312;
(*DONT_TOUCH="true"*) wire P0322;
(*DONT_TOUCH="true"*) wire P0332;
(*DONT_TOUCH="true"*) wire P0342;
(*DONT_TOUCH="true"*) wire P0352;
(*DONT_TOUCH="true"*) wire P0362;
(*DONT_TOUCH="true"*) wire P0372;
(*DONT_TOUCH="true"*) wire P0402;
(*DONT_TOUCH="true"*) wire P0412;
(*DONT_TOUCH="true"*) wire P0422;
(*DONT_TOUCH="true"*) wire P0432;
(*DONT_TOUCH="true"*) wire P0442;
(*DONT_TOUCH="true"*) wire P0452;
(*DONT_TOUCH="true"*) wire P0462;
(*DONT_TOUCH="true"*) wire P0472;
(*DONT_TOUCH="true"*) wire P0502;
(*DONT_TOUCH="true"*) wire P0512;
(*DONT_TOUCH="true"*) wire P0522;
(*DONT_TOUCH="true"*) wire P0532;
(*DONT_TOUCH="true"*) wire P0542;
(*DONT_TOUCH="true"*) wire P0552;
(*DONT_TOUCH="true"*) wire P0562;
(*DONT_TOUCH="true"*) wire P0572;
(*DONT_TOUCH="true"*) wire P0602;
(*DONT_TOUCH="true"*) wire P0612;
(*DONT_TOUCH="true"*) wire P0622;
(*DONT_TOUCH="true"*) wire P0632;
(*DONT_TOUCH="true"*) wire P0642;
(*DONT_TOUCH="true"*) wire P0652;
(*DONT_TOUCH="true"*) wire P0662;
(*DONT_TOUCH="true"*) wire P0672;
(*DONT_TOUCH="true"*) wire P0702;
(*DONT_TOUCH="true"*) wire P0712;
(*DONT_TOUCH="true"*) wire P0722;
(*DONT_TOUCH="true"*) wire P0732;
(*DONT_TOUCH="true"*) wire P0742;
(*DONT_TOUCH="true"*) wire P0752;
(*DONT_TOUCH="true"*) wire P0762;
(*DONT_TOUCH="true"*) wire P0772;
(*DONT_TOUCH="true"*) wire P1110;
(*DONT_TOUCH="true"*) wire P1120;
(*DONT_TOUCH="true"*) wire P1130;
(*DONT_TOUCH="true"*) wire P1210;
(*DONT_TOUCH="true"*) wire P1220;
(*DONT_TOUCH="true"*) wire P1230;
(*DONT_TOUCH="true"*) wire P1310;
(*DONT_TOUCH="true"*) wire P1320;
(*DONT_TOUCH="true"*) wire P1330;
(*DONT_TOUCH="true"*) wire P1111;
(*DONT_TOUCH="true"*) wire P1121;
(*DONT_TOUCH="true"*) wire P1131;
(*DONT_TOUCH="true"*) wire P1211;
(*DONT_TOUCH="true"*) wire P1221;
(*DONT_TOUCH="true"*) wire P1231;
(*DONT_TOUCH="true"*) wire P1311;
(*DONT_TOUCH="true"*) wire P1321;
(*DONT_TOUCH="true"*) wire P1331;
(*DONT_TOUCH="true"*) wire P1112;
(*DONT_TOUCH="true"*) wire P1122;
(*DONT_TOUCH="true"*) wire P1132;
(*DONT_TOUCH="true"*) wire P1212;
(*DONT_TOUCH="true"*) wire P1222;
(*DONT_TOUCH="true"*) wire P1232;
(*DONT_TOUCH="true"*) wire P1312;
(*DONT_TOUCH="true"*) wire P1322;
(*DONT_TOUCH="true"*) wire P1332;
(*DONT_TOUCH="true"*) wire P1113;
(*DONT_TOUCH="true"*) wire P1123;
(*DONT_TOUCH="true"*) wire P1133;
(*DONT_TOUCH="true"*) wire P1213;
(*DONT_TOUCH="true"*) wire P1223;
(*DONT_TOUCH="true"*) wire P1233;
(*DONT_TOUCH="true"*) wire P1313;
(*DONT_TOUCH="true"*) wire P1323;
(*DONT_TOUCH="true"*) wire P1333;
(*DONT_TOUCH="true"*) wire W00000,W00010,W00020,W00100,W00110,W00120,W00200,W00210,W00220;
(*DONT_TOUCH="true"*) wire W00001,W00011,W00021,W00101,W00111,W00121,W00201,W00211,W00221;
(*DONT_TOUCH="true"*) wire W00002,W00012,W00022,W00102,W00112,W00122,W00202,W00212,W00222;
(*DONT_TOUCH="true"*) wire W01000,W01010,W01020,W01100,W01110,W01120,W01200,W01210,W01220;
(*DONT_TOUCH="true"*) wire W01001,W01011,W01021,W01101,W01111,W01121,W01201,W01211,W01221;
(*DONT_TOUCH="true"*) wire W01002,W01012,W01022,W01102,W01112,W01122,W01202,W01212,W01222;
(*DONT_TOUCH="true"*) wire W02000,W02010,W02020,W02100,W02110,W02120,W02200,W02210,W02220;
(*DONT_TOUCH="true"*) wire W02001,W02011,W02021,W02101,W02111,W02121,W02201,W02211,W02221;
(*DONT_TOUCH="true"*) wire W02002,W02012,W02022,W02102,W02112,W02122,W02202,W02212,W02222;
(*DONT_TOUCH="true"*) wire W03000,W03010,W03020,W03100,W03110,W03120,W03200,W03210,W03220;
(*DONT_TOUCH="true"*) wire W03001,W03011,W03021,W03101,W03111,W03121,W03201,W03211,W03221;
(*DONT_TOUCH="true"*) wire W03002,W03012,W03022,W03102,W03112,W03122,W03202,W03212,W03222;
(*DONT_TOUCH="true"*) wire signed [4:0] c00000,c01000,c02000;
(*DONT_TOUCH="true"*) wire signed [4:0] c00010,c01010,c02010;
(*DONT_TOUCH="true"*) wire signed [4:0] c00020,c01020,c02020;
(*DONT_TOUCH="true"*) wire signed [4:0] c00030,c01030,c02030;
(*DONT_TOUCH="true"*) wire signed [4:0] c00040,c01040,c02040;
(*DONT_TOUCH="true"*) wire signed [4:0] c00050,c01050,c02050;
(*DONT_TOUCH="true"*) wire signed [4:0] c00100,c01100,c02100;
(*DONT_TOUCH="true"*) wire signed [4:0] c00110,c01110,c02110;
(*DONT_TOUCH="true"*) wire signed [4:0] c00120,c01120,c02120;
(*DONT_TOUCH="true"*) wire signed [4:0] c00130,c01130,c02130;
(*DONT_TOUCH="true"*) wire signed [4:0] c00140,c01140,c02140;
(*DONT_TOUCH="true"*) wire signed [4:0] c00150,c01150,c02150;
(*DONT_TOUCH="true"*) wire signed [4:0] c00200,c01200,c02200;
(*DONT_TOUCH="true"*) wire signed [4:0] c00210,c01210,c02210;
(*DONT_TOUCH="true"*) wire signed [4:0] c00220,c01220,c02220;
(*DONT_TOUCH="true"*) wire signed [4:0] c00230,c01230,c02230;
(*DONT_TOUCH="true"*) wire signed [4:0] c00240,c01240,c02240;
(*DONT_TOUCH="true"*) wire signed [4:0] c00250,c01250,c02250;
(*DONT_TOUCH="true"*) wire signed [4:0] c00300,c01300,c02300;
(*DONT_TOUCH="true"*) wire signed [4:0] c00310,c01310,c02310;
(*DONT_TOUCH="true"*) wire signed [4:0] c00320,c01320,c02320;
(*DONT_TOUCH="true"*) wire signed [4:0] c00330,c01330,c02330;
(*DONT_TOUCH="true"*) wire signed [4:0] c00340,c01340,c02340;
(*DONT_TOUCH="true"*) wire signed [4:0] c00350,c01350,c02350;
(*DONT_TOUCH="true"*) wire signed [4:0] c00400,c01400,c02400;
(*DONT_TOUCH="true"*) wire signed [4:0] c00410,c01410,c02410;
(*DONT_TOUCH="true"*) wire signed [4:0] c00420,c01420,c02420;
(*DONT_TOUCH="true"*) wire signed [4:0] c00430,c01430,c02430;
(*DONT_TOUCH="true"*) wire signed [4:0] c00440,c01440,c02440;
(*DONT_TOUCH="true"*) wire signed [4:0] c00450,c01450,c02450;
(*DONT_TOUCH="true"*) wire signed [4:0] c00500,c01500,c02500;
(*DONT_TOUCH="true"*) wire signed [4:0] c00510,c01510,c02510;
(*DONT_TOUCH="true"*) wire signed [4:0] c00520,c01520,c02520;
(*DONT_TOUCH="true"*) wire signed [4:0] c00530,c01530,c02530;
(*DONT_TOUCH="true"*) wire signed [4:0] c00540,c01540,c02540;
(*DONT_TOUCH="true"*) wire signed [4:0] c00550,c01550,c02550;
(*DONT_TOUCH="true"*) wire signed [4:0] c00001,c01001,c02001;
(*DONT_TOUCH="true"*) wire signed [4:0] c00011,c01011,c02011;
(*DONT_TOUCH="true"*) wire signed [4:0] c00021,c01021,c02021;
(*DONT_TOUCH="true"*) wire signed [4:0] c00031,c01031,c02031;
(*DONT_TOUCH="true"*) wire signed [4:0] c00041,c01041,c02041;
(*DONT_TOUCH="true"*) wire signed [4:0] c00051,c01051,c02051;
(*DONT_TOUCH="true"*) wire signed [4:0] c00101,c01101,c02101;
(*DONT_TOUCH="true"*) wire signed [4:0] c00111,c01111,c02111;
(*DONT_TOUCH="true"*) wire signed [4:0] c00121,c01121,c02121;
(*DONT_TOUCH="true"*) wire signed [4:0] c00131,c01131,c02131;
(*DONT_TOUCH="true"*) wire signed [4:0] c00141,c01141,c02141;
(*DONT_TOUCH="true"*) wire signed [4:0] c00151,c01151,c02151;
(*DONT_TOUCH="true"*) wire signed [4:0] c00201,c01201,c02201;
(*DONT_TOUCH="true"*) wire signed [4:0] c00211,c01211,c02211;
(*DONT_TOUCH="true"*) wire signed [4:0] c00221,c01221,c02221;
(*DONT_TOUCH="true"*) wire signed [4:0] c00231,c01231,c02231;
(*DONT_TOUCH="true"*) wire signed [4:0] c00241,c01241,c02241;
(*DONT_TOUCH="true"*) wire signed [4:0] c00251,c01251,c02251;
(*DONT_TOUCH="true"*) wire signed [4:0] c00301,c01301,c02301;
(*DONT_TOUCH="true"*) wire signed [4:0] c00311,c01311,c02311;
(*DONT_TOUCH="true"*) wire signed [4:0] c00321,c01321,c02321;
(*DONT_TOUCH="true"*) wire signed [4:0] c00331,c01331,c02331;
(*DONT_TOUCH="true"*) wire signed [4:0] c00341,c01341,c02341;
(*DONT_TOUCH="true"*) wire signed [4:0] c00351,c01351,c02351;
(*DONT_TOUCH="true"*) wire signed [4:0] c00401,c01401,c02401;
(*DONT_TOUCH="true"*) wire signed [4:0] c00411,c01411,c02411;
(*DONT_TOUCH="true"*) wire signed [4:0] c00421,c01421,c02421;
(*DONT_TOUCH="true"*) wire signed [4:0] c00431,c01431,c02431;
(*DONT_TOUCH="true"*) wire signed [4:0] c00441,c01441,c02441;
(*DONT_TOUCH="true"*) wire signed [4:0] c00451,c01451,c02451;
(*DONT_TOUCH="true"*) wire signed [4:0] c00501,c01501,c02501;
(*DONT_TOUCH="true"*) wire signed [4:0] c00511,c01511,c02511;
(*DONT_TOUCH="true"*) wire signed [4:0] c00521,c01521,c02521;
(*DONT_TOUCH="true"*) wire signed [4:0] c00531,c01531,c02531;
(*DONT_TOUCH="true"*) wire signed [4:0] c00541,c01541,c02541;
(*DONT_TOUCH="true"*) wire signed [4:0] c00551,c01551,c02551;
(*DONT_TOUCH="true"*) wire signed [4:0] c00002,c01002,c02002;
(*DONT_TOUCH="true"*) wire signed [4:0] c00012,c01012,c02012;
(*DONT_TOUCH="true"*) wire signed [4:0] c00022,c01022,c02022;
(*DONT_TOUCH="true"*) wire signed [4:0] c00032,c01032,c02032;
(*DONT_TOUCH="true"*) wire signed [4:0] c00042,c01042,c02042;
(*DONT_TOUCH="true"*) wire signed [4:0] c00052,c01052,c02052;
(*DONT_TOUCH="true"*) wire signed [4:0] c00102,c01102,c02102;
(*DONT_TOUCH="true"*) wire signed [4:0] c00112,c01112,c02112;
(*DONT_TOUCH="true"*) wire signed [4:0] c00122,c01122,c02122;
(*DONT_TOUCH="true"*) wire signed [4:0] c00132,c01132,c02132;
(*DONT_TOUCH="true"*) wire signed [4:0] c00142,c01142,c02142;
(*DONT_TOUCH="true"*) wire signed [4:0] c00152,c01152,c02152;
(*DONT_TOUCH="true"*) wire signed [4:0] c00202,c01202,c02202;
(*DONT_TOUCH="true"*) wire signed [4:0] c00212,c01212,c02212;
(*DONT_TOUCH="true"*) wire signed [4:0] c00222,c01222,c02222;
(*DONT_TOUCH="true"*) wire signed [4:0] c00232,c01232,c02232;
(*DONT_TOUCH="true"*) wire signed [4:0] c00242,c01242,c02242;
(*DONT_TOUCH="true"*) wire signed [4:0] c00252,c01252,c02252;
(*DONT_TOUCH="true"*) wire signed [4:0] c00302,c01302,c02302;
(*DONT_TOUCH="true"*) wire signed [4:0] c00312,c01312,c02312;
(*DONT_TOUCH="true"*) wire signed [4:0] c00322,c01322,c02322;
(*DONT_TOUCH="true"*) wire signed [4:0] c00332,c01332,c02332;
(*DONT_TOUCH="true"*) wire signed [4:0] c00342,c01342,c02342;
(*DONT_TOUCH="true"*) wire signed [4:0] c00352,c01352,c02352;
(*DONT_TOUCH="true"*) wire signed [4:0] c00402,c01402,c02402;
(*DONT_TOUCH="true"*) wire signed [4:0] c00412,c01412,c02412;
(*DONT_TOUCH="true"*) wire signed [4:0] c00422,c01422,c02422;
(*DONT_TOUCH="true"*) wire signed [4:0] c00432,c01432,c02432;
(*DONT_TOUCH="true"*) wire signed [4:0] c00442,c01442,c02442;
(*DONT_TOUCH="true"*) wire signed [4:0] c00452,c01452,c02452;
(*DONT_TOUCH="true"*) wire signed [4:0] c00502,c01502,c02502;
(*DONT_TOUCH="true"*) wire signed [4:0] c00512,c01512,c02512;
(*DONT_TOUCH="true"*) wire signed [4:0] c00522,c01522,c02522;
(*DONT_TOUCH="true"*) wire signed [4:0] c00532,c01532,c02532;
(*DONT_TOUCH="true"*) wire signed [4:0] c00542,c01542,c02542;
(*DONT_TOUCH="true"*) wire signed [4:0] c00552,c01552,c02552;
(*DONT_TOUCH="true"*) wire signed [4:0] c00003,c01003,c02003;
(*DONT_TOUCH="true"*) wire signed [4:0] c00013,c01013,c02013;
(*DONT_TOUCH="true"*) wire signed [4:0] c00023,c01023,c02023;
(*DONT_TOUCH="true"*) wire signed [4:0] c00033,c01033,c02033;
(*DONT_TOUCH="true"*) wire signed [4:0] c00043,c01043,c02043;
(*DONT_TOUCH="true"*) wire signed [4:0] c00053,c01053,c02053;
(*DONT_TOUCH="true"*) wire signed [4:0] c00103,c01103,c02103;
(*DONT_TOUCH="true"*) wire signed [4:0] c00113,c01113,c02113;
(*DONT_TOUCH="true"*) wire signed [4:0] c00123,c01123,c02123;
(*DONT_TOUCH="true"*) wire signed [4:0] c00133,c01133,c02133;
(*DONT_TOUCH="true"*) wire signed [4:0] c00143,c01143,c02143;
(*DONT_TOUCH="true"*) wire signed [4:0] c00153,c01153,c02153;
(*DONT_TOUCH="true"*) wire signed [4:0] c00203,c01203,c02203;
(*DONT_TOUCH="true"*) wire signed [4:0] c00213,c01213,c02213;
(*DONT_TOUCH="true"*) wire signed [4:0] c00223,c01223,c02223;
(*DONT_TOUCH="true"*) wire signed [4:0] c00233,c01233,c02233;
(*DONT_TOUCH="true"*) wire signed [4:0] c00243,c01243,c02243;
(*DONT_TOUCH="true"*) wire signed [4:0] c00253,c01253,c02253;
(*DONT_TOUCH="true"*) wire signed [4:0] c00303,c01303,c02303;
(*DONT_TOUCH="true"*) wire signed [4:0] c00313,c01313,c02313;
(*DONT_TOUCH="true"*) wire signed [4:0] c00323,c01323,c02323;
(*DONT_TOUCH="true"*) wire signed [4:0] c00333,c01333,c02333;
(*DONT_TOUCH="true"*) wire signed [4:0] c00343,c01343,c02343;
(*DONT_TOUCH="true"*) wire signed [4:0] c00353,c01353,c02353;
(*DONT_TOUCH="true"*) wire signed [4:0] c00403,c01403,c02403;
(*DONT_TOUCH="true"*) wire signed [4:0] c00413,c01413,c02413;
(*DONT_TOUCH="true"*) wire signed [4:0] c00423,c01423,c02423;
(*DONT_TOUCH="true"*) wire signed [4:0] c00433,c01433,c02433;
(*DONT_TOUCH="true"*) wire signed [4:0] c00443,c01443,c02443;
(*DONT_TOUCH="true"*) wire signed [4:0] c00453,c01453,c02453;
(*DONT_TOUCH="true"*) wire signed [4:0] c00503,c01503,c02503;
(*DONT_TOUCH="true"*) wire signed [4:0] c00513,c01513,c02513;
(*DONT_TOUCH="true"*) wire signed [4:0] c00523,c01523,c02523;
(*DONT_TOUCH="true"*) wire signed [4:0] c00533,c01533,c02533;
(*DONT_TOUCH="true"*) wire signed [4:0] c00543,c01543,c02543;
(*DONT_TOUCH="true"*) wire signed [4:0] c00553,c01553,c02553;
(*DONT_TOUCH="true"*) wire signed [6:0] C0000;
(*DONT_TOUCH="true"*) wire A0000;
(*DONT_TOUCH="true"*) wire signed [6:0] C0010;
(*DONT_TOUCH="true"*) wire A0010;
(*DONT_TOUCH="true"*) wire signed [6:0] C0020;
(*DONT_TOUCH="true"*) wire A0020;
(*DONT_TOUCH="true"*) wire signed [6:0] C0030;
(*DONT_TOUCH="true"*) wire A0030;
(*DONT_TOUCH="true"*) wire signed [6:0] C0040;
(*DONT_TOUCH="true"*) wire A0040;
(*DONT_TOUCH="true"*) wire signed [6:0] C0050;
(*DONT_TOUCH="true"*) wire A0050;
(*DONT_TOUCH="true"*) wire signed [6:0] C0100;
(*DONT_TOUCH="true"*) wire A0100;
(*DONT_TOUCH="true"*) wire signed [6:0] C0110;
(*DONT_TOUCH="true"*) wire A0110;
(*DONT_TOUCH="true"*) wire signed [6:0] C0120;
(*DONT_TOUCH="true"*) wire A0120;
(*DONT_TOUCH="true"*) wire signed [6:0] C0130;
(*DONT_TOUCH="true"*) wire A0130;
(*DONT_TOUCH="true"*) wire signed [6:0] C0140;
(*DONT_TOUCH="true"*) wire A0140;
(*DONT_TOUCH="true"*) wire signed [6:0] C0150;
(*DONT_TOUCH="true"*) wire A0150;
(*DONT_TOUCH="true"*) wire signed [6:0] C0200;
(*DONT_TOUCH="true"*) wire A0200;
(*DONT_TOUCH="true"*) wire signed [6:0] C0210;
(*DONT_TOUCH="true"*) wire A0210;
(*DONT_TOUCH="true"*) wire signed [6:0] C0220;
(*DONT_TOUCH="true"*) wire A0220;
(*DONT_TOUCH="true"*) wire signed [6:0] C0230;
(*DONT_TOUCH="true"*) wire A0230;
(*DONT_TOUCH="true"*) wire signed [6:0] C0240;
(*DONT_TOUCH="true"*) wire A0240;
(*DONT_TOUCH="true"*) wire signed [6:0] C0250;
(*DONT_TOUCH="true"*) wire A0250;
(*DONT_TOUCH="true"*) wire signed [6:0] C0300;
(*DONT_TOUCH="true"*) wire A0300;
(*DONT_TOUCH="true"*) wire signed [6:0] C0310;
(*DONT_TOUCH="true"*) wire A0310;
(*DONT_TOUCH="true"*) wire signed [6:0] C0320;
(*DONT_TOUCH="true"*) wire A0320;
(*DONT_TOUCH="true"*) wire signed [6:0] C0330;
(*DONT_TOUCH="true"*) wire A0330;
(*DONT_TOUCH="true"*) wire signed [6:0] C0340;
(*DONT_TOUCH="true"*) wire A0340;
(*DONT_TOUCH="true"*) wire signed [6:0] C0350;
(*DONT_TOUCH="true"*) wire A0350;
(*DONT_TOUCH="true"*) wire signed [6:0] C0400;
(*DONT_TOUCH="true"*) wire A0400;
(*DONT_TOUCH="true"*) wire signed [6:0] C0410;
(*DONT_TOUCH="true"*) wire A0410;
(*DONT_TOUCH="true"*) wire signed [6:0] C0420;
(*DONT_TOUCH="true"*) wire A0420;
(*DONT_TOUCH="true"*) wire signed [6:0] C0430;
(*DONT_TOUCH="true"*) wire A0430;
(*DONT_TOUCH="true"*) wire signed [6:0] C0440;
(*DONT_TOUCH="true"*) wire A0440;
(*DONT_TOUCH="true"*) wire signed [6:0] C0450;
(*DONT_TOUCH="true"*) wire A0450;
(*DONT_TOUCH="true"*) wire signed [6:0] C0500;
(*DONT_TOUCH="true"*) wire A0500;
(*DONT_TOUCH="true"*) wire signed [6:0] C0510;
(*DONT_TOUCH="true"*) wire A0510;
(*DONT_TOUCH="true"*) wire signed [6:0] C0520;
(*DONT_TOUCH="true"*) wire A0520;
(*DONT_TOUCH="true"*) wire signed [6:0] C0530;
(*DONT_TOUCH="true"*) wire A0530;
(*DONT_TOUCH="true"*) wire signed [6:0] C0540;
(*DONT_TOUCH="true"*) wire A0540;
(*DONT_TOUCH="true"*) wire signed [6:0] C0550;
(*DONT_TOUCH="true"*) wire A0550;
(*DONT_TOUCH="true"*) wire signed [6:0] C0001;
(*DONT_TOUCH="true"*) wire A0001;
(*DONT_TOUCH="true"*) wire signed [6:0] C0011;
(*DONT_TOUCH="true"*) wire A0011;
(*DONT_TOUCH="true"*) wire signed [6:0] C0021;
(*DONT_TOUCH="true"*) wire A0021;
(*DONT_TOUCH="true"*) wire signed [6:0] C0031;
(*DONT_TOUCH="true"*) wire A0031;
(*DONT_TOUCH="true"*) wire signed [6:0] C0041;
(*DONT_TOUCH="true"*) wire A0041;
(*DONT_TOUCH="true"*) wire signed [6:0] C0051;
(*DONT_TOUCH="true"*) wire A0051;
(*DONT_TOUCH="true"*) wire signed [6:0] C0101;
(*DONT_TOUCH="true"*) wire A0101;
(*DONT_TOUCH="true"*) wire signed [6:0] C0111;
(*DONT_TOUCH="true"*) wire A0111;
(*DONT_TOUCH="true"*) wire signed [6:0] C0121;
(*DONT_TOUCH="true"*) wire A0121;
(*DONT_TOUCH="true"*) wire signed [6:0] C0131;
(*DONT_TOUCH="true"*) wire A0131;
(*DONT_TOUCH="true"*) wire signed [6:0] C0141;
(*DONT_TOUCH="true"*) wire A0141;
(*DONT_TOUCH="true"*) wire signed [6:0] C0151;
(*DONT_TOUCH="true"*) wire A0151;
(*DONT_TOUCH="true"*) wire signed [6:0] C0201;
(*DONT_TOUCH="true"*) wire A0201;
(*DONT_TOUCH="true"*) wire signed [6:0] C0211;
(*DONT_TOUCH="true"*) wire A0211;
(*DONT_TOUCH="true"*) wire signed [6:0] C0221;
(*DONT_TOUCH="true"*) wire A0221;
(*DONT_TOUCH="true"*) wire signed [6:0] C0231;
(*DONT_TOUCH="true"*) wire A0231;
(*DONT_TOUCH="true"*) wire signed [6:0] C0241;
(*DONT_TOUCH="true"*) wire A0241;
(*DONT_TOUCH="true"*) wire signed [6:0] C0251;
(*DONT_TOUCH="true"*) wire A0251;
(*DONT_TOUCH="true"*) wire signed [6:0] C0301;
(*DONT_TOUCH="true"*) wire A0301;
(*DONT_TOUCH="true"*) wire signed [6:0] C0311;
(*DONT_TOUCH="true"*) wire A0311;
(*DONT_TOUCH="true"*) wire signed [6:0] C0321;
(*DONT_TOUCH="true"*) wire A0321;
(*DONT_TOUCH="true"*) wire signed [6:0] C0331;
(*DONT_TOUCH="true"*) wire A0331;
(*DONT_TOUCH="true"*) wire signed [6:0] C0341;
(*DONT_TOUCH="true"*) wire A0341;
(*DONT_TOUCH="true"*) wire signed [6:0] C0351;
(*DONT_TOUCH="true"*) wire A0351;
(*DONT_TOUCH="true"*) wire signed [6:0] C0401;
(*DONT_TOUCH="true"*) wire A0401;
(*DONT_TOUCH="true"*) wire signed [6:0] C0411;
(*DONT_TOUCH="true"*) wire A0411;
(*DONT_TOUCH="true"*) wire signed [6:0] C0421;
(*DONT_TOUCH="true"*) wire A0421;
(*DONT_TOUCH="true"*) wire signed [6:0] C0431;
(*DONT_TOUCH="true"*) wire A0431;
(*DONT_TOUCH="true"*) wire signed [6:0] C0441;
(*DONT_TOUCH="true"*) wire A0441;
(*DONT_TOUCH="true"*) wire signed [6:0] C0451;
(*DONT_TOUCH="true"*) wire A0451;
(*DONT_TOUCH="true"*) wire signed [6:0] C0501;
(*DONT_TOUCH="true"*) wire A0501;
(*DONT_TOUCH="true"*) wire signed [6:0] C0511;
(*DONT_TOUCH="true"*) wire A0511;
(*DONT_TOUCH="true"*) wire signed [6:0] C0521;
(*DONT_TOUCH="true"*) wire A0521;
(*DONT_TOUCH="true"*) wire signed [6:0] C0531;
(*DONT_TOUCH="true"*) wire A0531;
(*DONT_TOUCH="true"*) wire signed [6:0] C0541;
(*DONT_TOUCH="true"*) wire A0541;
(*DONT_TOUCH="true"*) wire signed [6:0] C0551;
(*DONT_TOUCH="true"*) wire A0551;
(*DONT_TOUCH="true"*) wire signed [6:0] C0002;
(*DONT_TOUCH="true"*) wire A0002;
(*DONT_TOUCH="true"*) wire signed [6:0] C0012;
(*DONT_TOUCH="true"*) wire A0012;
(*DONT_TOUCH="true"*) wire signed [6:0] C0022;
(*DONT_TOUCH="true"*) wire A0022;
(*DONT_TOUCH="true"*) wire signed [6:0] C0032;
(*DONT_TOUCH="true"*) wire A0032;
(*DONT_TOUCH="true"*) wire signed [6:0] C0042;
(*DONT_TOUCH="true"*) wire A0042;
(*DONT_TOUCH="true"*) wire signed [6:0] C0052;
(*DONT_TOUCH="true"*) wire A0052;
(*DONT_TOUCH="true"*) wire signed [6:0] C0102;
(*DONT_TOUCH="true"*) wire A0102;
(*DONT_TOUCH="true"*) wire signed [6:0] C0112;
(*DONT_TOUCH="true"*) wire A0112;
(*DONT_TOUCH="true"*) wire signed [6:0] C0122;
(*DONT_TOUCH="true"*) wire A0122;
(*DONT_TOUCH="true"*) wire signed [6:0] C0132;
(*DONT_TOUCH="true"*) wire A0132;
(*DONT_TOUCH="true"*) wire signed [6:0] C0142;
(*DONT_TOUCH="true"*) wire A0142;
(*DONT_TOUCH="true"*) wire signed [6:0] C0152;
(*DONT_TOUCH="true"*) wire A0152;
(*DONT_TOUCH="true"*) wire signed [6:0] C0202;
(*DONT_TOUCH="true"*) wire A0202;
(*DONT_TOUCH="true"*) wire signed [6:0] C0212;
(*DONT_TOUCH="true"*) wire A0212;
(*DONT_TOUCH="true"*) wire signed [6:0] C0222;
(*DONT_TOUCH="true"*) wire A0222;
(*DONT_TOUCH="true"*) wire signed [6:0] C0232;
(*DONT_TOUCH="true"*) wire A0232;
(*DONT_TOUCH="true"*) wire signed [6:0] C0242;
(*DONT_TOUCH="true"*) wire A0242;
(*DONT_TOUCH="true"*) wire signed [6:0] C0252;
(*DONT_TOUCH="true"*) wire A0252;
(*DONT_TOUCH="true"*) wire signed [6:0] C0302;
(*DONT_TOUCH="true"*) wire A0302;
(*DONT_TOUCH="true"*) wire signed [6:0] C0312;
(*DONT_TOUCH="true"*) wire A0312;
(*DONT_TOUCH="true"*) wire signed [6:0] C0322;
(*DONT_TOUCH="true"*) wire A0322;
(*DONT_TOUCH="true"*) wire signed [6:0] C0332;
(*DONT_TOUCH="true"*) wire A0332;
(*DONT_TOUCH="true"*) wire signed [6:0] C0342;
(*DONT_TOUCH="true"*) wire A0342;
(*DONT_TOUCH="true"*) wire signed [6:0] C0352;
(*DONT_TOUCH="true"*) wire A0352;
(*DONT_TOUCH="true"*) wire signed [6:0] C0402;
(*DONT_TOUCH="true"*) wire A0402;
(*DONT_TOUCH="true"*) wire signed [6:0] C0412;
(*DONT_TOUCH="true"*) wire A0412;
(*DONT_TOUCH="true"*) wire signed [6:0] C0422;
(*DONT_TOUCH="true"*) wire A0422;
(*DONT_TOUCH="true"*) wire signed [6:0] C0432;
(*DONT_TOUCH="true"*) wire A0432;
(*DONT_TOUCH="true"*) wire signed [6:0] C0442;
(*DONT_TOUCH="true"*) wire A0442;
(*DONT_TOUCH="true"*) wire signed [6:0] C0452;
(*DONT_TOUCH="true"*) wire A0452;
(*DONT_TOUCH="true"*) wire signed [6:0] C0502;
(*DONT_TOUCH="true"*) wire A0502;
(*DONT_TOUCH="true"*) wire signed [6:0] C0512;
(*DONT_TOUCH="true"*) wire A0512;
(*DONT_TOUCH="true"*) wire signed [6:0] C0522;
(*DONT_TOUCH="true"*) wire A0522;
(*DONT_TOUCH="true"*) wire signed [6:0] C0532;
(*DONT_TOUCH="true"*) wire A0532;
(*DONT_TOUCH="true"*) wire signed [6:0] C0542;
(*DONT_TOUCH="true"*) wire A0542;
(*DONT_TOUCH="true"*) wire signed [6:0] C0552;
(*DONT_TOUCH="true"*) wire A0552;
(*DONT_TOUCH="true"*) wire signed [6:0] C0003;
(*DONT_TOUCH="true"*) wire A0003;
(*DONT_TOUCH="true"*) wire signed [6:0] C0013;
(*DONT_TOUCH="true"*) wire A0013;
(*DONT_TOUCH="true"*) wire signed [6:0] C0023;
(*DONT_TOUCH="true"*) wire A0023;
(*DONT_TOUCH="true"*) wire signed [6:0] C0033;
(*DONT_TOUCH="true"*) wire A0033;
(*DONT_TOUCH="true"*) wire signed [6:0] C0043;
(*DONT_TOUCH="true"*) wire A0043;
(*DONT_TOUCH="true"*) wire signed [6:0] C0053;
(*DONT_TOUCH="true"*) wire A0053;
(*DONT_TOUCH="true"*) wire signed [6:0] C0103;
(*DONT_TOUCH="true"*) wire A0103;
(*DONT_TOUCH="true"*) wire signed [6:0] C0113;
(*DONT_TOUCH="true"*) wire A0113;
(*DONT_TOUCH="true"*) wire signed [6:0] C0123;
(*DONT_TOUCH="true"*) wire A0123;
(*DONT_TOUCH="true"*) wire signed [6:0] C0133;
(*DONT_TOUCH="true"*) wire A0133;
(*DONT_TOUCH="true"*) wire signed [6:0] C0143;
(*DONT_TOUCH="true"*) wire A0143;
(*DONT_TOUCH="true"*) wire signed [6:0] C0153;
(*DONT_TOUCH="true"*) wire A0153;
(*DONT_TOUCH="true"*) wire signed [6:0] C0203;
(*DONT_TOUCH="true"*) wire A0203;
(*DONT_TOUCH="true"*) wire signed [6:0] C0213;
(*DONT_TOUCH="true"*) wire A0213;
(*DONT_TOUCH="true"*) wire signed [6:0] C0223;
(*DONT_TOUCH="true"*) wire A0223;
(*DONT_TOUCH="true"*) wire signed [6:0] C0233;
(*DONT_TOUCH="true"*) wire A0233;
(*DONT_TOUCH="true"*) wire signed [6:0] C0243;
(*DONT_TOUCH="true"*) wire A0243;
(*DONT_TOUCH="true"*) wire signed [6:0] C0253;
(*DONT_TOUCH="true"*) wire A0253;
(*DONT_TOUCH="true"*) wire signed [6:0] C0303;
(*DONT_TOUCH="true"*) wire A0303;
(*DONT_TOUCH="true"*) wire signed [6:0] C0313;
(*DONT_TOUCH="true"*) wire A0313;
(*DONT_TOUCH="true"*) wire signed [6:0] C0323;
(*DONT_TOUCH="true"*) wire A0323;
(*DONT_TOUCH="true"*) wire signed [6:0] C0333;
(*DONT_TOUCH="true"*) wire A0333;
(*DONT_TOUCH="true"*) wire signed [6:0] C0343;
(*DONT_TOUCH="true"*) wire A0343;
(*DONT_TOUCH="true"*) wire signed [6:0] C0353;
(*DONT_TOUCH="true"*) wire A0353;
(*DONT_TOUCH="true"*) wire signed [6:0] C0403;
(*DONT_TOUCH="true"*) wire A0403;
(*DONT_TOUCH="true"*) wire signed [6:0] C0413;
(*DONT_TOUCH="true"*) wire A0413;
(*DONT_TOUCH="true"*) wire signed [6:0] C0423;
(*DONT_TOUCH="true"*) wire A0423;
(*DONT_TOUCH="true"*) wire signed [6:0] C0433;
(*DONT_TOUCH="true"*) wire A0433;
(*DONT_TOUCH="true"*) wire signed [6:0] C0443;
(*DONT_TOUCH="true"*) wire A0443;
(*DONT_TOUCH="true"*) wire signed [6:0] C0453;
(*DONT_TOUCH="true"*) wire A0453;
(*DONT_TOUCH="true"*) wire signed [6:0] C0503;
(*DONT_TOUCH="true"*) wire A0503;
(*DONT_TOUCH="true"*) wire signed [6:0] C0513;
(*DONT_TOUCH="true"*) wire A0513;
(*DONT_TOUCH="true"*) wire signed [6:0] C0523;
(*DONT_TOUCH="true"*) wire A0523;
(*DONT_TOUCH="true"*) wire signed [6:0] C0533;
(*DONT_TOUCH="true"*) wire A0533;
(*DONT_TOUCH="true"*) wire signed [6:0] C0543;
(*DONT_TOUCH="true"*) wire A0543;
(*DONT_TOUCH="true"*) wire signed [6:0] C0553;
(*DONT_TOUCH="true"*) wire A0553;
DFF_save_fm DFF_P0(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0000));
DFF_save_fm DFF_P1(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0010));
DFF_save_fm DFF_P2(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0020));
DFF_save_fm DFF_P3(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0030));
DFF_save_fm DFF_P4(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0040));
DFF_save_fm DFF_P5(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0050));
DFF_save_fm DFF_P6(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0060));
DFF_save_fm DFF_P7(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0070));
DFF_save_fm DFF_P8(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0100));
DFF_save_fm DFF_P9(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0110));
DFF_save_fm DFF_P10(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0120));
DFF_save_fm DFF_P11(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0130));
DFF_save_fm DFF_P12(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0140));
DFF_save_fm DFF_P13(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0150));
DFF_save_fm DFF_P14(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0160));
DFF_save_fm DFF_P15(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0170));
DFF_save_fm DFF_P16(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0200));
DFF_save_fm DFF_P17(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0210));
DFF_save_fm DFF_P18(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0220));
DFF_save_fm DFF_P19(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0230));
DFF_save_fm DFF_P20(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0240));
DFF_save_fm DFF_P21(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0250));
DFF_save_fm DFF_P22(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0260));
DFF_save_fm DFF_P23(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0270));
DFF_save_fm DFF_P24(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0300));
DFF_save_fm DFF_P25(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0310));
DFF_save_fm DFF_P26(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0320));
DFF_save_fm DFF_P27(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0330));
DFF_save_fm DFF_P28(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0340));
DFF_save_fm DFF_P29(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0350));
DFF_save_fm DFF_P30(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0360));
DFF_save_fm DFF_P31(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0370));
DFF_save_fm DFF_P32(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0400));
DFF_save_fm DFF_P33(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0410));
DFF_save_fm DFF_P34(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0420));
DFF_save_fm DFF_P35(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0430));
DFF_save_fm DFF_P36(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0440));
DFF_save_fm DFF_P37(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0450));
DFF_save_fm DFF_P38(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0460));
DFF_save_fm DFF_P39(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0470));
DFF_save_fm DFF_P40(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0500));
DFF_save_fm DFF_P41(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0510));
DFF_save_fm DFF_P42(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0520));
DFF_save_fm DFF_P43(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0530));
DFF_save_fm DFF_P44(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0540));
DFF_save_fm DFF_P45(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0550));
DFF_save_fm DFF_P46(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0560));
DFF_save_fm DFF_P47(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0570));
DFF_save_fm DFF_P48(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0600));
DFF_save_fm DFF_P49(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0610));
DFF_save_fm DFF_P50(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0620));
DFF_save_fm DFF_P51(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0630));
DFF_save_fm DFF_P52(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0640));
DFF_save_fm DFF_P53(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0650));
DFF_save_fm DFF_P54(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0660));
DFF_save_fm DFF_P55(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0670));
DFF_save_fm DFF_P56(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0700));
DFF_save_fm DFF_P57(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0710));
DFF_save_fm DFF_P58(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0720));
DFF_save_fm DFF_P59(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0730));
DFF_save_fm DFF_P60(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0740));
DFF_save_fm DFF_P61(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0750));
DFF_save_fm DFF_P62(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0760));
DFF_save_fm DFF_P63(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0770));
DFF_save_fm DFF_P64(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0001));
DFF_save_fm DFF_P65(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0011));
DFF_save_fm DFF_P66(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0021));
DFF_save_fm DFF_P67(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0031));
DFF_save_fm DFF_P68(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0041));
DFF_save_fm DFF_P69(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0051));
DFF_save_fm DFF_P70(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0061));
DFF_save_fm DFF_P71(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0071));
DFF_save_fm DFF_P72(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0101));
DFF_save_fm DFF_P73(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0111));
DFF_save_fm DFF_P74(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0121));
DFF_save_fm DFF_P75(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0131));
DFF_save_fm DFF_P76(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0141));
DFF_save_fm DFF_P77(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0151));
DFF_save_fm DFF_P78(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0161));
DFF_save_fm DFF_P79(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0171));
DFF_save_fm DFF_P80(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0201));
DFF_save_fm DFF_P81(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0211));
DFF_save_fm DFF_P82(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0221));
DFF_save_fm DFF_P83(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0231));
DFF_save_fm DFF_P84(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0241));
DFF_save_fm DFF_P85(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0251));
DFF_save_fm DFF_P86(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0261));
DFF_save_fm DFF_P87(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0271));
DFF_save_fm DFF_P88(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0301));
DFF_save_fm DFF_P89(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0311));
DFF_save_fm DFF_P90(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0321));
DFF_save_fm DFF_P91(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0331));
DFF_save_fm DFF_P92(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0341));
DFF_save_fm DFF_P93(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0351));
DFF_save_fm DFF_P94(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0361));
DFF_save_fm DFF_P95(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0371));
DFF_save_fm DFF_P96(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0401));
DFF_save_fm DFF_P97(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0411));
DFF_save_fm DFF_P98(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0421));
DFF_save_fm DFF_P99(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0431));
DFF_save_fm DFF_P100(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0441));
DFF_save_fm DFF_P101(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0451));
DFF_save_fm DFF_P102(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0461));
DFF_save_fm DFF_P103(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0471));
DFF_save_fm DFF_P104(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0501));
DFF_save_fm DFF_P105(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0511));
DFF_save_fm DFF_P106(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0521));
DFF_save_fm DFF_P107(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0531));
DFF_save_fm DFF_P108(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0541));
DFF_save_fm DFF_P109(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0551));
DFF_save_fm DFF_P110(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0561));
DFF_save_fm DFF_P111(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0571));
DFF_save_fm DFF_P112(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0601));
DFF_save_fm DFF_P113(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0611));
DFF_save_fm DFF_P114(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0621));
DFF_save_fm DFF_P115(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0631));
DFF_save_fm DFF_P116(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0641));
DFF_save_fm DFF_P117(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0651));
DFF_save_fm DFF_P118(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0661));
DFF_save_fm DFF_P119(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0671));
DFF_save_fm DFF_P120(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0701));
DFF_save_fm DFF_P121(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0711));
DFF_save_fm DFF_P122(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0721));
DFF_save_fm DFF_P123(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0731));
DFF_save_fm DFF_P124(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0741));
DFF_save_fm DFF_P125(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0751));
DFF_save_fm DFF_P126(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0761));
DFF_save_fm DFF_P127(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0771));
DFF_save_fm DFF_P128(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0002));
DFF_save_fm DFF_P129(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0012));
DFF_save_fm DFF_P130(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0022));
DFF_save_fm DFF_P131(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0032));
DFF_save_fm DFF_P132(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0042));
DFF_save_fm DFF_P133(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0052));
DFF_save_fm DFF_P134(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0062));
DFF_save_fm DFF_P135(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0072));
DFF_save_fm DFF_P136(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0102));
DFF_save_fm DFF_P137(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0112));
DFF_save_fm DFF_P138(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0122));
DFF_save_fm DFF_P139(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0132));
DFF_save_fm DFF_P140(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0142));
DFF_save_fm DFF_P141(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0152));
DFF_save_fm DFF_P142(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0162));
DFF_save_fm DFF_P143(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0172));
DFF_save_fm DFF_P144(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0202));
DFF_save_fm DFF_P145(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0212));
DFF_save_fm DFF_P146(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0222));
DFF_save_fm DFF_P147(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0232));
DFF_save_fm DFF_P148(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0242));
DFF_save_fm DFF_P149(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0252));
DFF_save_fm DFF_P150(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0262));
DFF_save_fm DFF_P151(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0272));
DFF_save_fm DFF_P152(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0302));
DFF_save_fm DFF_P153(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0312));
DFF_save_fm DFF_P154(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0322));
DFF_save_fm DFF_P155(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0332));
DFF_save_fm DFF_P156(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0342));
DFF_save_fm DFF_P157(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0352));
DFF_save_fm DFF_P158(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0362));
DFF_save_fm DFF_P159(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0372));
DFF_save_fm DFF_P160(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0402));
DFF_save_fm DFF_P161(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0412));
DFF_save_fm DFF_P162(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0422));
DFF_save_fm DFF_P163(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0432));
DFF_save_fm DFF_P164(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0442));
DFF_save_fm DFF_P165(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0452));
DFF_save_fm DFF_P166(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0462));
DFF_save_fm DFF_P167(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0472));
DFF_save_fm DFF_P168(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0502));
DFF_save_fm DFF_P169(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0512));
DFF_save_fm DFF_P170(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0522));
DFF_save_fm DFF_P171(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0532));
DFF_save_fm DFF_P172(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0542));
DFF_save_fm DFF_P173(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0552));
DFF_save_fm DFF_P174(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0562));
DFF_save_fm DFF_P175(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0572));
DFF_save_fm DFF_P176(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0602));
DFF_save_fm DFF_P177(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0612));
DFF_save_fm DFF_P178(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0622));
DFF_save_fm DFF_P179(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0632));
DFF_save_fm DFF_P180(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0642));
DFF_save_fm DFF_P181(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0652));
DFF_save_fm DFF_P182(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0662));
DFF_save_fm DFF_P183(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0672));
DFF_save_fm DFF_P184(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0702));
DFF_save_fm DFF_P185(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0712));
DFF_save_fm DFF_P186(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0722));
DFF_save_fm DFF_P187(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0732));
DFF_save_fm DFF_P188(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0742));
DFF_save_fm DFF_P189(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0752));
DFF_save_fm DFF_P190(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0762));
DFF_save_fm DFF_P191(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0772));
DFF_save_fm DFF_W0(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00000));
DFF_save_fm DFF_W1(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00010));
DFF_save_fm DFF_W2(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00020));
DFF_save_fm DFF_W3(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00100));
DFF_save_fm DFF_W4(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00110));
DFF_save_fm DFF_W5(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00120));
DFF_save_fm DFF_W6(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00200));
DFF_save_fm DFF_W7(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00210));
DFF_save_fm DFF_W8(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00220));
DFF_save_fm DFF_W9(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00001));
DFF_save_fm DFF_W10(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00011));
DFF_save_fm DFF_W11(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00021));
DFF_save_fm DFF_W12(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00101));
DFF_save_fm DFF_W13(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00111));
DFF_save_fm DFF_W14(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00121));
DFF_save_fm DFF_W15(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00201));
DFF_save_fm DFF_W16(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00211));
DFF_save_fm DFF_W17(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00221));
DFF_save_fm DFF_W18(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00002));
DFF_save_fm DFF_W19(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00012));
DFF_save_fm DFF_W20(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00022));
DFF_save_fm DFF_W21(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00102));
DFF_save_fm DFF_W22(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00112));
DFF_save_fm DFF_W23(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00122));
DFF_save_fm DFF_W24(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00202));
DFF_save_fm DFF_W25(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00212));
DFF_save_fm DFF_W26(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00222));
DFF_save_fm DFF_W27(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01000));
DFF_save_fm DFF_W28(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01010));
DFF_save_fm DFF_W29(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01020));
DFF_save_fm DFF_W30(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01100));
DFF_save_fm DFF_W31(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01110));
DFF_save_fm DFF_W32(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01120));
DFF_save_fm DFF_W33(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01200));
DFF_save_fm DFF_W34(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01210));
DFF_save_fm DFF_W35(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01220));
DFF_save_fm DFF_W36(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01001));
DFF_save_fm DFF_W37(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01011));
DFF_save_fm DFF_W38(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01021));
DFF_save_fm DFF_W39(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01101));
DFF_save_fm DFF_W40(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01111));
DFF_save_fm DFF_W41(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01121));
DFF_save_fm DFF_W42(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01201));
DFF_save_fm DFF_W43(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01211));
DFF_save_fm DFF_W44(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01221));
DFF_save_fm DFF_W45(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01002));
DFF_save_fm DFF_W46(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01012));
DFF_save_fm DFF_W47(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01022));
DFF_save_fm DFF_W48(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01102));
DFF_save_fm DFF_W49(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01112));
DFF_save_fm DFF_W50(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01122));
DFF_save_fm DFF_W51(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01202));
DFF_save_fm DFF_W52(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01212));
DFF_save_fm DFF_W53(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01222));
DFF_save_fm DFF_W54(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02000));
DFF_save_fm DFF_W55(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02010));
DFF_save_fm DFF_W56(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02020));
DFF_save_fm DFF_W57(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02100));
DFF_save_fm DFF_W58(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02110));
DFF_save_fm DFF_W59(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02120));
DFF_save_fm DFF_W60(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02200));
DFF_save_fm DFF_W61(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02210));
DFF_save_fm DFF_W62(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02220));
DFF_save_fm DFF_W63(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02001));
DFF_save_fm DFF_W64(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02011));
DFF_save_fm DFF_W65(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02021));
DFF_save_fm DFF_W66(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02101));
DFF_save_fm DFF_W67(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02111));
DFF_save_fm DFF_W68(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02121));
DFF_save_fm DFF_W69(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02201));
DFF_save_fm DFF_W70(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02211));
DFF_save_fm DFF_W71(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02221));
DFF_save_fm DFF_W72(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02002));
DFF_save_fm DFF_W73(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02012));
DFF_save_fm DFF_W74(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02022));
DFF_save_fm DFF_W75(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02102));
DFF_save_fm DFF_W76(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02112));
DFF_save_fm DFF_W77(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02122));
DFF_save_fm DFF_W78(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02202));
DFF_save_fm DFF_W79(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02212));
DFF_save_fm DFF_W80(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02222));
DFF_save_fm DFF_W81(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03000));
DFF_save_fm DFF_W82(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03010));
DFF_save_fm DFF_W83(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03020));
DFF_save_fm DFF_W84(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03100));
DFF_save_fm DFF_W85(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03110));
DFF_save_fm DFF_W86(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03120));
DFF_save_fm DFF_W87(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03200));
DFF_save_fm DFF_W88(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03210));
DFF_save_fm DFF_W89(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03220));
DFF_save_fm DFF_W90(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03001));
DFF_save_fm DFF_W91(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03011));
DFF_save_fm DFF_W92(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03021));
DFF_save_fm DFF_W93(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03101));
DFF_save_fm DFF_W94(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03111));
DFF_save_fm DFF_W95(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03121));
DFF_save_fm DFF_W96(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03201));
DFF_save_fm DFF_W97(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03211));
DFF_save_fm DFF_W98(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03221));
DFF_save_fm DFF_W99(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03002));
DFF_save_fm DFF_W100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03012));
DFF_save_fm DFF_W101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03022));
DFF_save_fm DFF_W102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03102));
DFF_save_fm DFF_W103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03112));
DFF_save_fm DFF_W104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03122));
DFF_save_fm DFF_W105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W03202));
DFF_save_fm DFF_W106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03212));
DFF_save_fm DFF_W107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W03222));
ninexnine_unit ninexnine_unit_0(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00000)
);

ninexnine_unit ninexnine_unit_1(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01000)
);

ninexnine_unit ninexnine_unit_2(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02000)
);

assign C0000=c00000+c01000+c02000;
assign A0000=(C0000>=0)?1:0;

ninexnine_unit ninexnine_unit_3(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00010)
);

ninexnine_unit ninexnine_unit_4(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01010)
);

ninexnine_unit ninexnine_unit_5(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02010)
);

assign C0010=c00010+c01010+c02010;
assign A0010=(C0010>=0)?1:0;

ninexnine_unit ninexnine_unit_6(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00020)
);

ninexnine_unit ninexnine_unit_7(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01020)
);

ninexnine_unit ninexnine_unit_8(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02020)
);

assign C0020=c00020+c01020+c02020;
assign A0020=(C0020>=0)?1:0;

ninexnine_unit ninexnine_unit_9(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00030)
);

ninexnine_unit ninexnine_unit_10(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01030)
);

ninexnine_unit ninexnine_unit_11(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02030)
);

assign C0030=c00030+c01030+c02030;
assign A0030=(C0030>=0)?1:0;

ninexnine_unit ninexnine_unit_12(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00040)
);

ninexnine_unit ninexnine_unit_13(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01040)
);

ninexnine_unit ninexnine_unit_14(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02040)
);

assign C0040=c00040+c01040+c02040;
assign A0040=(C0040>=0)?1:0;

ninexnine_unit ninexnine_unit_15(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00050)
);

ninexnine_unit ninexnine_unit_16(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01050)
);

ninexnine_unit ninexnine_unit_17(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02050)
);

assign C0050=c00050+c01050+c02050;
assign A0050=(C0050>=0)?1:0;

ninexnine_unit ninexnine_unit_18(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00100)
);

ninexnine_unit ninexnine_unit_19(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01100)
);

ninexnine_unit ninexnine_unit_20(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02100)
);

assign C0100=c00100+c01100+c02100;
assign A0100=(C0100>=0)?1:0;

ninexnine_unit ninexnine_unit_21(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00110)
);

ninexnine_unit ninexnine_unit_22(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01110)
);

ninexnine_unit ninexnine_unit_23(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02110)
);

assign C0110=c00110+c01110+c02110;
assign A0110=(C0110>=0)?1:0;

ninexnine_unit ninexnine_unit_24(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00120)
);

ninexnine_unit ninexnine_unit_25(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01120)
);

ninexnine_unit ninexnine_unit_26(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02120)
);

assign C0120=c00120+c01120+c02120;
assign A0120=(C0120>=0)?1:0;

ninexnine_unit ninexnine_unit_27(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00130)
);

ninexnine_unit ninexnine_unit_28(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01130)
);

ninexnine_unit ninexnine_unit_29(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02130)
);

assign C0130=c00130+c01130+c02130;
assign A0130=(C0130>=0)?1:0;

ninexnine_unit ninexnine_unit_30(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00140)
);

ninexnine_unit ninexnine_unit_31(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01140)
);

ninexnine_unit ninexnine_unit_32(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02140)
);

assign C0140=c00140+c01140+c02140;
assign A0140=(C0140>=0)?1:0;

ninexnine_unit ninexnine_unit_33(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00150)
);

ninexnine_unit ninexnine_unit_34(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01150)
);

ninexnine_unit ninexnine_unit_35(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02150)
);

assign C0150=c00150+c01150+c02150;
assign A0150=(C0150>=0)?1:0;

ninexnine_unit ninexnine_unit_36(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00200)
);

ninexnine_unit ninexnine_unit_37(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01200)
);

ninexnine_unit ninexnine_unit_38(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02200)
);

assign C0200=c00200+c01200+c02200;
assign A0200=(C0200>=0)?1:0;

ninexnine_unit ninexnine_unit_39(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00210)
);

ninexnine_unit ninexnine_unit_40(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01210)
);

ninexnine_unit ninexnine_unit_41(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02210)
);

assign C0210=c00210+c01210+c02210;
assign A0210=(C0210>=0)?1:0;

ninexnine_unit ninexnine_unit_42(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00220)
);

ninexnine_unit ninexnine_unit_43(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01220)
);

ninexnine_unit ninexnine_unit_44(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02220)
);

assign C0220=c00220+c01220+c02220;
assign A0220=(C0220>=0)?1:0;

ninexnine_unit ninexnine_unit_45(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00230)
);

ninexnine_unit ninexnine_unit_46(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01230)
);

ninexnine_unit ninexnine_unit_47(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02230)
);

assign C0230=c00230+c01230+c02230;
assign A0230=(C0230>=0)?1:0;

ninexnine_unit ninexnine_unit_48(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00240)
);

ninexnine_unit ninexnine_unit_49(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01240)
);

ninexnine_unit ninexnine_unit_50(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02240)
);

assign C0240=c00240+c01240+c02240;
assign A0240=(C0240>=0)?1:0;

ninexnine_unit ninexnine_unit_51(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00250)
);

ninexnine_unit ninexnine_unit_52(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01250)
);

ninexnine_unit ninexnine_unit_53(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02250)
);

assign C0250=c00250+c01250+c02250;
assign A0250=(C0250>=0)?1:0;

ninexnine_unit ninexnine_unit_54(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00300)
);

ninexnine_unit ninexnine_unit_55(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01300)
);

ninexnine_unit ninexnine_unit_56(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02300)
);

assign C0300=c00300+c01300+c02300;
assign A0300=(C0300>=0)?1:0;

ninexnine_unit ninexnine_unit_57(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00310)
);

ninexnine_unit ninexnine_unit_58(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01310)
);

ninexnine_unit ninexnine_unit_59(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02310)
);

assign C0310=c00310+c01310+c02310;
assign A0310=(C0310>=0)?1:0;

ninexnine_unit ninexnine_unit_60(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00320)
);

ninexnine_unit ninexnine_unit_61(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01320)
);

ninexnine_unit ninexnine_unit_62(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02320)
);

assign C0320=c00320+c01320+c02320;
assign A0320=(C0320>=0)?1:0;

ninexnine_unit ninexnine_unit_63(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00330)
);

ninexnine_unit ninexnine_unit_64(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01330)
);

ninexnine_unit ninexnine_unit_65(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02330)
);

assign C0330=c00330+c01330+c02330;
assign A0330=(C0330>=0)?1:0;

ninexnine_unit ninexnine_unit_66(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00340)
);

ninexnine_unit ninexnine_unit_67(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01340)
);

ninexnine_unit ninexnine_unit_68(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02340)
);

assign C0340=c00340+c01340+c02340;
assign A0340=(C0340>=0)?1:0;

ninexnine_unit ninexnine_unit_69(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00350)
);

ninexnine_unit ninexnine_unit_70(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01350)
);

ninexnine_unit ninexnine_unit_71(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02350)
);

assign C0350=c00350+c01350+c02350;
assign A0350=(C0350>=0)?1:0;

ninexnine_unit ninexnine_unit_72(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00400)
);

ninexnine_unit ninexnine_unit_73(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01400)
);

ninexnine_unit ninexnine_unit_74(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02400)
);

assign C0400=c00400+c01400+c02400;
assign A0400=(C0400>=0)?1:0;

ninexnine_unit ninexnine_unit_75(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00410)
);

ninexnine_unit ninexnine_unit_76(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01410)
);

ninexnine_unit ninexnine_unit_77(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02410)
);

assign C0410=c00410+c01410+c02410;
assign A0410=(C0410>=0)?1:0;

ninexnine_unit ninexnine_unit_78(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00420)
);

ninexnine_unit ninexnine_unit_79(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01420)
);

ninexnine_unit ninexnine_unit_80(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02420)
);

assign C0420=c00420+c01420+c02420;
assign A0420=(C0420>=0)?1:0;

ninexnine_unit ninexnine_unit_81(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00430)
);

ninexnine_unit ninexnine_unit_82(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01430)
);

ninexnine_unit ninexnine_unit_83(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02430)
);

assign C0430=c00430+c01430+c02430;
assign A0430=(C0430>=0)?1:0;

ninexnine_unit ninexnine_unit_84(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00440)
);

ninexnine_unit ninexnine_unit_85(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01440)
);

ninexnine_unit ninexnine_unit_86(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02440)
);

assign C0440=c00440+c01440+c02440;
assign A0440=(C0440>=0)?1:0;

ninexnine_unit ninexnine_unit_87(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00450)
);

ninexnine_unit ninexnine_unit_88(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01450)
);

ninexnine_unit ninexnine_unit_89(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02450)
);

assign C0450=c00450+c01450+c02450;
assign A0450=(C0450>=0)?1:0;

ninexnine_unit ninexnine_unit_90(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00500)
);

ninexnine_unit ninexnine_unit_91(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01500)
);

ninexnine_unit ninexnine_unit_92(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02500)
);

assign C0500=c00500+c01500+c02500;
assign A0500=(C0500>=0)?1:0;

ninexnine_unit ninexnine_unit_93(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00510)
);

ninexnine_unit ninexnine_unit_94(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01510)
);

ninexnine_unit ninexnine_unit_95(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02510)
);

assign C0510=c00510+c01510+c02510;
assign A0510=(C0510>=0)?1:0;

ninexnine_unit ninexnine_unit_96(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00520)
);

ninexnine_unit ninexnine_unit_97(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01520)
);

ninexnine_unit ninexnine_unit_98(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02520)
);

assign C0520=c00520+c01520+c02520;
assign A0520=(C0520>=0)?1:0;

ninexnine_unit ninexnine_unit_99(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00530)
);

ninexnine_unit ninexnine_unit_100(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01530)
);

ninexnine_unit ninexnine_unit_101(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02530)
);

assign C0530=c00530+c01530+c02530;
assign A0530=(C0530>=0)?1:0;

ninexnine_unit ninexnine_unit_102(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00540)
);

ninexnine_unit ninexnine_unit_103(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01540)
);

ninexnine_unit ninexnine_unit_104(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02540)
);

assign C0540=c00540+c01540+c02540;
assign A0540=(C0540>=0)?1:0;

ninexnine_unit ninexnine_unit_105(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00550)
);

ninexnine_unit ninexnine_unit_106(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01550)
);

ninexnine_unit ninexnine_unit_107(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02550)
);

assign C0550=c00550+c01550+c02550;
assign A0550=(C0550>=0)?1:0;

ninexnine_unit ninexnine_unit_108(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00001)
);

ninexnine_unit ninexnine_unit_109(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01001)
);

ninexnine_unit ninexnine_unit_110(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02001)
);

assign C0001=c00001+c01001+c02001;
assign A0001=(C0001>=0)?1:0;

ninexnine_unit ninexnine_unit_111(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00011)
);

ninexnine_unit ninexnine_unit_112(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01011)
);

ninexnine_unit ninexnine_unit_113(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02011)
);

assign C0011=c00011+c01011+c02011;
assign A0011=(C0011>=0)?1:0;

ninexnine_unit ninexnine_unit_114(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00021)
);

ninexnine_unit ninexnine_unit_115(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01021)
);

ninexnine_unit ninexnine_unit_116(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02021)
);

assign C0021=c00021+c01021+c02021;
assign A0021=(C0021>=0)?1:0;

ninexnine_unit ninexnine_unit_117(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00031)
);

ninexnine_unit ninexnine_unit_118(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01031)
);

ninexnine_unit ninexnine_unit_119(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02031)
);

assign C0031=c00031+c01031+c02031;
assign A0031=(C0031>=0)?1:0;

ninexnine_unit ninexnine_unit_120(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00041)
);

ninexnine_unit ninexnine_unit_121(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01041)
);

ninexnine_unit ninexnine_unit_122(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02041)
);

assign C0041=c00041+c01041+c02041;
assign A0041=(C0041>=0)?1:0;

ninexnine_unit ninexnine_unit_123(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00051)
);

ninexnine_unit ninexnine_unit_124(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01051)
);

ninexnine_unit ninexnine_unit_125(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02051)
);

assign C0051=c00051+c01051+c02051;
assign A0051=(C0051>=0)?1:0;

ninexnine_unit ninexnine_unit_126(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00101)
);

ninexnine_unit ninexnine_unit_127(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01101)
);

ninexnine_unit ninexnine_unit_128(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02101)
);

assign C0101=c00101+c01101+c02101;
assign A0101=(C0101>=0)?1:0;

ninexnine_unit ninexnine_unit_129(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00111)
);

ninexnine_unit ninexnine_unit_130(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01111)
);

ninexnine_unit ninexnine_unit_131(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02111)
);

assign C0111=c00111+c01111+c02111;
assign A0111=(C0111>=0)?1:0;

ninexnine_unit ninexnine_unit_132(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00121)
);

ninexnine_unit ninexnine_unit_133(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01121)
);

ninexnine_unit ninexnine_unit_134(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02121)
);

assign C0121=c00121+c01121+c02121;
assign A0121=(C0121>=0)?1:0;

ninexnine_unit ninexnine_unit_135(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00131)
);

ninexnine_unit ninexnine_unit_136(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01131)
);

ninexnine_unit ninexnine_unit_137(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02131)
);

assign C0131=c00131+c01131+c02131;
assign A0131=(C0131>=0)?1:0;

ninexnine_unit ninexnine_unit_138(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00141)
);

ninexnine_unit ninexnine_unit_139(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01141)
);

ninexnine_unit ninexnine_unit_140(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02141)
);

assign C0141=c00141+c01141+c02141;
assign A0141=(C0141>=0)?1:0;

ninexnine_unit ninexnine_unit_141(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00151)
);

ninexnine_unit ninexnine_unit_142(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01151)
);

ninexnine_unit ninexnine_unit_143(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02151)
);

assign C0151=c00151+c01151+c02151;
assign A0151=(C0151>=0)?1:0;

ninexnine_unit ninexnine_unit_144(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00201)
);

ninexnine_unit ninexnine_unit_145(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01201)
);

ninexnine_unit ninexnine_unit_146(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02201)
);

assign C0201=c00201+c01201+c02201;
assign A0201=(C0201>=0)?1:0;

ninexnine_unit ninexnine_unit_147(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00211)
);

ninexnine_unit ninexnine_unit_148(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01211)
);

ninexnine_unit ninexnine_unit_149(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02211)
);

assign C0211=c00211+c01211+c02211;
assign A0211=(C0211>=0)?1:0;

ninexnine_unit ninexnine_unit_150(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00221)
);

ninexnine_unit ninexnine_unit_151(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01221)
);

ninexnine_unit ninexnine_unit_152(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02221)
);

assign C0221=c00221+c01221+c02221;
assign A0221=(C0221>=0)?1:0;

ninexnine_unit ninexnine_unit_153(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00231)
);

ninexnine_unit ninexnine_unit_154(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01231)
);

ninexnine_unit ninexnine_unit_155(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02231)
);

assign C0231=c00231+c01231+c02231;
assign A0231=(C0231>=0)?1:0;

ninexnine_unit ninexnine_unit_156(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00241)
);

ninexnine_unit ninexnine_unit_157(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01241)
);

ninexnine_unit ninexnine_unit_158(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02241)
);

assign C0241=c00241+c01241+c02241;
assign A0241=(C0241>=0)?1:0;

ninexnine_unit ninexnine_unit_159(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00251)
);

ninexnine_unit ninexnine_unit_160(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01251)
);

ninexnine_unit ninexnine_unit_161(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02251)
);

assign C0251=c00251+c01251+c02251;
assign A0251=(C0251>=0)?1:0;

ninexnine_unit ninexnine_unit_162(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00301)
);

ninexnine_unit ninexnine_unit_163(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01301)
);

ninexnine_unit ninexnine_unit_164(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02301)
);

assign C0301=c00301+c01301+c02301;
assign A0301=(C0301>=0)?1:0;

ninexnine_unit ninexnine_unit_165(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00311)
);

ninexnine_unit ninexnine_unit_166(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01311)
);

ninexnine_unit ninexnine_unit_167(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02311)
);

assign C0311=c00311+c01311+c02311;
assign A0311=(C0311>=0)?1:0;

ninexnine_unit ninexnine_unit_168(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00321)
);

ninexnine_unit ninexnine_unit_169(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01321)
);

ninexnine_unit ninexnine_unit_170(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02321)
);

assign C0321=c00321+c01321+c02321;
assign A0321=(C0321>=0)?1:0;

ninexnine_unit ninexnine_unit_171(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00331)
);

ninexnine_unit ninexnine_unit_172(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01331)
);

ninexnine_unit ninexnine_unit_173(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02331)
);

assign C0331=c00331+c01331+c02331;
assign A0331=(C0331>=0)?1:0;

ninexnine_unit ninexnine_unit_174(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00341)
);

ninexnine_unit ninexnine_unit_175(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01341)
);

ninexnine_unit ninexnine_unit_176(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02341)
);

assign C0341=c00341+c01341+c02341;
assign A0341=(C0341>=0)?1:0;

ninexnine_unit ninexnine_unit_177(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00351)
);

ninexnine_unit ninexnine_unit_178(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01351)
);

ninexnine_unit ninexnine_unit_179(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02351)
);

assign C0351=c00351+c01351+c02351;
assign A0351=(C0351>=0)?1:0;

ninexnine_unit ninexnine_unit_180(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00401)
);

ninexnine_unit ninexnine_unit_181(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01401)
);

ninexnine_unit ninexnine_unit_182(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02401)
);

assign C0401=c00401+c01401+c02401;
assign A0401=(C0401>=0)?1:0;

ninexnine_unit ninexnine_unit_183(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00411)
);

ninexnine_unit ninexnine_unit_184(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01411)
);

ninexnine_unit ninexnine_unit_185(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02411)
);

assign C0411=c00411+c01411+c02411;
assign A0411=(C0411>=0)?1:0;

ninexnine_unit ninexnine_unit_186(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00421)
);

ninexnine_unit ninexnine_unit_187(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01421)
);

ninexnine_unit ninexnine_unit_188(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02421)
);

assign C0421=c00421+c01421+c02421;
assign A0421=(C0421>=0)?1:0;

ninexnine_unit ninexnine_unit_189(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00431)
);

ninexnine_unit ninexnine_unit_190(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01431)
);

ninexnine_unit ninexnine_unit_191(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02431)
);

assign C0431=c00431+c01431+c02431;
assign A0431=(C0431>=0)?1:0;

ninexnine_unit ninexnine_unit_192(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00441)
);

ninexnine_unit ninexnine_unit_193(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01441)
);

ninexnine_unit ninexnine_unit_194(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02441)
);

assign C0441=c00441+c01441+c02441;
assign A0441=(C0441>=0)?1:0;

ninexnine_unit ninexnine_unit_195(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00451)
);

ninexnine_unit ninexnine_unit_196(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01451)
);

ninexnine_unit ninexnine_unit_197(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02451)
);

assign C0451=c00451+c01451+c02451;
assign A0451=(C0451>=0)?1:0;

ninexnine_unit ninexnine_unit_198(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00501)
);

ninexnine_unit ninexnine_unit_199(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01501)
);

ninexnine_unit ninexnine_unit_200(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02501)
);

assign C0501=c00501+c01501+c02501;
assign A0501=(C0501>=0)?1:0;

ninexnine_unit ninexnine_unit_201(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00511)
);

ninexnine_unit ninexnine_unit_202(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01511)
);

ninexnine_unit ninexnine_unit_203(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02511)
);

assign C0511=c00511+c01511+c02511;
assign A0511=(C0511>=0)?1:0;

ninexnine_unit ninexnine_unit_204(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00521)
);

ninexnine_unit ninexnine_unit_205(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01521)
);

ninexnine_unit ninexnine_unit_206(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02521)
);

assign C0521=c00521+c01521+c02521;
assign A0521=(C0521>=0)?1:0;

ninexnine_unit ninexnine_unit_207(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00531)
);

ninexnine_unit ninexnine_unit_208(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01531)
);

ninexnine_unit ninexnine_unit_209(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02531)
);

assign C0531=c00531+c01531+c02531;
assign A0531=(C0531>=0)?1:0;

ninexnine_unit ninexnine_unit_210(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00541)
);

ninexnine_unit ninexnine_unit_211(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01541)
);

ninexnine_unit ninexnine_unit_212(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02541)
);

assign C0541=c00541+c01541+c02541;
assign A0541=(C0541>=0)?1:0;

ninexnine_unit ninexnine_unit_213(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00551)
);

ninexnine_unit ninexnine_unit_214(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01551)
);

ninexnine_unit ninexnine_unit_215(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02551)
);

assign C0551=c00551+c01551+c02551;
assign A0551=(C0551>=0)?1:0;

ninexnine_unit ninexnine_unit_216(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00002)
);

ninexnine_unit ninexnine_unit_217(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01002)
);

ninexnine_unit ninexnine_unit_218(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02002)
);

assign C0002=c00002+c01002+c02002;
assign A0002=(C0002>=0)?1:0;

ninexnine_unit ninexnine_unit_219(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00012)
);

ninexnine_unit ninexnine_unit_220(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01012)
);

ninexnine_unit ninexnine_unit_221(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02012)
);

assign C0012=c00012+c01012+c02012;
assign A0012=(C0012>=0)?1:0;

ninexnine_unit ninexnine_unit_222(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00022)
);

ninexnine_unit ninexnine_unit_223(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01022)
);

ninexnine_unit ninexnine_unit_224(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02022)
);

assign C0022=c00022+c01022+c02022;
assign A0022=(C0022>=0)?1:0;

ninexnine_unit ninexnine_unit_225(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00032)
);

ninexnine_unit ninexnine_unit_226(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01032)
);

ninexnine_unit ninexnine_unit_227(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02032)
);

assign C0032=c00032+c01032+c02032;
assign A0032=(C0032>=0)?1:0;

ninexnine_unit ninexnine_unit_228(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00042)
);

ninexnine_unit ninexnine_unit_229(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01042)
);

ninexnine_unit ninexnine_unit_230(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02042)
);

assign C0042=c00042+c01042+c02042;
assign A0042=(C0042>=0)?1:0;

ninexnine_unit ninexnine_unit_231(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00052)
);

ninexnine_unit ninexnine_unit_232(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01052)
);

ninexnine_unit ninexnine_unit_233(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02052)
);

assign C0052=c00052+c01052+c02052;
assign A0052=(C0052>=0)?1:0;

ninexnine_unit ninexnine_unit_234(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00102)
);

ninexnine_unit ninexnine_unit_235(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01102)
);

ninexnine_unit ninexnine_unit_236(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02102)
);

assign C0102=c00102+c01102+c02102;
assign A0102=(C0102>=0)?1:0;

ninexnine_unit ninexnine_unit_237(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00112)
);

ninexnine_unit ninexnine_unit_238(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01112)
);

ninexnine_unit ninexnine_unit_239(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02112)
);

assign C0112=c00112+c01112+c02112;
assign A0112=(C0112>=0)?1:0;

ninexnine_unit ninexnine_unit_240(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00122)
);

ninexnine_unit ninexnine_unit_241(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01122)
);

ninexnine_unit ninexnine_unit_242(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02122)
);

assign C0122=c00122+c01122+c02122;
assign A0122=(C0122>=0)?1:0;

ninexnine_unit ninexnine_unit_243(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00132)
);

ninexnine_unit ninexnine_unit_244(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01132)
);

ninexnine_unit ninexnine_unit_245(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02132)
);

assign C0132=c00132+c01132+c02132;
assign A0132=(C0132>=0)?1:0;

ninexnine_unit ninexnine_unit_246(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00142)
);

ninexnine_unit ninexnine_unit_247(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01142)
);

ninexnine_unit ninexnine_unit_248(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02142)
);

assign C0142=c00142+c01142+c02142;
assign A0142=(C0142>=0)?1:0;

ninexnine_unit ninexnine_unit_249(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00152)
);

ninexnine_unit ninexnine_unit_250(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01152)
);

ninexnine_unit ninexnine_unit_251(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02152)
);

assign C0152=c00152+c01152+c02152;
assign A0152=(C0152>=0)?1:0;

ninexnine_unit ninexnine_unit_252(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00202)
);

ninexnine_unit ninexnine_unit_253(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01202)
);

ninexnine_unit ninexnine_unit_254(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02202)
);

assign C0202=c00202+c01202+c02202;
assign A0202=(C0202>=0)?1:0;

ninexnine_unit ninexnine_unit_255(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00212)
);

ninexnine_unit ninexnine_unit_256(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01212)
);

ninexnine_unit ninexnine_unit_257(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02212)
);

assign C0212=c00212+c01212+c02212;
assign A0212=(C0212>=0)?1:0;

ninexnine_unit ninexnine_unit_258(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00222)
);

ninexnine_unit ninexnine_unit_259(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01222)
);

ninexnine_unit ninexnine_unit_260(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02222)
);

assign C0222=c00222+c01222+c02222;
assign A0222=(C0222>=0)?1:0;

ninexnine_unit ninexnine_unit_261(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00232)
);

ninexnine_unit ninexnine_unit_262(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01232)
);

ninexnine_unit ninexnine_unit_263(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02232)
);

assign C0232=c00232+c01232+c02232;
assign A0232=(C0232>=0)?1:0;

ninexnine_unit ninexnine_unit_264(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00242)
);

ninexnine_unit ninexnine_unit_265(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01242)
);

ninexnine_unit ninexnine_unit_266(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02242)
);

assign C0242=c00242+c01242+c02242;
assign A0242=(C0242>=0)?1:0;

ninexnine_unit ninexnine_unit_267(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00252)
);

ninexnine_unit ninexnine_unit_268(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01252)
);

ninexnine_unit ninexnine_unit_269(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02252)
);

assign C0252=c00252+c01252+c02252;
assign A0252=(C0252>=0)?1:0;

ninexnine_unit ninexnine_unit_270(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00302)
);

ninexnine_unit ninexnine_unit_271(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01302)
);

ninexnine_unit ninexnine_unit_272(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02302)
);

assign C0302=c00302+c01302+c02302;
assign A0302=(C0302>=0)?1:0;

ninexnine_unit ninexnine_unit_273(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00312)
);

ninexnine_unit ninexnine_unit_274(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01312)
);

ninexnine_unit ninexnine_unit_275(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02312)
);

assign C0312=c00312+c01312+c02312;
assign A0312=(C0312>=0)?1:0;

ninexnine_unit ninexnine_unit_276(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00322)
);

ninexnine_unit ninexnine_unit_277(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01322)
);

ninexnine_unit ninexnine_unit_278(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02322)
);

assign C0322=c00322+c01322+c02322;
assign A0322=(C0322>=0)?1:0;

ninexnine_unit ninexnine_unit_279(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00332)
);

ninexnine_unit ninexnine_unit_280(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01332)
);

ninexnine_unit ninexnine_unit_281(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02332)
);

assign C0332=c00332+c01332+c02332;
assign A0332=(C0332>=0)?1:0;

ninexnine_unit ninexnine_unit_282(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00342)
);

ninexnine_unit ninexnine_unit_283(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01342)
);

ninexnine_unit ninexnine_unit_284(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02342)
);

assign C0342=c00342+c01342+c02342;
assign A0342=(C0342>=0)?1:0;

ninexnine_unit ninexnine_unit_285(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00352)
);

ninexnine_unit ninexnine_unit_286(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01352)
);

ninexnine_unit ninexnine_unit_287(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02352)
);

assign C0352=c00352+c01352+c02352;
assign A0352=(C0352>=0)?1:0;

ninexnine_unit ninexnine_unit_288(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00402)
);

ninexnine_unit ninexnine_unit_289(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01402)
);

ninexnine_unit ninexnine_unit_290(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02402)
);

assign C0402=c00402+c01402+c02402;
assign A0402=(C0402>=0)?1:0;

ninexnine_unit ninexnine_unit_291(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00412)
);

ninexnine_unit ninexnine_unit_292(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01412)
);

ninexnine_unit ninexnine_unit_293(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02412)
);

assign C0412=c00412+c01412+c02412;
assign A0412=(C0412>=0)?1:0;

ninexnine_unit ninexnine_unit_294(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00422)
);

ninexnine_unit ninexnine_unit_295(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01422)
);

ninexnine_unit ninexnine_unit_296(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02422)
);

assign C0422=c00422+c01422+c02422;
assign A0422=(C0422>=0)?1:0;

ninexnine_unit ninexnine_unit_297(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00432)
);

ninexnine_unit ninexnine_unit_298(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01432)
);

ninexnine_unit ninexnine_unit_299(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02432)
);

assign C0432=c00432+c01432+c02432;
assign A0432=(C0432>=0)?1:0;

ninexnine_unit ninexnine_unit_300(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00442)
);

ninexnine_unit ninexnine_unit_301(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01442)
);

ninexnine_unit ninexnine_unit_302(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02442)
);

assign C0442=c00442+c01442+c02442;
assign A0442=(C0442>=0)?1:0;

ninexnine_unit ninexnine_unit_303(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00452)
);

ninexnine_unit ninexnine_unit_304(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01452)
);

ninexnine_unit ninexnine_unit_305(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02452)
);

assign C0452=c00452+c01452+c02452;
assign A0452=(C0452>=0)?1:0;

ninexnine_unit ninexnine_unit_306(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00502)
);

ninexnine_unit ninexnine_unit_307(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01502)
);

ninexnine_unit ninexnine_unit_308(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02502)
);

assign C0502=c00502+c01502+c02502;
assign A0502=(C0502>=0)?1:0;

ninexnine_unit ninexnine_unit_309(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00512)
);

ninexnine_unit ninexnine_unit_310(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01512)
);

ninexnine_unit ninexnine_unit_311(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02512)
);

assign C0512=c00512+c01512+c02512;
assign A0512=(C0512>=0)?1:0;

ninexnine_unit ninexnine_unit_312(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00522)
);

ninexnine_unit ninexnine_unit_313(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01522)
);

ninexnine_unit ninexnine_unit_314(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02522)
);

assign C0522=c00522+c01522+c02522;
assign A0522=(C0522>=0)?1:0;

ninexnine_unit ninexnine_unit_315(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00532)
);

ninexnine_unit ninexnine_unit_316(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01532)
);

ninexnine_unit ninexnine_unit_317(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02532)
);

assign C0532=c00532+c01532+c02532;
assign A0532=(C0532>=0)?1:0;

ninexnine_unit ninexnine_unit_318(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00542)
);

ninexnine_unit ninexnine_unit_319(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01542)
);

ninexnine_unit ninexnine_unit_320(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02542)
);

assign C0542=c00542+c01542+c02542;
assign A0542=(C0542>=0)?1:0;

ninexnine_unit ninexnine_unit_321(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00552)
);

ninexnine_unit ninexnine_unit_322(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01552)
);

ninexnine_unit ninexnine_unit_323(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02552)
);

assign C0552=c00552+c01552+c02552;
assign A0552=(C0552>=0)?1:0;

ninexnine_unit ninexnine_unit_324(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00003)
);

ninexnine_unit ninexnine_unit_325(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01003)
);

ninexnine_unit ninexnine_unit_326(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02003)
);

assign C0003=c00003+c01003+c02003;
assign A0003=(C0003>=0)?1:0;

ninexnine_unit ninexnine_unit_327(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00013)
);

ninexnine_unit ninexnine_unit_328(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01013)
);

ninexnine_unit ninexnine_unit_329(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02013)
);

assign C0013=c00013+c01013+c02013;
assign A0013=(C0013>=0)?1:0;

ninexnine_unit ninexnine_unit_330(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00023)
);

ninexnine_unit ninexnine_unit_331(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01023)
);

ninexnine_unit ninexnine_unit_332(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02023)
);

assign C0023=c00023+c01023+c02023;
assign A0023=(C0023>=0)?1:0;

ninexnine_unit ninexnine_unit_333(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00033)
);

ninexnine_unit ninexnine_unit_334(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01033)
);

ninexnine_unit ninexnine_unit_335(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02033)
);

assign C0033=c00033+c01033+c02033;
assign A0033=(C0033>=0)?1:0;

ninexnine_unit ninexnine_unit_336(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00043)
);

ninexnine_unit ninexnine_unit_337(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01043)
);

ninexnine_unit ninexnine_unit_338(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02043)
);

assign C0043=c00043+c01043+c02043;
assign A0043=(C0043>=0)?1:0;

ninexnine_unit ninexnine_unit_339(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00053)
);

ninexnine_unit ninexnine_unit_340(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01053)
);

ninexnine_unit ninexnine_unit_341(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02053)
);

assign C0053=c00053+c01053+c02053;
assign A0053=(C0053>=0)?1:0;

ninexnine_unit ninexnine_unit_342(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00103)
);

ninexnine_unit ninexnine_unit_343(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01103)
);

ninexnine_unit ninexnine_unit_344(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02103)
);

assign C0103=c00103+c01103+c02103;
assign A0103=(C0103>=0)?1:0;

ninexnine_unit ninexnine_unit_345(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00113)
);

ninexnine_unit ninexnine_unit_346(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01113)
);

ninexnine_unit ninexnine_unit_347(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02113)
);

assign C0113=c00113+c01113+c02113;
assign A0113=(C0113>=0)?1:0;

ninexnine_unit ninexnine_unit_348(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00123)
);

ninexnine_unit ninexnine_unit_349(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01123)
);

ninexnine_unit ninexnine_unit_350(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02123)
);

assign C0123=c00123+c01123+c02123;
assign A0123=(C0123>=0)?1:0;

ninexnine_unit ninexnine_unit_351(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00133)
);

ninexnine_unit ninexnine_unit_352(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01133)
);

ninexnine_unit ninexnine_unit_353(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02133)
);

assign C0133=c00133+c01133+c02133;
assign A0133=(C0133>=0)?1:0;

ninexnine_unit ninexnine_unit_354(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00143)
);

ninexnine_unit ninexnine_unit_355(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01143)
);

ninexnine_unit ninexnine_unit_356(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02143)
);

assign C0143=c00143+c01143+c02143;
assign A0143=(C0143>=0)?1:0;

ninexnine_unit ninexnine_unit_357(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00153)
);

ninexnine_unit ninexnine_unit_358(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01153)
);

ninexnine_unit ninexnine_unit_359(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02153)
);

assign C0153=c00153+c01153+c02153;
assign A0153=(C0153>=0)?1:0;

ninexnine_unit ninexnine_unit_360(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00203)
);

ninexnine_unit ninexnine_unit_361(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01203)
);

ninexnine_unit ninexnine_unit_362(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02203)
);

assign C0203=c00203+c01203+c02203;
assign A0203=(C0203>=0)?1:0;

ninexnine_unit ninexnine_unit_363(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00213)
);

ninexnine_unit ninexnine_unit_364(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01213)
);

ninexnine_unit ninexnine_unit_365(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02213)
);

assign C0213=c00213+c01213+c02213;
assign A0213=(C0213>=0)?1:0;

ninexnine_unit ninexnine_unit_366(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00223)
);

ninexnine_unit ninexnine_unit_367(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01223)
);

ninexnine_unit ninexnine_unit_368(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02223)
);

assign C0223=c00223+c01223+c02223;
assign A0223=(C0223>=0)?1:0;

ninexnine_unit ninexnine_unit_369(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00233)
);

ninexnine_unit ninexnine_unit_370(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01233)
);

ninexnine_unit ninexnine_unit_371(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02233)
);

assign C0233=c00233+c01233+c02233;
assign A0233=(C0233>=0)?1:0;

ninexnine_unit ninexnine_unit_372(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00243)
);

ninexnine_unit ninexnine_unit_373(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01243)
);

ninexnine_unit ninexnine_unit_374(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02243)
);

assign C0243=c00243+c01243+c02243;
assign A0243=(C0243>=0)?1:0;

ninexnine_unit ninexnine_unit_375(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00253)
);

ninexnine_unit ninexnine_unit_376(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01253)
);

ninexnine_unit ninexnine_unit_377(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02253)
);

assign C0253=c00253+c01253+c02253;
assign A0253=(C0253>=0)?1:0;

ninexnine_unit ninexnine_unit_378(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00303)
);

ninexnine_unit ninexnine_unit_379(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01303)
);

ninexnine_unit ninexnine_unit_380(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02303)
);

assign C0303=c00303+c01303+c02303;
assign A0303=(C0303>=0)?1:0;

ninexnine_unit ninexnine_unit_381(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00313)
);

ninexnine_unit ninexnine_unit_382(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01313)
);

ninexnine_unit ninexnine_unit_383(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02313)
);

assign C0313=c00313+c01313+c02313;
assign A0313=(C0313>=0)?1:0;

ninexnine_unit ninexnine_unit_384(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00323)
);

ninexnine_unit ninexnine_unit_385(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01323)
);

ninexnine_unit ninexnine_unit_386(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02323)
);

assign C0323=c00323+c01323+c02323;
assign A0323=(C0323>=0)?1:0;

ninexnine_unit ninexnine_unit_387(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00333)
);

ninexnine_unit ninexnine_unit_388(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01333)
);

ninexnine_unit ninexnine_unit_389(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02333)
);

assign C0333=c00333+c01333+c02333;
assign A0333=(C0333>=0)?1:0;

ninexnine_unit ninexnine_unit_390(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00343)
);

ninexnine_unit ninexnine_unit_391(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01343)
);

ninexnine_unit ninexnine_unit_392(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02343)
);

assign C0343=c00343+c01343+c02343;
assign A0343=(C0343>=0)?1:0;

ninexnine_unit ninexnine_unit_393(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00353)
);

ninexnine_unit ninexnine_unit_394(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01353)
);

ninexnine_unit ninexnine_unit_395(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02353)
);

assign C0353=c00353+c01353+c02353;
assign A0353=(C0353>=0)?1:0;

ninexnine_unit ninexnine_unit_396(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00403)
);

ninexnine_unit ninexnine_unit_397(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01403)
);

ninexnine_unit ninexnine_unit_398(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02403)
);

assign C0403=c00403+c01403+c02403;
assign A0403=(C0403>=0)?1:0;

ninexnine_unit ninexnine_unit_399(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00413)
);

ninexnine_unit ninexnine_unit_400(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01413)
);

ninexnine_unit ninexnine_unit_401(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02413)
);

assign C0413=c00413+c01413+c02413;
assign A0413=(C0413>=0)?1:0;

ninexnine_unit ninexnine_unit_402(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00423)
);

ninexnine_unit ninexnine_unit_403(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01423)
);

ninexnine_unit ninexnine_unit_404(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02423)
);

assign C0423=c00423+c01423+c02423;
assign A0423=(C0423>=0)?1:0;

ninexnine_unit ninexnine_unit_405(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00433)
);

ninexnine_unit ninexnine_unit_406(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01433)
);

ninexnine_unit ninexnine_unit_407(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02433)
);

assign C0433=c00433+c01433+c02433;
assign A0433=(C0433>=0)?1:0;

ninexnine_unit ninexnine_unit_408(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00443)
);

ninexnine_unit ninexnine_unit_409(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01443)
);

ninexnine_unit ninexnine_unit_410(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02443)
);

assign C0443=c00443+c01443+c02443;
assign A0443=(C0443>=0)?1:0;

ninexnine_unit ninexnine_unit_411(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00453)
);

ninexnine_unit ninexnine_unit_412(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01453)
);

ninexnine_unit ninexnine_unit_413(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02453)
);

assign C0453=c00453+c01453+c02453;
assign A0453=(C0453>=0)?1:0;

ninexnine_unit ninexnine_unit_414(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00503)
);

ninexnine_unit ninexnine_unit_415(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01503)
);

ninexnine_unit ninexnine_unit_416(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02503)
);

assign C0503=c00503+c01503+c02503;
assign A0503=(C0503>=0)?1:0;

ninexnine_unit ninexnine_unit_417(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00513)
);

ninexnine_unit ninexnine_unit_418(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01513)
);

ninexnine_unit ninexnine_unit_419(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02513)
);

assign C0513=c00513+c01513+c02513;
assign A0513=(C0513>=0)?1:0;

ninexnine_unit ninexnine_unit_420(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00523)
);

ninexnine_unit ninexnine_unit_421(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01523)
);

ninexnine_unit ninexnine_unit_422(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02523)
);

assign C0523=c00523+c01523+c02523;
assign A0523=(C0523>=0)?1:0;

ninexnine_unit ninexnine_unit_423(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00533)
);

ninexnine_unit ninexnine_unit_424(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01533)
);

ninexnine_unit ninexnine_unit_425(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02533)
);

assign C0533=c00533+c01533+c02533;
assign A0533=(C0533>=0)?1:0;

ninexnine_unit ninexnine_unit_426(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00543)
);

ninexnine_unit ninexnine_unit_427(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01543)
);

ninexnine_unit ninexnine_unit_428(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02543)
);

assign C0543=c00543+c01543+c02543;
assign A0543=(C0543>=0)?1:0;

ninexnine_unit ninexnine_unit_429(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W03000),
				.b1(W03010),
				.b2(W03020),
				.b3(W03100),
				.b4(W03110),
				.b5(W03120),
				.b6(W03200),
				.b7(W03210),
				.b8(W03220),
				.c(c00553)
);

ninexnine_unit ninexnine_unit_430(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W03001),
				.b1(W03011),
				.b2(W03021),
				.b3(W03101),
				.b4(W03111),
				.b5(W03121),
				.b6(W03201),
				.b7(W03211),
				.b8(W03221),
				.c(c01553)
);

ninexnine_unit ninexnine_unit_431(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W03002),
				.b1(W03012),
				.b2(W03022),
				.b3(W03102),
				.b4(W03112),
				.b5(W03122),
				.b6(W03202),
				.b7(W03212),
				.b8(W03222),
				.c(c02553)
);

assign C0553=c00553+c01553+c02553;
assign A0553=(C0553>=0)?1:0;

maxpool maxpool_0(
				.clk(clk),
				.rstn(rstn),
				.a0(A0000),
				.a1(A0010),
				.a2(A0100),
				.a3(A0110),
				.p(P1110)
);

maxpool maxpool_1(
				.clk(clk),
				.rstn(rstn),
				.a0(A0020),
				.a1(A0030),
				.a2(A0120),
				.a3(A0130),
				.p(P1120)
);

maxpool maxpool_2(
				.clk(clk),
				.rstn(rstn),
				.a0(A0040),
				.a1(A0050),
				.a2(A0140),
				.a3(A0150),
				.p(P1130)
);

maxpool maxpool_3(
				.clk(clk),
				.rstn(rstn),
				.a0(A0200),
				.a1(A0210),
				.a2(A0300),
				.a3(A0310),
				.p(P1210)
);

maxpool maxpool_4(
				.clk(clk),
				.rstn(rstn),
				.a0(A0220),
				.a1(A0230),
				.a2(A0320),
				.a3(A0330),
				.p(P1220)
);

maxpool maxpool_5(
				.clk(clk),
				.rstn(rstn),
				.a0(A0240),
				.a1(A0250),
				.a2(A0340),
				.a3(A0350),
				.p(P1230)
);

maxpool maxpool_6(
				.clk(clk),
				.rstn(rstn),
				.a0(A0400),
				.a1(A0410),
				.a2(A0500),
				.a3(A0510),
				.p(P1310)
);

maxpool maxpool_7(
				.clk(clk),
				.rstn(rstn),
				.a0(A0420),
				.a1(A0430),
				.a2(A0520),
				.a3(A0530),
				.p(P1320)
);

maxpool maxpool_8(
				.clk(clk),
				.rstn(rstn),
				.a0(A0440),
				.a1(A0450),
				.a2(A0540),
				.a3(A0550),
				.p(P1330)
);

maxpool maxpool_9(
				.clk(clk),
				.rstn(rstn),
				.a0(A0001),
				.a1(A0011),
				.a2(A0101),
				.a3(A0111),
				.p(P1111)
);

maxpool maxpool_10(
				.clk(clk),
				.rstn(rstn),
				.a0(A0021),
				.a1(A0031),
				.a2(A0121),
				.a3(A0131),
				.p(P1121)
);

maxpool maxpool_11(
				.clk(clk),
				.rstn(rstn),
				.a0(A0041),
				.a1(A0051),
				.a2(A0141),
				.a3(A0151),
				.p(P1131)
);

maxpool maxpool_12(
				.clk(clk),
				.rstn(rstn),
				.a0(A0201),
				.a1(A0211),
				.a2(A0301),
				.a3(A0311),
				.p(P1211)
);

maxpool maxpool_13(
				.clk(clk),
				.rstn(rstn),
				.a0(A0221),
				.a1(A0231),
				.a2(A0321),
				.a3(A0331),
				.p(P1221)
);

maxpool maxpool_14(
				.clk(clk),
				.rstn(rstn),
				.a0(A0241),
				.a1(A0251),
				.a2(A0341),
				.a3(A0351),
				.p(P1231)
);

maxpool maxpool_15(
				.clk(clk),
				.rstn(rstn),
				.a0(A0401),
				.a1(A0411),
				.a2(A0501),
				.a3(A0511),
				.p(P1311)
);

maxpool maxpool_16(
				.clk(clk),
				.rstn(rstn),
				.a0(A0421),
				.a1(A0431),
				.a2(A0521),
				.a3(A0531),
				.p(P1321)
);

maxpool maxpool_17(
				.clk(clk),
				.rstn(rstn),
				.a0(A0441),
				.a1(A0451),
				.a2(A0541),
				.a3(A0551),
				.p(P1331)
);

maxpool maxpool_18(
				.clk(clk),
				.rstn(rstn),
				.a0(A0002),
				.a1(A0012),
				.a2(A0102),
				.a3(A0112),
				.p(P1112)
);

maxpool maxpool_19(
				.clk(clk),
				.rstn(rstn),
				.a0(A0022),
				.a1(A0032),
				.a2(A0122),
				.a3(A0132),
				.p(P1122)
);

maxpool maxpool_20(
				.clk(clk),
				.rstn(rstn),
				.a0(A0042),
				.a1(A0052),
				.a2(A0142),
				.a3(A0152),
				.p(P1132)
);

maxpool maxpool_21(
				.clk(clk),
				.rstn(rstn),
				.a0(A0202),
				.a1(A0212),
				.a2(A0302),
				.a3(A0312),
				.p(P1212)
);

maxpool maxpool_22(
				.clk(clk),
				.rstn(rstn),
				.a0(A0222),
				.a1(A0232),
				.a2(A0322),
				.a3(A0332),
				.p(P1222)
);

maxpool maxpool_23(
				.clk(clk),
				.rstn(rstn),
				.a0(A0242),
				.a1(A0252),
				.a2(A0342),
				.a3(A0352),
				.p(P1232)
);

maxpool maxpool_24(
				.clk(clk),
				.rstn(rstn),
				.a0(A0402),
				.a1(A0412),
				.a2(A0502),
				.a3(A0512),
				.p(P1312)
);

maxpool maxpool_25(
				.clk(clk),
				.rstn(rstn),
				.a0(A0422),
				.a1(A0432),
				.a2(A0522),
				.a3(A0532),
				.p(P1322)
);

maxpool maxpool_26(
				.clk(clk),
				.rstn(rstn),
				.a0(A0442),
				.a1(A0452),
				.a2(A0542),
				.a3(A0552),
				.p(P1332)
);

maxpool maxpool_27(
				.clk(clk),
				.rstn(rstn),
				.a0(A0003),
				.a1(A0013),
				.a2(A0103),
				.a3(A0113),
				.p(P1113)
);

maxpool maxpool_28(
				.clk(clk),
				.rstn(rstn),
				.a0(A0023),
				.a1(A0033),
				.a2(A0123),
				.a3(A0133),
				.p(P1123)
);

maxpool maxpool_29(
				.clk(clk),
				.rstn(rstn),
				.a0(A0043),
				.a1(A0053),
				.a2(A0143),
				.a3(A0153),
				.p(P1133)
);

maxpool maxpool_30(
				.clk(clk),
				.rstn(rstn),
				.a0(A0203),
				.a1(A0213),
				.a2(A0303),
				.a3(A0313),
				.p(P1213)
);

maxpool maxpool_31(
				.clk(clk),
				.rstn(rstn),
				.a0(A0223),
				.a1(A0233),
				.a2(A0323),
				.a3(A0333),
				.p(P1223)
);

maxpool maxpool_32(
				.clk(clk),
				.rstn(rstn),
				.a0(A0243),
				.a1(A0253),
				.a2(A0343),
				.a3(A0353),
				.p(P1233)
);

maxpool maxpool_33(
				.clk(clk),
				.rstn(rstn),
				.a0(A0403),
				.a1(A0413),
				.a2(A0503),
				.a3(A0513),
				.p(P1313)
);

maxpool maxpool_34(
				.clk(clk),
				.rstn(rstn),
				.a0(A0423),
				.a1(A0433),
				.a2(A0523),
				.a3(A0533),
				.p(P1323)
);

maxpool maxpool_35(
				.clk(clk),
				.rstn(rstn),
				.a0(A0443),
				.a1(A0453),
				.a2(A0543),
				.a3(A0553),
				.p(P1333)
);

//layer0 done, begain next layer
(*DONT_TOUCH="true"*) wire P1000;
(*DONT_TOUCH="true"*) wire P1010;
(*DONT_TOUCH="true"*) wire P1020;
(*DONT_TOUCH="true"*) wire P1030;
(*DONT_TOUCH="true"*) wire P1100;
(*DONT_TOUCH="true"*) wire P1200;
(*DONT_TOUCH="true"*) wire P1300;
(*DONT_TOUCH="true"*) wire P1001;
(*DONT_TOUCH="true"*) wire P1011;
(*DONT_TOUCH="true"*) wire P1021;
(*DONT_TOUCH="true"*) wire P1031;
(*DONT_TOUCH="true"*) wire P1101;
(*DONT_TOUCH="true"*) wire P1201;
(*DONT_TOUCH="true"*) wire P1301;
(*DONT_TOUCH="true"*) wire P1002;
(*DONT_TOUCH="true"*) wire P1012;
(*DONT_TOUCH="true"*) wire P1022;
(*DONT_TOUCH="true"*) wire P1032;
(*DONT_TOUCH="true"*) wire P1102;
(*DONT_TOUCH="true"*) wire P1202;
(*DONT_TOUCH="true"*) wire P1302;
(*DONT_TOUCH="true"*) wire P1003;
(*DONT_TOUCH="true"*) wire P1013;
(*DONT_TOUCH="true"*) wire P1023;
(*DONT_TOUCH="true"*) wire P1033;
(*DONT_TOUCH="true"*) wire P1103;
(*DONT_TOUCH="true"*) wire P1203;
(*DONT_TOUCH="true"*) wire P1303;
(*DONT_TOUCH="true"*) wire P2000;
(*DONT_TOUCH="true"*) wire W10000,W10010,W10020,W10100,W10110,W10120,W10200,W10210,W10220;
(*DONT_TOUCH="true"*) wire W10001,W10011,W10021,W10101,W10111,W10121,W10201,W10211,W10221;
(*DONT_TOUCH="true"*) wire W10002,W10012,W10022,W10102,W10112,W10122,W10202,W10212,W10222;
(*DONT_TOUCH="true"*) wire W10003,W10013,W10023,W10103,W10113,W10123,W10203,W10213,W10223;
(*DONT_TOUCH="true"*) wire signed [4:0] c10000,c11000,c12000,c13000;
(*DONT_TOUCH="true"*) wire signed [4:0] c10010,c11010,c12010,c13010;
(*DONT_TOUCH="true"*) wire signed [4:0] c10020,c11020,c12020,c13020;
(*DONT_TOUCH="true"*) wire signed [4:0] c10100,c11100,c12100,c13100;
(*DONT_TOUCH="true"*) wire signed [4:0] c10110,c11110,c12110,c13110;
(*DONT_TOUCH="true"*) wire signed [4:0] c10120,c11120,c12120,c13120;
(*DONT_TOUCH="true"*) wire signed [4:0] c10200,c11200,c12200,c13200;
(*DONT_TOUCH="true"*) wire signed [4:0] c10210,c11210,c12210,c13210;
(*DONT_TOUCH="true"*) wire signed [4:0] c10220,c11220,c12220,c13220;
(*DONT_TOUCH="true"*) wire signed [6:0] C1000;
(*DONT_TOUCH="true"*) wire A1000;
(*DONT_TOUCH="true"*) wire signed [6:0] C1010;
(*DONT_TOUCH="true"*) wire A1010;
(*DONT_TOUCH="true"*) wire signed [6:0] C1100;
(*DONT_TOUCH="true"*) wire A1100;
(*DONT_TOUCH="true"*) wire signed [6:0] C1110;
(*DONT_TOUCH="true"*) wire A1110;
DFF_save_fm DFF_P192(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1000));
DFF_save_fm DFF_P193(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1010));
DFF_save_fm DFF_P194(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1020));
DFF_save_fm DFF_P195(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1030));
DFF_save_fm DFF_P196(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1100));
DFF_save_fm DFF_P197(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1200));
DFF_save_fm DFF_P198(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1300));
DFF_save_fm DFF_P199(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1001));
DFF_save_fm DFF_P200(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1011));
DFF_save_fm DFF_P201(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1021));
DFF_save_fm DFF_P202(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1031));
DFF_save_fm DFF_P203(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1101));
DFF_save_fm DFF_P204(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1201));
DFF_save_fm DFF_P205(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1301));
DFF_save_fm DFF_P206(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1002));
DFF_save_fm DFF_P207(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1012));
DFF_save_fm DFF_P208(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1022));
DFF_save_fm DFF_P209(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1032));
DFF_save_fm DFF_P210(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1102));
DFF_save_fm DFF_P211(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1202));
DFF_save_fm DFF_P212(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1302));
DFF_save_fm DFF_P213(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1003));
DFF_save_fm DFF_P214(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1013));
DFF_save_fm DFF_P215(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1023));
DFF_save_fm DFF_P216(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1033));
DFF_save_fm DFF_P217(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1103));
DFF_save_fm DFF_P218(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1203));
DFF_save_fm DFF_P219(.clk(clk),.rstn(rstn),.reset_value(1),.q(P1303));
DFF_save_fm DFF_W108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10000));
DFF_save_fm DFF_W109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10010));
DFF_save_fm DFF_W110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10020));
DFF_save_fm DFF_W111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10100));
DFF_save_fm DFF_W112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10110));
DFF_save_fm DFF_W113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10120));
DFF_save_fm DFF_W114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10200));
DFF_save_fm DFF_W115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10210));
DFF_save_fm DFF_W116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10220));
DFF_save_fm DFF_W117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10001));
DFF_save_fm DFF_W118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10011));
DFF_save_fm DFF_W119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10021));
DFF_save_fm DFF_W120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10101));
DFF_save_fm DFF_W121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10111));
DFF_save_fm DFF_W122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10121));
DFF_save_fm DFF_W123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10201));
DFF_save_fm DFF_W124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10211));
DFF_save_fm DFF_W125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10221));
DFF_save_fm DFF_W126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10002));
DFF_save_fm DFF_W127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10012));
DFF_save_fm DFF_W128(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10022));
DFF_save_fm DFF_W129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10102));
DFF_save_fm DFF_W130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10112));
DFF_save_fm DFF_W131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10122));
DFF_save_fm DFF_W132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10202));
DFF_save_fm DFF_W133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10212));
DFF_save_fm DFF_W134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10222));
DFF_save_fm DFF_W135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10003));
DFF_save_fm DFF_W136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10013));
DFF_save_fm DFF_W137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10023));
DFF_save_fm DFF_W138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10103));
DFF_save_fm DFF_W139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10113));
DFF_save_fm DFF_W140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10123));
DFF_save_fm DFF_W141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10203));
DFF_save_fm DFF_W142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10213));
DFF_save_fm DFF_W143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10223));
ninexnine_unit ninexnine_unit_432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10000)
);

ninexnine_unit ninexnine_unit_433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11000)
);

ninexnine_unit ninexnine_unit_434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12000)
);

ninexnine_unit ninexnine_unit_435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1003),
				.a1(P1013),
				.a2(P1023),
				.a3(P1103),
				.a4(P1113),
				.a5(P1123),
				.a6(P1203),
				.a7(P1213),
				.a8(P1223),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13000)
);

assign C1000=c10000+c11000+c12000+c13000;
assign A1000=(C1000>=0)?1:0;

ninexnine_unit ninexnine_unit_436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10010)
);

ninexnine_unit ninexnine_unit_437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11010)
);

ninexnine_unit ninexnine_unit_438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12010)
);

ninexnine_unit ninexnine_unit_439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1013),
				.a1(P1023),
				.a2(P1033),
				.a3(P1113),
				.a4(P1123),
				.a5(P1133),
				.a6(P1213),
				.a7(P1223),
				.a8(P1233),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13010)
);

assign C1010=c10010+c11010+c12010+c13010;
assign A1010=(C1010>=0)?1:0;

ninexnine_unit ninexnine_unit_440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10100)
);

ninexnine_unit ninexnine_unit_441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11100)
);

ninexnine_unit ninexnine_unit_442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12100)
);

ninexnine_unit ninexnine_unit_443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1103),
				.a1(P1113),
				.a2(P1123),
				.a3(P1203),
				.a4(P1213),
				.a5(P1223),
				.a6(P1303),
				.a7(P1313),
				.a8(P1323),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13100)
);

assign C1100=c10100+c11100+c12100+c13100;
assign A1100=(C1100>=0)?1:0;

ninexnine_unit ninexnine_unit_444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10110)
);

ninexnine_unit ninexnine_unit_445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11110)
);

ninexnine_unit ninexnine_unit_446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12110)
);

ninexnine_unit ninexnine_unit_447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1113),
				.a1(P1123),
				.a2(P1133),
				.a3(P1213),
				.a4(P1223),
				.a5(P1233),
				.a6(P1313),
				.a7(P1323),
				.a8(P1333),
				.b0(W10003),
				.b1(W10013),
				.b2(W10023),
				.b3(W10103),
				.b4(W10113),
				.b5(W10123),
				.b6(W10203),
				.b7(W10213),
				.b8(W10223),
				.c(c13110)
);

assign C1110=c10110+c11110+c12110+c13110;
assign A1110=(C1110>=0)?1:0;

maxpool maxpool_36(
				.clk(clk),
				.rstn(rstn),
				.a0(A1000),
				.a1(A1010),
				.a2(A1100),
				.a3(A1110),
				.p(P2000)
);

//layer1 done, begain next layer
