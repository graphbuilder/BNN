module tb_test_layer2(

);
reg clk,rstn;
test_layer2 test_layer2(
clk,
rstn
);
reg mem[14*14*4-1:0];
always #5 clk=~clk;
initial
begin
clk=0;
rstn=0;
$readmemb("D:/work/PROJ_5/proj_2/src/to_csma/test_tb/answer_layer_2.txt",mem);
#10;
rstn=1;
end
reg [31:0]count;
always@(posedge clk or negedge rstn)
	if(~rstn)
		count<=0;
	else
		count<=count+1;

reg Pass_0;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_0<=0;
	else if(count>=2)
		begin
			if(tb_test_layer2.test_layer2.P3000==mem[0])
				Pass_0<=1;
			else
				Pass_0<=0;
		end

reg Pass_1;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_1<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3010==mem[1])&&(Pass_0))
				Pass_1<=1;
			else
				Pass_1<=0;
		end

reg Pass_2;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_2<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3020==mem[2])&&(Pass_1))
				Pass_2<=1;
			else
				Pass_2<=0;
		end

reg Pass_3;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_3<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3030==mem[3])&&(Pass_2))
				Pass_3<=1;
			else
				Pass_3<=0;
		end

reg Pass_4;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_4<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3040==mem[4])&&(Pass_3))
				Pass_4<=1;
			else
				Pass_4<=0;
		end

reg Pass_5;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_5<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3100==mem[5])&&(Pass_4))
				Pass_5<=1;
			else
				Pass_5<=0;
		end

reg Pass_6;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_6<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3110==mem[6])&&(Pass_5))
				Pass_6<=1;
			else
				Pass_6<=0;
		end

reg Pass_7;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_7<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3120==mem[7])&&(Pass_6))
				Pass_7<=1;
			else
				Pass_7<=0;
		end

reg Pass_8;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_8<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3130==mem[8])&&(Pass_7))
				Pass_8<=1;
			else
				Pass_8<=0;
		end

reg Pass_9;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_9<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3140==mem[9])&&(Pass_8))
				Pass_9<=1;
			else
				Pass_9<=0;
		end

reg Pass_10;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_10<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3200==mem[10])&&(Pass_9))
				Pass_10<=1;
			else
				Pass_10<=0;
		end

reg Pass_11;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_11<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3210==mem[11])&&(Pass_10))
				Pass_11<=1;
			else
				Pass_11<=0;
		end

reg Pass_12;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_12<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3220==mem[12])&&(Pass_11))
				Pass_12<=1;
			else
				Pass_12<=0;
		end

reg Pass_13;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_13<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3230==mem[13])&&(Pass_12))
				Pass_13<=1;
			else
				Pass_13<=0;
		end

reg Pass_14;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_14<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3240==mem[14])&&(Pass_13))
				Pass_14<=1;
			else
				Pass_14<=0;
		end

reg Pass_15;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_15<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3300==mem[15])&&(Pass_14))
				Pass_15<=1;
			else
				Pass_15<=0;
		end

reg Pass_16;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_16<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3310==mem[16])&&(Pass_15))
				Pass_16<=1;
			else
				Pass_16<=0;
		end

reg Pass_17;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_17<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3320==mem[17])&&(Pass_16))
				Pass_17<=1;
			else
				Pass_17<=0;
		end

reg Pass_18;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_18<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3330==mem[18])&&(Pass_17))
				Pass_18<=1;
			else
				Pass_18<=0;
		end

reg Pass_19;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_19<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3340==mem[19])&&(Pass_18))
				Pass_19<=1;
			else
				Pass_19<=0;
		end

reg Pass_20;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_20<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3400==mem[20])&&(Pass_19))
				Pass_20<=1;
			else
				Pass_20<=0;
		end

reg Pass_21;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_21<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3410==mem[21])&&(Pass_20))
				Pass_21<=1;
			else
				Pass_21<=0;
		end

reg Pass_22;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_22<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3420==mem[22])&&(Pass_21))
				Pass_22<=1;
			else
				Pass_22<=0;
		end

reg Pass_23;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_23<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3430==mem[23])&&(Pass_22))
				Pass_23<=1;
			else
				Pass_23<=0;
		end

reg Pass_24;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_24<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3440==mem[24])&&(Pass_23))
				Pass_24<=1;
			else
				Pass_24<=0;
		end

reg Pass_25;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_25<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3001==mem[25])&&(Pass_24))
				Pass_25<=1;
			else
				Pass_25<=0;
		end

reg Pass_26;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_26<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3011==mem[26])&&(Pass_25))
				Pass_26<=1;
			else
				Pass_26<=0;
		end

reg Pass_27;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_27<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3021==mem[27])&&(Pass_26))
				Pass_27<=1;
			else
				Pass_27<=0;
		end

reg Pass_28;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_28<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3031==mem[28])&&(Pass_27))
				Pass_28<=1;
			else
				Pass_28<=0;
		end

reg Pass_29;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_29<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3041==mem[29])&&(Pass_28))
				Pass_29<=1;
			else
				Pass_29<=0;
		end

reg Pass_30;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_30<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3101==mem[30])&&(Pass_29))
				Pass_30<=1;
			else
				Pass_30<=0;
		end

reg Pass_31;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_31<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3111==mem[31])&&(Pass_30))
				Pass_31<=1;
			else
				Pass_31<=0;
		end

reg Pass_32;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_32<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3121==mem[32])&&(Pass_31))
				Pass_32<=1;
			else
				Pass_32<=0;
		end

reg Pass_33;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_33<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3131==mem[33])&&(Pass_32))
				Pass_33<=1;
			else
				Pass_33<=0;
		end

reg Pass_34;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_34<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3141==mem[34])&&(Pass_33))
				Pass_34<=1;
			else
				Pass_34<=0;
		end

reg Pass_35;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_35<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3201==mem[35])&&(Pass_34))
				Pass_35<=1;
			else
				Pass_35<=0;
		end

reg Pass_36;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_36<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3211==mem[36])&&(Pass_35))
				Pass_36<=1;
			else
				Pass_36<=0;
		end

reg Pass_37;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_37<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3221==mem[37])&&(Pass_36))
				Pass_37<=1;
			else
				Pass_37<=0;
		end

reg Pass_38;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_38<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3231==mem[38])&&(Pass_37))
				Pass_38<=1;
			else
				Pass_38<=0;
		end

reg Pass_39;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_39<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3241==mem[39])&&(Pass_38))
				Pass_39<=1;
			else
				Pass_39<=0;
		end

reg Pass_40;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_40<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3301==mem[40])&&(Pass_39))
				Pass_40<=1;
			else
				Pass_40<=0;
		end

reg Pass_41;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_41<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3311==mem[41])&&(Pass_40))
				Pass_41<=1;
			else
				Pass_41<=0;
		end

reg Pass_42;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_42<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3321==mem[42])&&(Pass_41))
				Pass_42<=1;
			else
				Pass_42<=0;
		end

reg Pass_43;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_43<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3331==mem[43])&&(Pass_42))
				Pass_43<=1;
			else
				Pass_43<=0;
		end

reg Pass_44;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_44<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3341==mem[44])&&(Pass_43))
				Pass_44<=1;
			else
				Pass_44<=0;
		end

reg Pass_45;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_45<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3401==mem[45])&&(Pass_44))
				Pass_45<=1;
			else
				Pass_45<=0;
		end

reg Pass_46;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_46<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3411==mem[46])&&(Pass_45))
				Pass_46<=1;
			else
				Pass_46<=0;
		end

reg Pass_47;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_47<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3421==mem[47])&&(Pass_46))
				Pass_47<=1;
			else
				Pass_47<=0;
		end

reg Pass_48;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_48<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3431==mem[48])&&(Pass_47))
				Pass_48<=1;
			else
				Pass_48<=0;
		end

reg Pass_49;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_49<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3441==mem[49])&&(Pass_48))
				Pass_49<=1;
			else
				Pass_49<=0;
		end

reg Pass_50;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_50<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3002==mem[50])&&(Pass_49))
				Pass_50<=1;
			else
				Pass_50<=0;
		end

reg Pass_51;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_51<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3012==mem[51])&&(Pass_50))
				Pass_51<=1;
			else
				Pass_51<=0;
		end

reg Pass_52;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_52<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3022==mem[52])&&(Pass_51))
				Pass_52<=1;
			else
				Pass_52<=0;
		end

reg Pass_53;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_53<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3032==mem[53])&&(Pass_52))
				Pass_53<=1;
			else
				Pass_53<=0;
		end

reg Pass_54;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_54<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3042==mem[54])&&(Pass_53))
				Pass_54<=1;
			else
				Pass_54<=0;
		end

reg Pass_55;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_55<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3102==mem[55])&&(Pass_54))
				Pass_55<=1;
			else
				Pass_55<=0;
		end

reg Pass_56;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_56<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3112==mem[56])&&(Pass_55))
				Pass_56<=1;
			else
				Pass_56<=0;
		end

reg Pass_57;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_57<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3122==mem[57])&&(Pass_56))
				Pass_57<=1;
			else
				Pass_57<=0;
		end

reg Pass_58;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_58<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3132==mem[58])&&(Pass_57))
				Pass_58<=1;
			else
				Pass_58<=0;
		end

reg Pass_59;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_59<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3142==mem[59])&&(Pass_58))
				Pass_59<=1;
			else
				Pass_59<=0;
		end

reg Pass_60;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_60<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3202==mem[60])&&(Pass_59))
				Pass_60<=1;
			else
				Pass_60<=0;
		end

reg Pass_61;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_61<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3212==mem[61])&&(Pass_60))
				Pass_61<=1;
			else
				Pass_61<=0;
		end

reg Pass_62;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_62<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3222==mem[62])&&(Pass_61))
				Pass_62<=1;
			else
				Pass_62<=0;
		end

reg Pass_63;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_63<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3232==mem[63])&&(Pass_62))
				Pass_63<=1;
			else
				Pass_63<=0;
		end

reg Pass_64;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_64<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3242==mem[64])&&(Pass_63))
				Pass_64<=1;
			else
				Pass_64<=0;
		end

reg Pass_65;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_65<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3302==mem[65])&&(Pass_64))
				Pass_65<=1;
			else
				Pass_65<=0;
		end

reg Pass_66;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_66<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3312==mem[66])&&(Pass_65))
				Pass_66<=1;
			else
				Pass_66<=0;
		end

reg Pass_67;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_67<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3322==mem[67])&&(Pass_66))
				Pass_67<=1;
			else
				Pass_67<=0;
		end

reg Pass_68;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_68<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3332==mem[68])&&(Pass_67))
				Pass_68<=1;
			else
				Pass_68<=0;
		end

reg Pass_69;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_69<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3342==mem[69])&&(Pass_68))
				Pass_69<=1;
			else
				Pass_69<=0;
		end

reg Pass_70;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_70<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3402==mem[70])&&(Pass_69))
				Pass_70<=1;
			else
				Pass_70<=0;
		end

reg Pass_71;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_71<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3412==mem[71])&&(Pass_70))
				Pass_71<=1;
			else
				Pass_71<=0;
		end

reg Pass_72;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_72<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3422==mem[72])&&(Pass_71))
				Pass_72<=1;
			else
				Pass_72<=0;
		end

reg Pass_73;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_73<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3432==mem[73])&&(Pass_72))
				Pass_73<=1;
			else
				Pass_73<=0;
		end

reg Pass_74;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_74<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3442==mem[74])&&(Pass_73))
				Pass_74<=1;
			else
				Pass_74<=0;
		end

reg Pass_75;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_75<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3003==mem[75])&&(Pass_74))
				Pass_75<=1;
			else
				Pass_75<=0;
		end

reg Pass_76;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_76<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3013==mem[76])&&(Pass_75))
				Pass_76<=1;
			else
				Pass_76<=0;
		end

reg Pass_77;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_77<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3023==mem[77])&&(Pass_76))
				Pass_77<=1;
			else
				Pass_77<=0;
		end

reg Pass_78;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_78<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3033==mem[78])&&(Pass_77))
				Pass_78<=1;
			else
				Pass_78<=0;
		end

reg Pass_79;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_79<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3043==mem[79])&&(Pass_78))
				Pass_79<=1;
			else
				Pass_79<=0;
		end

reg Pass_80;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_80<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3103==mem[80])&&(Pass_79))
				Pass_80<=1;
			else
				Pass_80<=0;
		end

reg Pass_81;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_81<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3113==mem[81])&&(Pass_80))
				Pass_81<=1;
			else
				Pass_81<=0;
		end

reg Pass_82;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_82<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3123==mem[82])&&(Pass_81))
				Pass_82<=1;
			else
				Pass_82<=0;
		end

reg Pass_83;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_83<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3133==mem[83])&&(Pass_82))
				Pass_83<=1;
			else
				Pass_83<=0;
		end

reg Pass_84;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_84<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3143==mem[84])&&(Pass_83))
				Pass_84<=1;
			else
				Pass_84<=0;
		end

reg Pass_85;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_85<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3203==mem[85])&&(Pass_84))
				Pass_85<=1;
			else
				Pass_85<=0;
		end

reg Pass_86;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_86<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3213==mem[86])&&(Pass_85))
				Pass_86<=1;
			else
				Pass_86<=0;
		end

reg Pass_87;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_87<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3223==mem[87])&&(Pass_86))
				Pass_87<=1;
			else
				Pass_87<=0;
		end

reg Pass_88;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_88<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3233==mem[88])&&(Pass_87))
				Pass_88<=1;
			else
				Pass_88<=0;
		end

reg Pass_89;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_89<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3243==mem[89])&&(Pass_88))
				Pass_89<=1;
			else
				Pass_89<=0;
		end

reg Pass_90;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_90<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3303==mem[90])&&(Pass_89))
				Pass_90<=1;
			else
				Pass_90<=0;
		end

reg Pass_91;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_91<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3313==mem[91])&&(Pass_90))
				Pass_91<=1;
			else
				Pass_91<=0;
		end

reg Pass_92;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_92<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3323==mem[92])&&(Pass_91))
				Pass_92<=1;
			else
				Pass_92<=0;
		end

reg Pass_93;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_93<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3333==mem[93])&&(Pass_92))
				Pass_93<=1;
			else
				Pass_93<=0;
		end

reg Pass_94;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_94<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3343==mem[94])&&(Pass_93))
				Pass_94<=1;
			else
				Pass_94<=0;
		end

reg Pass_95;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_95<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3403==mem[95])&&(Pass_94))
				Pass_95<=1;
			else
				Pass_95<=0;
		end

reg Pass_96;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_96<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3413==mem[96])&&(Pass_95))
				Pass_96<=1;
			else
				Pass_96<=0;
		end

reg Pass_97;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_97<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3423==mem[97])&&(Pass_96))
				Pass_97<=1;
			else
				Pass_97<=0;
		end

reg Pass_98;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_98<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3433==mem[98])&&(Pass_97))
				Pass_98<=1;
			else
				Pass_98<=0;
		end

reg Pass_99;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_99<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3443==mem[99])&&(Pass_98))
				Pass_99<=1;
			else
				Pass_99<=0;
		end

reg Pass_100;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_100<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3004==mem[100])&&(Pass_99))
				Pass_100<=1;
			else
				Pass_100<=0;
		end

reg Pass_101;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_101<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3014==mem[101])&&(Pass_100))
				Pass_101<=1;
			else
				Pass_101<=0;
		end

reg Pass_102;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_102<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3024==mem[102])&&(Pass_101))
				Pass_102<=1;
			else
				Pass_102<=0;
		end

reg Pass_103;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_103<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3034==mem[103])&&(Pass_102))
				Pass_103<=1;
			else
				Pass_103<=0;
		end

reg Pass_104;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_104<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3044==mem[104])&&(Pass_103))
				Pass_104<=1;
			else
				Pass_104<=0;
		end

reg Pass_105;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_105<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3104==mem[105])&&(Pass_104))
				Pass_105<=1;
			else
				Pass_105<=0;
		end

reg Pass_106;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_106<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3114==mem[106])&&(Pass_105))
				Pass_106<=1;
			else
				Pass_106<=0;
		end

reg Pass_107;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_107<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3124==mem[107])&&(Pass_106))
				Pass_107<=1;
			else
				Pass_107<=0;
		end

reg Pass_108;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_108<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3134==mem[108])&&(Pass_107))
				Pass_108<=1;
			else
				Pass_108<=0;
		end

reg Pass_109;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_109<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3144==mem[109])&&(Pass_108))
				Pass_109<=1;
			else
				Pass_109<=0;
		end

reg Pass_110;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_110<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3204==mem[110])&&(Pass_109))
				Pass_110<=1;
			else
				Pass_110<=0;
		end

reg Pass_111;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_111<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3214==mem[111])&&(Pass_110))
				Pass_111<=1;
			else
				Pass_111<=0;
		end

reg Pass_112;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_112<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3224==mem[112])&&(Pass_111))
				Pass_112<=1;
			else
				Pass_112<=0;
		end

reg Pass_113;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_113<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3234==mem[113])&&(Pass_112))
				Pass_113<=1;
			else
				Pass_113<=0;
		end

reg Pass_114;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_114<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3244==mem[114])&&(Pass_113))
				Pass_114<=1;
			else
				Pass_114<=0;
		end

reg Pass_115;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_115<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3304==mem[115])&&(Pass_114))
				Pass_115<=1;
			else
				Pass_115<=0;
		end

reg Pass_116;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_116<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3314==mem[116])&&(Pass_115))
				Pass_116<=1;
			else
				Pass_116<=0;
		end

reg Pass_117;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_117<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3324==mem[117])&&(Pass_116))
				Pass_117<=1;
			else
				Pass_117<=0;
		end

reg Pass_118;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_118<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3334==mem[118])&&(Pass_117))
				Pass_118<=1;
			else
				Pass_118<=0;
		end

reg Pass_119;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_119<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3344==mem[119])&&(Pass_118))
				Pass_119<=1;
			else
				Pass_119<=0;
		end

reg Pass_120;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_120<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3404==mem[120])&&(Pass_119))
				Pass_120<=1;
			else
				Pass_120<=0;
		end

reg Pass_121;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_121<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3414==mem[121])&&(Pass_120))
				Pass_121<=1;
			else
				Pass_121<=0;
		end

reg Pass_122;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_122<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3424==mem[122])&&(Pass_121))
				Pass_122<=1;
			else
				Pass_122<=0;
		end

reg Pass_123;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_123<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3434==mem[123])&&(Pass_122))
				Pass_123<=1;
			else
				Pass_123<=0;
		end

reg Pass_124;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_124<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3444==mem[124])&&(Pass_123))
				Pass_124<=1;
			else
				Pass_124<=0;
		end

reg Pass_125;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_125<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3005==mem[125])&&(Pass_124))
				Pass_125<=1;
			else
				Pass_125<=0;
		end

reg Pass_126;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_126<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3015==mem[126])&&(Pass_125))
				Pass_126<=1;
			else
				Pass_126<=0;
		end

reg Pass_127;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_127<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3025==mem[127])&&(Pass_126))
				Pass_127<=1;
			else
				Pass_127<=0;
		end

reg Pass_128;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_128<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3035==mem[128])&&(Pass_127))
				Pass_128<=1;
			else
				Pass_128<=0;
		end

reg Pass_129;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_129<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3045==mem[129])&&(Pass_128))
				Pass_129<=1;
			else
				Pass_129<=0;
		end

reg Pass_130;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_130<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3105==mem[130])&&(Pass_129))
				Pass_130<=1;
			else
				Pass_130<=0;
		end

reg Pass_131;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_131<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3115==mem[131])&&(Pass_130))
				Pass_131<=1;
			else
				Pass_131<=0;
		end

reg Pass_132;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_132<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3125==mem[132])&&(Pass_131))
				Pass_132<=1;
			else
				Pass_132<=0;
		end

reg Pass_133;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_133<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3135==mem[133])&&(Pass_132))
				Pass_133<=1;
			else
				Pass_133<=0;
		end

reg Pass_134;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_134<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3145==mem[134])&&(Pass_133))
				Pass_134<=1;
			else
				Pass_134<=0;
		end

reg Pass_135;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_135<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3205==mem[135])&&(Pass_134))
				Pass_135<=1;
			else
				Pass_135<=0;
		end

reg Pass_136;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_136<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3215==mem[136])&&(Pass_135))
				Pass_136<=1;
			else
				Pass_136<=0;
		end

reg Pass_137;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_137<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3225==mem[137])&&(Pass_136))
				Pass_137<=1;
			else
				Pass_137<=0;
		end

reg Pass_138;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_138<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3235==mem[138])&&(Pass_137))
				Pass_138<=1;
			else
				Pass_138<=0;
		end

reg Pass_139;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_139<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3245==mem[139])&&(Pass_138))
				Pass_139<=1;
			else
				Pass_139<=0;
		end

reg Pass_140;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_140<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3305==mem[140])&&(Pass_139))
				Pass_140<=1;
			else
				Pass_140<=0;
		end

reg Pass_141;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_141<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3315==mem[141])&&(Pass_140))
				Pass_141<=1;
			else
				Pass_141<=0;
		end

reg Pass_142;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_142<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3325==mem[142])&&(Pass_141))
				Pass_142<=1;
			else
				Pass_142<=0;
		end

reg Pass_143;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_143<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3335==mem[143])&&(Pass_142))
				Pass_143<=1;
			else
				Pass_143<=0;
		end

reg Pass_144;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_144<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3345==mem[144])&&(Pass_143))
				Pass_144<=1;
			else
				Pass_144<=0;
		end

reg Pass_145;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_145<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3405==mem[145])&&(Pass_144))
				Pass_145<=1;
			else
				Pass_145<=0;
		end

reg Pass_146;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_146<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3415==mem[146])&&(Pass_145))
				Pass_146<=1;
			else
				Pass_146<=0;
		end

reg Pass_147;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_147<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3425==mem[147])&&(Pass_146))
				Pass_147<=1;
			else
				Pass_147<=0;
		end

reg Pass_148;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_148<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3435==mem[148])&&(Pass_147))
				Pass_148<=1;
			else
				Pass_148<=0;
		end

reg Pass_149;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_149<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3445==mem[149])&&(Pass_148))
				Pass_149<=1;
			else
				Pass_149<=0;
		end

reg Pass_150;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_150<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3006==mem[150])&&(Pass_149))
				Pass_150<=1;
			else
				Pass_150<=0;
		end

reg Pass_151;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_151<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3016==mem[151])&&(Pass_150))
				Pass_151<=1;
			else
				Pass_151<=0;
		end

reg Pass_152;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_152<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3026==mem[152])&&(Pass_151))
				Pass_152<=1;
			else
				Pass_152<=0;
		end

reg Pass_153;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_153<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3036==mem[153])&&(Pass_152))
				Pass_153<=1;
			else
				Pass_153<=0;
		end

reg Pass_154;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_154<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3046==mem[154])&&(Pass_153))
				Pass_154<=1;
			else
				Pass_154<=0;
		end

reg Pass_155;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_155<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3106==mem[155])&&(Pass_154))
				Pass_155<=1;
			else
				Pass_155<=0;
		end

reg Pass_156;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_156<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3116==mem[156])&&(Pass_155))
				Pass_156<=1;
			else
				Pass_156<=0;
		end

reg Pass_157;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_157<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3126==mem[157])&&(Pass_156))
				Pass_157<=1;
			else
				Pass_157<=0;
		end

reg Pass_158;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_158<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3136==mem[158])&&(Pass_157))
				Pass_158<=1;
			else
				Pass_158<=0;
		end

reg Pass_159;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_159<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3146==mem[159])&&(Pass_158))
				Pass_159<=1;
			else
				Pass_159<=0;
		end

reg Pass_160;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_160<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3206==mem[160])&&(Pass_159))
				Pass_160<=1;
			else
				Pass_160<=0;
		end

reg Pass_161;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_161<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3216==mem[161])&&(Pass_160))
				Pass_161<=1;
			else
				Pass_161<=0;
		end

reg Pass_162;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_162<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3226==mem[162])&&(Pass_161))
				Pass_162<=1;
			else
				Pass_162<=0;
		end

reg Pass_163;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_163<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3236==mem[163])&&(Pass_162))
				Pass_163<=1;
			else
				Pass_163<=0;
		end

reg Pass_164;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_164<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3246==mem[164])&&(Pass_163))
				Pass_164<=1;
			else
				Pass_164<=0;
		end

reg Pass_165;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_165<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3306==mem[165])&&(Pass_164))
				Pass_165<=1;
			else
				Pass_165<=0;
		end

reg Pass_166;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_166<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3316==mem[166])&&(Pass_165))
				Pass_166<=1;
			else
				Pass_166<=0;
		end

reg Pass_167;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_167<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3326==mem[167])&&(Pass_166))
				Pass_167<=1;
			else
				Pass_167<=0;
		end

reg Pass_168;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_168<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3336==mem[168])&&(Pass_167))
				Pass_168<=1;
			else
				Pass_168<=0;
		end

reg Pass_169;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_169<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3346==mem[169])&&(Pass_168))
				Pass_169<=1;
			else
				Pass_169<=0;
		end

reg Pass_170;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_170<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3406==mem[170])&&(Pass_169))
				Pass_170<=1;
			else
				Pass_170<=0;
		end

reg Pass_171;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_171<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3416==mem[171])&&(Pass_170))
				Pass_171<=1;
			else
				Pass_171<=0;
		end

reg Pass_172;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_172<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3426==mem[172])&&(Pass_171))
				Pass_172<=1;
			else
				Pass_172<=0;
		end

reg Pass_173;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_173<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3436==mem[173])&&(Pass_172))
				Pass_173<=1;
			else
				Pass_173<=0;
		end

reg Pass_174;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_174<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3446==mem[174])&&(Pass_173))
				Pass_174<=1;
			else
				Pass_174<=0;
		end

reg Pass_175;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_175<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3007==mem[175])&&(Pass_174))
				Pass_175<=1;
			else
				Pass_175<=0;
		end

reg Pass_176;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_176<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3017==mem[176])&&(Pass_175))
				Pass_176<=1;
			else
				Pass_176<=0;
		end

reg Pass_177;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_177<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3027==mem[177])&&(Pass_176))
				Pass_177<=1;
			else
				Pass_177<=0;
		end

reg Pass_178;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_178<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3037==mem[178])&&(Pass_177))
				Pass_178<=1;
			else
				Pass_178<=0;
		end

reg Pass_179;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_179<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3047==mem[179])&&(Pass_178))
				Pass_179<=1;
			else
				Pass_179<=0;
		end

reg Pass_180;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_180<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3107==mem[180])&&(Pass_179))
				Pass_180<=1;
			else
				Pass_180<=0;
		end

reg Pass_181;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_181<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3117==mem[181])&&(Pass_180))
				Pass_181<=1;
			else
				Pass_181<=0;
		end

reg Pass_182;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_182<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3127==mem[182])&&(Pass_181))
				Pass_182<=1;
			else
				Pass_182<=0;
		end

reg Pass_183;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_183<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3137==mem[183])&&(Pass_182))
				Pass_183<=1;
			else
				Pass_183<=0;
		end

reg Pass_184;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_184<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3147==mem[184])&&(Pass_183))
				Pass_184<=1;
			else
				Pass_184<=0;
		end

reg Pass_185;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_185<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3207==mem[185])&&(Pass_184))
				Pass_185<=1;
			else
				Pass_185<=0;
		end

reg Pass_186;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_186<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3217==mem[186])&&(Pass_185))
				Pass_186<=1;
			else
				Pass_186<=0;
		end

reg Pass_187;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_187<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3227==mem[187])&&(Pass_186))
				Pass_187<=1;
			else
				Pass_187<=0;
		end

reg Pass_188;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_188<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3237==mem[188])&&(Pass_187))
				Pass_188<=1;
			else
				Pass_188<=0;
		end

reg Pass_189;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_189<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3247==mem[189])&&(Pass_188))
				Pass_189<=1;
			else
				Pass_189<=0;
		end

reg Pass_190;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_190<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3307==mem[190])&&(Pass_189))
				Pass_190<=1;
			else
				Pass_190<=0;
		end

reg Pass_191;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_191<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3317==mem[191])&&(Pass_190))
				Pass_191<=1;
			else
				Pass_191<=0;
		end

reg Pass_192;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_192<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3327==mem[192])&&(Pass_191))
				Pass_192<=1;
			else
				Pass_192<=0;
		end

reg Pass_193;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_193<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3337==mem[193])&&(Pass_192))
				Pass_193<=1;
			else
				Pass_193<=0;
		end

reg Pass_194;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_194<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3347==mem[194])&&(Pass_193))
				Pass_194<=1;
			else
				Pass_194<=0;
		end

reg Pass_195;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_195<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3407==mem[195])&&(Pass_194))
				Pass_195<=1;
			else
				Pass_195<=0;
		end

reg Pass_196;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_196<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3417==mem[196])&&(Pass_195))
				Pass_196<=1;
			else
				Pass_196<=0;
		end

reg Pass_197;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_197<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3427==mem[197])&&(Pass_196))
				Pass_197<=1;
			else
				Pass_197<=0;
		end

reg Pass_198;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_198<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3437==mem[198])&&(Pass_197))
				Pass_198<=1;
			else
				Pass_198<=0;
		end

reg Pass_199;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_199<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3447==mem[199])&&(Pass_198))
				Pass_199<=1;
			else
				Pass_199<=0;
		end

reg Pass_200;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_200<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3008==mem[200])&&(Pass_199))
				Pass_200<=1;
			else
				Pass_200<=0;
		end

reg Pass_201;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_201<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3018==mem[201])&&(Pass_200))
				Pass_201<=1;
			else
				Pass_201<=0;
		end

reg Pass_202;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_202<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3028==mem[202])&&(Pass_201))
				Pass_202<=1;
			else
				Pass_202<=0;
		end

reg Pass_203;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_203<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3038==mem[203])&&(Pass_202))
				Pass_203<=1;
			else
				Pass_203<=0;
		end

reg Pass_204;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_204<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3048==mem[204])&&(Pass_203))
				Pass_204<=1;
			else
				Pass_204<=0;
		end

reg Pass_205;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_205<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3108==mem[205])&&(Pass_204))
				Pass_205<=1;
			else
				Pass_205<=0;
		end

reg Pass_206;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_206<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3118==mem[206])&&(Pass_205))
				Pass_206<=1;
			else
				Pass_206<=0;
		end

reg Pass_207;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_207<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3128==mem[207])&&(Pass_206))
				Pass_207<=1;
			else
				Pass_207<=0;
		end

reg Pass_208;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_208<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3138==mem[208])&&(Pass_207))
				Pass_208<=1;
			else
				Pass_208<=0;
		end

reg Pass_209;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_209<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3148==mem[209])&&(Pass_208))
				Pass_209<=1;
			else
				Pass_209<=0;
		end

reg Pass_210;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_210<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3208==mem[210])&&(Pass_209))
				Pass_210<=1;
			else
				Pass_210<=0;
		end

reg Pass_211;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_211<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3218==mem[211])&&(Pass_210))
				Pass_211<=1;
			else
				Pass_211<=0;
		end

reg Pass_212;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_212<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3228==mem[212])&&(Pass_211))
				Pass_212<=1;
			else
				Pass_212<=0;
		end

reg Pass_213;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_213<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3238==mem[213])&&(Pass_212))
				Pass_213<=1;
			else
				Pass_213<=0;
		end

reg Pass_214;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_214<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3248==mem[214])&&(Pass_213))
				Pass_214<=1;
			else
				Pass_214<=0;
		end

reg Pass_215;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_215<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3308==mem[215])&&(Pass_214))
				Pass_215<=1;
			else
				Pass_215<=0;
		end

reg Pass_216;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_216<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3318==mem[216])&&(Pass_215))
				Pass_216<=1;
			else
				Pass_216<=0;
		end

reg Pass_217;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_217<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3328==mem[217])&&(Pass_216))
				Pass_217<=1;
			else
				Pass_217<=0;
		end

reg Pass_218;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_218<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3338==mem[218])&&(Pass_217))
				Pass_218<=1;
			else
				Pass_218<=0;
		end

reg Pass_219;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_219<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3348==mem[219])&&(Pass_218))
				Pass_219<=1;
			else
				Pass_219<=0;
		end

reg Pass_220;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_220<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3408==mem[220])&&(Pass_219))
				Pass_220<=1;
			else
				Pass_220<=0;
		end

reg Pass_221;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_221<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3418==mem[221])&&(Pass_220))
				Pass_221<=1;
			else
				Pass_221<=0;
		end

reg Pass_222;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_222<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3428==mem[222])&&(Pass_221))
				Pass_222<=1;
			else
				Pass_222<=0;
		end

reg Pass_223;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_223<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3438==mem[223])&&(Pass_222))
				Pass_223<=1;
			else
				Pass_223<=0;
		end

reg Pass_224;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_224<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3448==mem[224])&&(Pass_223))
				Pass_224<=1;
			else
				Pass_224<=0;
		end

reg Pass_225;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_225<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3009==mem[225])&&(Pass_224))
				Pass_225<=1;
			else
				Pass_225<=0;
		end

reg Pass_226;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_226<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3019==mem[226])&&(Pass_225))
				Pass_226<=1;
			else
				Pass_226<=0;
		end

reg Pass_227;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_227<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3029==mem[227])&&(Pass_226))
				Pass_227<=1;
			else
				Pass_227<=0;
		end

reg Pass_228;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_228<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3039==mem[228])&&(Pass_227))
				Pass_228<=1;
			else
				Pass_228<=0;
		end

reg Pass_229;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_229<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3049==mem[229])&&(Pass_228))
				Pass_229<=1;
			else
				Pass_229<=0;
		end

reg Pass_230;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_230<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3109==mem[230])&&(Pass_229))
				Pass_230<=1;
			else
				Pass_230<=0;
		end

reg Pass_231;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_231<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3119==mem[231])&&(Pass_230))
				Pass_231<=1;
			else
				Pass_231<=0;
		end

reg Pass_232;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_232<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3129==mem[232])&&(Pass_231))
				Pass_232<=1;
			else
				Pass_232<=0;
		end

reg Pass_233;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_233<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3139==mem[233])&&(Pass_232))
				Pass_233<=1;
			else
				Pass_233<=0;
		end

reg Pass_234;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_234<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3149==mem[234])&&(Pass_233))
				Pass_234<=1;
			else
				Pass_234<=0;
		end

reg Pass_235;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_235<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3209==mem[235])&&(Pass_234))
				Pass_235<=1;
			else
				Pass_235<=0;
		end

reg Pass_236;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_236<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3219==mem[236])&&(Pass_235))
				Pass_236<=1;
			else
				Pass_236<=0;
		end

reg Pass_237;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_237<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3229==mem[237])&&(Pass_236))
				Pass_237<=1;
			else
				Pass_237<=0;
		end

reg Pass_238;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_238<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3239==mem[238])&&(Pass_237))
				Pass_238<=1;
			else
				Pass_238<=0;
		end

reg Pass_239;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_239<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3249==mem[239])&&(Pass_238))
				Pass_239<=1;
			else
				Pass_239<=0;
		end

reg Pass_240;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_240<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3309==mem[240])&&(Pass_239))
				Pass_240<=1;
			else
				Pass_240<=0;
		end

reg Pass_241;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_241<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3319==mem[241])&&(Pass_240))
				Pass_241<=1;
			else
				Pass_241<=0;
		end

reg Pass_242;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_242<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3329==mem[242])&&(Pass_241))
				Pass_242<=1;
			else
				Pass_242<=0;
		end

reg Pass_243;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_243<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3339==mem[243])&&(Pass_242))
				Pass_243<=1;
			else
				Pass_243<=0;
		end

reg Pass_244;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_244<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3349==mem[244])&&(Pass_243))
				Pass_244<=1;
			else
				Pass_244<=0;
		end

reg Pass_245;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_245<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3409==mem[245])&&(Pass_244))
				Pass_245<=1;
			else
				Pass_245<=0;
		end

reg Pass_246;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_246<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3419==mem[246])&&(Pass_245))
				Pass_246<=1;
			else
				Pass_246<=0;
		end

reg Pass_247;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_247<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3429==mem[247])&&(Pass_246))
				Pass_247<=1;
			else
				Pass_247<=0;
		end

reg Pass_248;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_248<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3439==mem[248])&&(Pass_247))
				Pass_248<=1;
			else
				Pass_248<=0;
		end

reg Pass_249;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_249<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P3449==mem[249])&&(Pass_248))
				Pass_249<=1;
			else
				Pass_249<=0;
		end

reg Pass_250;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_250<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P300A==mem[250])&&(Pass_249))
				Pass_250<=1;
			else
				Pass_250<=0;
		end

reg Pass_251;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_251<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P301A==mem[251])&&(Pass_250))
				Pass_251<=1;
			else
				Pass_251<=0;
		end

reg Pass_252;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_252<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P302A==mem[252])&&(Pass_251))
				Pass_252<=1;
			else
				Pass_252<=0;
		end

reg Pass_253;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_253<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P303A==mem[253])&&(Pass_252))
				Pass_253<=1;
			else
				Pass_253<=0;
		end

reg Pass_254;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_254<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P304A==mem[254])&&(Pass_253))
				Pass_254<=1;
			else
				Pass_254<=0;
		end

reg Pass_255;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_255<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P310A==mem[255])&&(Pass_254))
				Pass_255<=1;
			else
				Pass_255<=0;
		end

reg Pass_256;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_256<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P311A==mem[256])&&(Pass_255))
				Pass_256<=1;
			else
				Pass_256<=0;
		end

reg Pass_257;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_257<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P312A==mem[257])&&(Pass_256))
				Pass_257<=1;
			else
				Pass_257<=0;
		end

reg Pass_258;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_258<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P313A==mem[258])&&(Pass_257))
				Pass_258<=1;
			else
				Pass_258<=0;
		end

reg Pass_259;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_259<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P314A==mem[259])&&(Pass_258))
				Pass_259<=1;
			else
				Pass_259<=0;
		end

reg Pass_260;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_260<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P320A==mem[260])&&(Pass_259))
				Pass_260<=1;
			else
				Pass_260<=0;
		end

reg Pass_261;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_261<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P321A==mem[261])&&(Pass_260))
				Pass_261<=1;
			else
				Pass_261<=0;
		end

reg Pass_262;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_262<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P322A==mem[262])&&(Pass_261))
				Pass_262<=1;
			else
				Pass_262<=0;
		end

reg Pass_263;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_263<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P323A==mem[263])&&(Pass_262))
				Pass_263<=1;
			else
				Pass_263<=0;
		end

reg Pass_264;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_264<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P324A==mem[264])&&(Pass_263))
				Pass_264<=1;
			else
				Pass_264<=0;
		end

reg Pass_265;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_265<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P330A==mem[265])&&(Pass_264))
				Pass_265<=1;
			else
				Pass_265<=0;
		end

reg Pass_266;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_266<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P331A==mem[266])&&(Pass_265))
				Pass_266<=1;
			else
				Pass_266<=0;
		end

reg Pass_267;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_267<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P332A==mem[267])&&(Pass_266))
				Pass_267<=1;
			else
				Pass_267<=0;
		end

reg Pass_268;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_268<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P333A==mem[268])&&(Pass_267))
				Pass_268<=1;
			else
				Pass_268<=0;
		end

reg Pass_269;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_269<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P334A==mem[269])&&(Pass_268))
				Pass_269<=1;
			else
				Pass_269<=0;
		end

reg Pass_270;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_270<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P340A==mem[270])&&(Pass_269))
				Pass_270<=1;
			else
				Pass_270<=0;
		end

reg Pass_271;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_271<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P341A==mem[271])&&(Pass_270))
				Pass_271<=1;
			else
				Pass_271<=0;
		end

reg Pass_272;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_272<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P342A==mem[272])&&(Pass_271))
				Pass_272<=1;
			else
				Pass_272<=0;
		end

reg Pass_273;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_273<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P343A==mem[273])&&(Pass_272))
				Pass_273<=1;
			else
				Pass_273<=0;
		end

reg Pass_274;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_274<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P344A==mem[274])&&(Pass_273))
				Pass_274<=1;
			else
				Pass_274<=0;
		end

reg Pass_275;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_275<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P300B==mem[275])&&(Pass_274))
				Pass_275<=1;
			else
				Pass_275<=0;
		end

reg Pass_276;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_276<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P301B==mem[276])&&(Pass_275))
				Pass_276<=1;
			else
				Pass_276<=0;
		end

reg Pass_277;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_277<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P302B==mem[277])&&(Pass_276))
				Pass_277<=1;
			else
				Pass_277<=0;
		end

reg Pass_278;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_278<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P303B==mem[278])&&(Pass_277))
				Pass_278<=1;
			else
				Pass_278<=0;
		end

reg Pass_279;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_279<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P304B==mem[279])&&(Pass_278))
				Pass_279<=1;
			else
				Pass_279<=0;
		end

reg Pass_280;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_280<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P310B==mem[280])&&(Pass_279))
				Pass_280<=1;
			else
				Pass_280<=0;
		end

reg Pass_281;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_281<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P311B==mem[281])&&(Pass_280))
				Pass_281<=1;
			else
				Pass_281<=0;
		end

reg Pass_282;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_282<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P312B==mem[282])&&(Pass_281))
				Pass_282<=1;
			else
				Pass_282<=0;
		end

reg Pass_283;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_283<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P313B==mem[283])&&(Pass_282))
				Pass_283<=1;
			else
				Pass_283<=0;
		end

reg Pass_284;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_284<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P314B==mem[284])&&(Pass_283))
				Pass_284<=1;
			else
				Pass_284<=0;
		end

reg Pass_285;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_285<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P320B==mem[285])&&(Pass_284))
				Pass_285<=1;
			else
				Pass_285<=0;
		end

reg Pass_286;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_286<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P321B==mem[286])&&(Pass_285))
				Pass_286<=1;
			else
				Pass_286<=0;
		end

reg Pass_287;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_287<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P322B==mem[287])&&(Pass_286))
				Pass_287<=1;
			else
				Pass_287<=0;
		end

reg Pass_288;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_288<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P323B==mem[288])&&(Pass_287))
				Pass_288<=1;
			else
				Pass_288<=0;
		end

reg Pass_289;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_289<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P324B==mem[289])&&(Pass_288))
				Pass_289<=1;
			else
				Pass_289<=0;
		end

reg Pass_290;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_290<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P330B==mem[290])&&(Pass_289))
				Pass_290<=1;
			else
				Pass_290<=0;
		end

reg Pass_291;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_291<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P331B==mem[291])&&(Pass_290))
				Pass_291<=1;
			else
				Pass_291<=0;
		end

reg Pass_292;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_292<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P332B==mem[292])&&(Pass_291))
				Pass_292<=1;
			else
				Pass_292<=0;
		end

reg Pass_293;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_293<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P333B==mem[293])&&(Pass_292))
				Pass_293<=1;
			else
				Pass_293<=0;
		end

reg Pass_294;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_294<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P334B==mem[294])&&(Pass_293))
				Pass_294<=1;
			else
				Pass_294<=0;
		end

reg Pass_295;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_295<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P340B==mem[295])&&(Pass_294))
				Pass_295<=1;
			else
				Pass_295<=0;
		end

reg Pass_296;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_296<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P341B==mem[296])&&(Pass_295))
				Pass_296<=1;
			else
				Pass_296<=0;
		end

reg Pass_297;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_297<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P342B==mem[297])&&(Pass_296))
				Pass_297<=1;
			else
				Pass_297<=0;
		end

reg Pass_298;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_298<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P343B==mem[298])&&(Pass_297))
				Pass_298<=1;
			else
				Pass_298<=0;
		end

reg Pass_299;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_299<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P344B==mem[299])&&(Pass_298))
				Pass_299<=1;
			else
				Pass_299<=0;
		end

reg Pass_300;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_300<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P300C==mem[300])&&(Pass_299))
				Pass_300<=1;
			else
				Pass_300<=0;
		end

reg Pass_301;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_301<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P301C==mem[301])&&(Pass_300))
				Pass_301<=1;
			else
				Pass_301<=0;
		end

reg Pass_302;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_302<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P302C==mem[302])&&(Pass_301))
				Pass_302<=1;
			else
				Pass_302<=0;
		end

reg Pass_303;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_303<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P303C==mem[303])&&(Pass_302))
				Pass_303<=1;
			else
				Pass_303<=0;
		end

reg Pass_304;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_304<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P304C==mem[304])&&(Pass_303))
				Pass_304<=1;
			else
				Pass_304<=0;
		end

reg Pass_305;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_305<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P310C==mem[305])&&(Pass_304))
				Pass_305<=1;
			else
				Pass_305<=0;
		end

reg Pass_306;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_306<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P311C==mem[306])&&(Pass_305))
				Pass_306<=1;
			else
				Pass_306<=0;
		end

reg Pass_307;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_307<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P312C==mem[307])&&(Pass_306))
				Pass_307<=1;
			else
				Pass_307<=0;
		end

reg Pass_308;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_308<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P313C==mem[308])&&(Pass_307))
				Pass_308<=1;
			else
				Pass_308<=0;
		end

reg Pass_309;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_309<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P314C==mem[309])&&(Pass_308))
				Pass_309<=1;
			else
				Pass_309<=0;
		end

reg Pass_310;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_310<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P320C==mem[310])&&(Pass_309))
				Pass_310<=1;
			else
				Pass_310<=0;
		end

reg Pass_311;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_311<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P321C==mem[311])&&(Pass_310))
				Pass_311<=1;
			else
				Pass_311<=0;
		end

reg Pass_312;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_312<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P322C==mem[312])&&(Pass_311))
				Pass_312<=1;
			else
				Pass_312<=0;
		end

reg Pass_313;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_313<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P323C==mem[313])&&(Pass_312))
				Pass_313<=1;
			else
				Pass_313<=0;
		end

reg Pass_314;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_314<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P324C==mem[314])&&(Pass_313))
				Pass_314<=1;
			else
				Pass_314<=0;
		end

reg Pass_315;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_315<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P330C==mem[315])&&(Pass_314))
				Pass_315<=1;
			else
				Pass_315<=0;
		end

reg Pass_316;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_316<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P331C==mem[316])&&(Pass_315))
				Pass_316<=1;
			else
				Pass_316<=0;
		end

reg Pass_317;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_317<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P332C==mem[317])&&(Pass_316))
				Pass_317<=1;
			else
				Pass_317<=0;
		end

reg Pass_318;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_318<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P333C==mem[318])&&(Pass_317))
				Pass_318<=1;
			else
				Pass_318<=0;
		end

reg Pass_319;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_319<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P334C==mem[319])&&(Pass_318))
				Pass_319<=1;
			else
				Pass_319<=0;
		end

reg Pass_320;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_320<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P340C==mem[320])&&(Pass_319))
				Pass_320<=1;
			else
				Pass_320<=0;
		end

reg Pass_321;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_321<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P341C==mem[321])&&(Pass_320))
				Pass_321<=1;
			else
				Pass_321<=0;
		end

reg Pass_322;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_322<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P342C==mem[322])&&(Pass_321))
				Pass_322<=1;
			else
				Pass_322<=0;
		end

reg Pass_323;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_323<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P343C==mem[323])&&(Pass_322))
				Pass_323<=1;
			else
				Pass_323<=0;
		end

reg Pass_324;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_324<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P344C==mem[324])&&(Pass_323))
				Pass_324<=1;
			else
				Pass_324<=0;
		end

reg Pass_325;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_325<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P300D==mem[325])&&(Pass_324))
				Pass_325<=1;
			else
				Pass_325<=0;
		end

reg Pass_326;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_326<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P301D==mem[326])&&(Pass_325))
				Pass_326<=1;
			else
				Pass_326<=0;
		end

reg Pass_327;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_327<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P302D==mem[327])&&(Pass_326))
				Pass_327<=1;
			else
				Pass_327<=0;
		end

reg Pass_328;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_328<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P303D==mem[328])&&(Pass_327))
				Pass_328<=1;
			else
				Pass_328<=0;
		end

reg Pass_329;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_329<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P304D==mem[329])&&(Pass_328))
				Pass_329<=1;
			else
				Pass_329<=0;
		end

reg Pass_330;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_330<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P310D==mem[330])&&(Pass_329))
				Pass_330<=1;
			else
				Pass_330<=0;
		end

reg Pass_331;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_331<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P311D==mem[331])&&(Pass_330))
				Pass_331<=1;
			else
				Pass_331<=0;
		end

reg Pass_332;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_332<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P312D==mem[332])&&(Pass_331))
				Pass_332<=1;
			else
				Pass_332<=0;
		end

reg Pass_333;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_333<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P313D==mem[333])&&(Pass_332))
				Pass_333<=1;
			else
				Pass_333<=0;
		end

reg Pass_334;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_334<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P314D==mem[334])&&(Pass_333))
				Pass_334<=1;
			else
				Pass_334<=0;
		end

reg Pass_335;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_335<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P320D==mem[335])&&(Pass_334))
				Pass_335<=1;
			else
				Pass_335<=0;
		end

reg Pass_336;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_336<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P321D==mem[336])&&(Pass_335))
				Pass_336<=1;
			else
				Pass_336<=0;
		end

reg Pass_337;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_337<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P322D==mem[337])&&(Pass_336))
				Pass_337<=1;
			else
				Pass_337<=0;
		end

reg Pass_338;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_338<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P323D==mem[338])&&(Pass_337))
				Pass_338<=1;
			else
				Pass_338<=0;
		end

reg Pass_339;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_339<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P324D==mem[339])&&(Pass_338))
				Pass_339<=1;
			else
				Pass_339<=0;
		end

reg Pass_340;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_340<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P330D==mem[340])&&(Pass_339))
				Pass_340<=1;
			else
				Pass_340<=0;
		end

reg Pass_341;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_341<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P331D==mem[341])&&(Pass_340))
				Pass_341<=1;
			else
				Pass_341<=0;
		end

reg Pass_342;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_342<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P332D==mem[342])&&(Pass_341))
				Pass_342<=1;
			else
				Pass_342<=0;
		end

reg Pass_343;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_343<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P333D==mem[343])&&(Pass_342))
				Pass_343<=1;
			else
				Pass_343<=0;
		end

reg Pass_344;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_344<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P334D==mem[344])&&(Pass_343))
				Pass_344<=1;
			else
				Pass_344<=0;
		end

reg Pass_345;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_345<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P340D==mem[345])&&(Pass_344))
				Pass_345<=1;
			else
				Pass_345<=0;
		end

reg Pass_346;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_346<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P341D==mem[346])&&(Pass_345))
				Pass_346<=1;
			else
				Pass_346<=0;
		end

reg Pass_347;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_347<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P342D==mem[347])&&(Pass_346))
				Pass_347<=1;
			else
				Pass_347<=0;
		end

reg Pass_348;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_348<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P343D==mem[348])&&(Pass_347))
				Pass_348<=1;
			else
				Pass_348<=0;
		end

reg Pass_349;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_349<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P344D==mem[349])&&(Pass_348))
				Pass_349<=1;
			else
				Pass_349<=0;
		end

reg Pass_350;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_350<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P300E==mem[350])&&(Pass_349))
				Pass_350<=1;
			else
				Pass_350<=0;
		end

reg Pass_351;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_351<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P301E==mem[351])&&(Pass_350))
				Pass_351<=1;
			else
				Pass_351<=0;
		end

reg Pass_352;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_352<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P302E==mem[352])&&(Pass_351))
				Pass_352<=1;
			else
				Pass_352<=0;
		end

reg Pass_353;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_353<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P303E==mem[353])&&(Pass_352))
				Pass_353<=1;
			else
				Pass_353<=0;
		end

reg Pass_354;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_354<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P304E==mem[354])&&(Pass_353))
				Pass_354<=1;
			else
				Pass_354<=0;
		end

reg Pass_355;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_355<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P310E==mem[355])&&(Pass_354))
				Pass_355<=1;
			else
				Pass_355<=0;
		end

reg Pass_356;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_356<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P311E==mem[356])&&(Pass_355))
				Pass_356<=1;
			else
				Pass_356<=0;
		end

reg Pass_357;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_357<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P312E==mem[357])&&(Pass_356))
				Pass_357<=1;
			else
				Pass_357<=0;
		end

reg Pass_358;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_358<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P313E==mem[358])&&(Pass_357))
				Pass_358<=1;
			else
				Pass_358<=0;
		end

reg Pass_359;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_359<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P314E==mem[359])&&(Pass_358))
				Pass_359<=1;
			else
				Pass_359<=0;
		end

reg Pass_360;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_360<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P320E==mem[360])&&(Pass_359))
				Pass_360<=1;
			else
				Pass_360<=0;
		end

reg Pass_361;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_361<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P321E==mem[361])&&(Pass_360))
				Pass_361<=1;
			else
				Pass_361<=0;
		end

reg Pass_362;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_362<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P322E==mem[362])&&(Pass_361))
				Pass_362<=1;
			else
				Pass_362<=0;
		end

reg Pass_363;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_363<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P323E==mem[363])&&(Pass_362))
				Pass_363<=1;
			else
				Pass_363<=0;
		end

reg Pass_364;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_364<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P324E==mem[364])&&(Pass_363))
				Pass_364<=1;
			else
				Pass_364<=0;
		end

reg Pass_365;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_365<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P330E==mem[365])&&(Pass_364))
				Pass_365<=1;
			else
				Pass_365<=0;
		end

reg Pass_366;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_366<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P331E==mem[366])&&(Pass_365))
				Pass_366<=1;
			else
				Pass_366<=0;
		end

reg Pass_367;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_367<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P332E==mem[367])&&(Pass_366))
				Pass_367<=1;
			else
				Pass_367<=0;
		end

reg Pass_368;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_368<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P333E==mem[368])&&(Pass_367))
				Pass_368<=1;
			else
				Pass_368<=0;
		end

reg Pass_369;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_369<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P334E==mem[369])&&(Pass_368))
				Pass_369<=1;
			else
				Pass_369<=0;
		end

reg Pass_370;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_370<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P340E==mem[370])&&(Pass_369))
				Pass_370<=1;
			else
				Pass_370<=0;
		end

reg Pass_371;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_371<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P341E==mem[371])&&(Pass_370))
				Pass_371<=1;
			else
				Pass_371<=0;
		end

reg Pass_372;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_372<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P342E==mem[372])&&(Pass_371))
				Pass_372<=1;
			else
				Pass_372<=0;
		end

reg Pass_373;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_373<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P343E==mem[373])&&(Pass_372))
				Pass_373<=1;
			else
				Pass_373<=0;
		end

reg Pass_374;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_374<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P344E==mem[374])&&(Pass_373))
				Pass_374<=1;
			else
				Pass_374<=0;
		end

reg Pass_375;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_375<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P300F==mem[375])&&(Pass_374))
				Pass_375<=1;
			else
				Pass_375<=0;
		end

reg Pass_376;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_376<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P301F==mem[376])&&(Pass_375))
				Pass_376<=1;
			else
				Pass_376<=0;
		end

reg Pass_377;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_377<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P302F==mem[377])&&(Pass_376))
				Pass_377<=1;
			else
				Pass_377<=0;
		end

reg Pass_378;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_378<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P303F==mem[378])&&(Pass_377))
				Pass_378<=1;
			else
				Pass_378<=0;
		end

reg Pass_379;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_379<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P304F==mem[379])&&(Pass_378))
				Pass_379<=1;
			else
				Pass_379<=0;
		end

reg Pass_380;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_380<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P310F==mem[380])&&(Pass_379))
				Pass_380<=1;
			else
				Pass_380<=0;
		end

reg Pass_381;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_381<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P311F==mem[381])&&(Pass_380))
				Pass_381<=1;
			else
				Pass_381<=0;
		end

reg Pass_382;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_382<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P312F==mem[382])&&(Pass_381))
				Pass_382<=1;
			else
				Pass_382<=0;
		end

reg Pass_383;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_383<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P313F==mem[383])&&(Pass_382))
				Pass_383<=1;
			else
				Pass_383<=0;
		end

reg Pass_384;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_384<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P314F==mem[384])&&(Pass_383))
				Pass_384<=1;
			else
				Pass_384<=0;
		end

reg Pass_385;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_385<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P320F==mem[385])&&(Pass_384))
				Pass_385<=1;
			else
				Pass_385<=0;
		end

reg Pass_386;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_386<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P321F==mem[386])&&(Pass_385))
				Pass_386<=1;
			else
				Pass_386<=0;
		end

reg Pass_387;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_387<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P322F==mem[387])&&(Pass_386))
				Pass_387<=1;
			else
				Pass_387<=0;
		end

reg Pass_388;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_388<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P323F==mem[388])&&(Pass_387))
				Pass_388<=1;
			else
				Pass_388<=0;
		end

reg Pass_389;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_389<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P324F==mem[389])&&(Pass_388))
				Pass_389<=1;
			else
				Pass_389<=0;
		end

reg Pass_390;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_390<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P330F==mem[390])&&(Pass_389))
				Pass_390<=1;
			else
				Pass_390<=0;
		end

reg Pass_391;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_391<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P331F==mem[391])&&(Pass_390))
				Pass_391<=1;
			else
				Pass_391<=0;
		end

reg Pass_392;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_392<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P332F==mem[392])&&(Pass_391))
				Pass_392<=1;
			else
				Pass_392<=0;
		end

reg Pass_393;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_393<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P333F==mem[393])&&(Pass_392))
				Pass_393<=1;
			else
				Pass_393<=0;
		end

reg Pass_394;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_394<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P334F==mem[394])&&(Pass_393))
				Pass_394<=1;
			else
				Pass_394<=0;
		end

reg Pass_395;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_395<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P340F==mem[395])&&(Pass_394))
				Pass_395<=1;
			else
				Pass_395<=0;
		end

reg Pass_396;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_396<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P341F==mem[396])&&(Pass_395))
				Pass_396<=1;
			else
				Pass_396<=0;
		end

reg Pass_397;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_397<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P342F==mem[397])&&(Pass_396))
				Pass_397<=1;
			else
				Pass_397<=0;
		end

reg Pass_398;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_398<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P343F==mem[398])&&(Pass_397))
				Pass_398<=1;
			else
				Pass_398<=0;
		end

reg Pass_399;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_399<=0;
	else if(count>=2)
		begin
			if((tb_test_layer2.test_layer2.P344F==mem[399])&&(Pass_398))
				Pass_399<=1;
			else
				Pass_399<=0;
		end

always@(posedge clk)
if(Pass_0&&Pass_1&&Pass_2&&Pass_3&&Pass_4&&Pass_5&&Pass_6&&Pass_7&&Pass_8&&Pass_9&&Pass_10&&Pass_11&&Pass_12&&Pass_13&&Pass_14&&Pass_15&&Pass_16&&Pass_17&&Pass_18&&Pass_19&&Pass_20&&Pass_21&&Pass_22&&Pass_23&&Pass_24&&Pass_25&&Pass_26&&Pass_27&&Pass_28&&Pass_29&&Pass_30&&Pass_31&&Pass_32&&Pass_33&&Pass_34&&Pass_35&&Pass_36&&Pass_37&&Pass_38&&Pass_39&&Pass_40&&Pass_41&&Pass_42&&Pass_43&&Pass_44&&Pass_45&&Pass_46&&Pass_47&&Pass_48&&Pass_49&&Pass_50&&Pass_51&&Pass_52&&Pass_53&&Pass_54&&Pass_55&&Pass_56&&Pass_57&&Pass_58&&Pass_59&&Pass_60&&Pass_61&&Pass_62&&Pass_63&&Pass_64&&Pass_65&&Pass_66&&Pass_67&&Pass_68&&Pass_69&&Pass_70&&Pass_71&&Pass_72&&Pass_73&&Pass_74&&Pass_75&&Pass_76&&Pass_77&&Pass_78&&Pass_79&&Pass_80&&Pass_81&&Pass_82&&Pass_83&&Pass_84&&Pass_85&&Pass_86&&Pass_87&&Pass_88&&Pass_89&&Pass_90&&Pass_91&&Pass_92&&Pass_93&&Pass_94&&Pass_95&&Pass_96&&Pass_97&&Pass_98&&Pass_99&&Pass_100&&Pass_101&&Pass_102&&Pass_103&&Pass_104&&Pass_105&&Pass_106&&Pass_107&&Pass_108&&Pass_109&&Pass_110&&Pass_111&&Pass_112&&Pass_113&&Pass_114&&Pass_115&&Pass_116&&Pass_117&&Pass_118&&Pass_119&&Pass_120&&Pass_121&&Pass_122&&Pass_123&&Pass_124&&Pass_125&&Pass_126&&Pass_127&&Pass_128&&Pass_129&&Pass_130&&Pass_131&&Pass_132&&Pass_133&&Pass_134&&Pass_135&&Pass_136&&Pass_137&&Pass_138&&Pass_139&&Pass_140&&Pass_141&&Pass_142&&Pass_143&&Pass_144&&Pass_145&&Pass_146&&Pass_147&&Pass_148&&Pass_149&&Pass_150&&Pass_151&&Pass_152&&Pass_153&&Pass_154&&Pass_155&&Pass_156&&Pass_157&&Pass_158&&Pass_159&&Pass_160&&Pass_161&&Pass_162&&Pass_163&&Pass_164&&Pass_165&&Pass_166&&Pass_167&&Pass_168&&Pass_169&&Pass_170&&Pass_171&&Pass_172&&Pass_173&&Pass_174&&Pass_175&&Pass_176&&Pass_177&&Pass_178&&Pass_179&&Pass_180&&Pass_181&&Pass_182&&Pass_183&&Pass_184&&Pass_185&&Pass_186&&Pass_187&&Pass_188&&Pass_189&&Pass_190&&Pass_191&&Pass_192&&Pass_193&&Pass_194&&Pass_195&&Pass_196&&Pass_197&&Pass_198&&Pass_199&&Pass_200&&Pass_201&&Pass_202&&Pass_203&&Pass_204&&Pass_205&&Pass_206&&Pass_207&&Pass_208&&Pass_209&&Pass_210&&Pass_211&&Pass_212&&Pass_213&&Pass_214&&Pass_215&&Pass_216&&Pass_217&&Pass_218&&Pass_219&&Pass_220&&Pass_221&&Pass_222&&Pass_223&&Pass_224&&Pass_225&&Pass_226&&Pass_227&&Pass_228&&Pass_229&&Pass_230&&Pass_231&&Pass_232&&Pass_233&&Pass_234&&Pass_235&&Pass_236&&Pass_237&&Pass_238&&Pass_239&&Pass_240&&Pass_241&&Pass_242&&Pass_243&&Pass_244&&Pass_245&&Pass_246&&Pass_247&&Pass_248&&Pass_249&&Pass_250&&Pass_251&&Pass_252&&Pass_253&&Pass_254&&Pass_255&&Pass_256&&Pass_257&&Pass_258&&Pass_259&&Pass_260&&Pass_261&&Pass_262&&Pass_263&&Pass_264&&Pass_265&&Pass_266&&Pass_267&&Pass_268&&Pass_269&&Pass_270&&Pass_271&&Pass_272&&Pass_273&&Pass_274&&Pass_275&&Pass_276&&Pass_277&&Pass_278&&Pass_279&&Pass_280&&Pass_281&&Pass_282&&Pass_283&&Pass_284&&Pass_285&&Pass_286&&Pass_287&&Pass_288&&Pass_289&&Pass_290&&Pass_291&&Pass_292&&Pass_293&&Pass_294&&Pass_295&&Pass_296&&Pass_297&&Pass_298&&Pass_299&&Pass_300&&Pass_301&&Pass_302&&Pass_303&&Pass_304&&Pass_305&&Pass_306&&Pass_307&&Pass_308&&Pass_309&&Pass_310&&Pass_311&&Pass_312&&Pass_313&&Pass_314&&Pass_315&&Pass_316&&Pass_317&&Pass_318&&Pass_319&&Pass_320&&Pass_321&&Pass_322&&Pass_323&&Pass_324&&Pass_325&&Pass_326&&Pass_327&&Pass_328&&Pass_329&&Pass_330&&Pass_331&&Pass_332&&Pass_333&&Pass_334&&Pass_335&&Pass_336&&Pass_337&&Pass_338&&Pass_339&&Pass_340&&Pass_341&&Pass_342&&Pass_343&&Pass_344&&Pass_345&&Pass_346&&Pass_347&&Pass_348&&Pass_349&&Pass_350&&Pass_351&&Pass_352&&Pass_353&&Pass_354&&Pass_355&&Pass_356&&Pass_357&&Pass_358&&Pass_359&&Pass_360&&Pass_361&&Pass_362&&Pass_363&&Pass_364&&Pass_365&&Pass_366&&Pass_367&&Pass_368&&Pass_369&&Pass_370&&Pass_371&&Pass_372&&Pass_373&&Pass_374&&Pass_375&&Pass_376&&Pass_377&&Pass_378&&Pass_379&&Pass_380&&Pass_381&&Pass_382&&Pass_383&&Pass_384&&Pass_385&&Pass_386&&Pass_387&&Pass_388&&Pass_389&&Pass_390&&Pass_391&&Pass_392&&Pass_393&&Pass_394&&Pass_395&&Pass_396&&Pass_397&&Pass_398&&Pass_399)
begin
$display("PASS");
$finish;
end

endmodule
